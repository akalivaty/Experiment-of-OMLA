//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n560, new_n561, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n631, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OR2_X1    g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g043(.A(KEYINPUT3), .B(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(G137), .A3(new_n461), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n468), .A2(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n469), .A2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  AND2_X1   g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  NOR2_X1   g060(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n486));
  OAI211_X1 g061(.A(G138), .B(new_n461), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n469), .A2(new_n489), .A3(G138), .A4(new_n461), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(G126), .A2(G2105), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n492), .B1(new_n463), .B2(new_n464), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n461), .A2(G114), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT66), .ZN(new_n497));
  NOR3_X1   g072(.A1(new_n493), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  OAI211_X1 g073(.A(G126), .B(G2105), .C1(new_n485), .C2(new_n486), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(G114), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(G2105), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n500), .A2(new_n502), .A3(G2104), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT66), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n491), .B1(new_n498), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT67), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n497), .B1(new_n493), .B2(new_n496), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n499), .A2(new_n503), .A3(KEYINPUT66), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(KEYINPUT67), .A3(new_n491), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n507), .A2(new_n511), .ZN(G164));
  OR2_X1    g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OR2_X1    g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  NOR2_X1   g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  AND2_X1   g099(.A1(KEYINPUT5), .A2(G543), .ZN(new_n525));
  AND2_X1   g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n524), .A2(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G88), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n522), .A2(new_n523), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT68), .ZN(new_n531));
  OR3_X1    g106(.A1(new_n518), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n518), .B2(new_n530), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(G166));
  INV_X1    g109(.A(G543), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n535), .B1(new_n519), .B2(new_n520), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT69), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n537), .A2(G51), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n539));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT7), .ZN(new_n541));
  INV_X1    g116(.A(G89), .ZN(new_n542));
  OAI211_X1 g117(.A(new_n539), .B(new_n541), .C1(new_n542), .C2(new_n528), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n538), .A2(new_n543), .ZN(G168));
  AND2_X1   g119(.A1(new_n537), .A2(G52), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  INV_X1    g121(.A(G90), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n546), .A2(new_n517), .B1(new_n547), .B2(new_n528), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(G171));
  AOI22_X1  g124(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n517), .ZN(new_n551));
  INV_X1    g126(.A(new_n528), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n551), .A2(KEYINPUT70), .B1(G81), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n537), .A2(G43), .ZN(new_n554));
  OAI211_X1 g129(.A(new_n553), .B(new_n554), .C1(KEYINPUT70), .C2(new_n551), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT71), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  INV_X1    g137(.A(KEYINPUT73), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n528), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n515), .A2(new_n521), .A3(KEYINPUT73), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n564), .A2(G91), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT72), .ZN(new_n567));
  INV_X1    g142(.A(G53), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n567), .B(KEYINPUT9), .C1(new_n522), .C2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(KEYINPUT9), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n536), .A2(G53), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n515), .A2(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n525), .A2(new_n524), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT74), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n566), .B(new_n572), .C1(new_n578), .C2(new_n517), .ZN(G299));
  OR2_X1    g154(.A1(new_n545), .A2(new_n548), .ZN(G301));
  INV_X1    g155(.A(G168), .ZN(G286));
  INV_X1    g156(.A(G166), .ZN(G303));
  NAND3_X1  g157(.A1(new_n564), .A2(G87), .A3(new_n565), .ZN(new_n583));
  INV_X1    g158(.A(G74), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n575), .A2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(new_n536), .B2(G49), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT75), .ZN(G288));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n513), .B2(new_n514), .ZN(new_n590));
  INV_X1    g165(.A(G73), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n591), .A2(new_n535), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n594));
  AOI21_X1  g169(.A(new_n594), .B1(new_n536), .B2(G48), .ZN(new_n595));
  OAI211_X1 g170(.A(G48), .B(G543), .C1(new_n526), .C2(new_n527), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n596), .A2(KEYINPUT77), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n593), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n564), .A2(G86), .A3(new_n565), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT76), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g176(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT76), .A4(G86), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n598), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G305));
  NAND2_X1  g179(.A1(new_n537), .A2(G47), .ZN(new_n605));
  NAND2_X1  g180(.A1(G72), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G60), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n575), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(G651), .A2(new_n608), .B1(new_n552), .B2(G85), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n605), .A2(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  AND2_X1   g186(.A1(new_n577), .A2(G66), .ZN(new_n612));
  AND2_X1   g187(.A1(G79), .A2(G543), .ZN(new_n613));
  OAI21_X1  g188(.A(G651), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n537), .A2(G54), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT79), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n614), .A2(KEYINPUT79), .A3(new_n615), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n564), .A2(G92), .A3(new_n565), .ZN(new_n621));
  XOR2_X1   g196(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  AND2_X1   g198(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n611), .B1(new_n624), .B2(G868), .ZN(G284));
  OAI21_X1  g200(.A(new_n611), .B1(new_n624), .B2(G868), .ZN(G321));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(G299), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n628), .B1(new_n627), .B2(G168), .ZN(G297));
  OAI21_X1  g204(.A(new_n628), .B1(new_n627), .B2(G168), .ZN(G280));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n624), .B1(new_n631), .B2(G860), .ZN(G148));
  NAND2_X1  g207(.A1(new_n624), .A2(new_n631), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G868), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n469), .A2(new_n472), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  INV_X1    g215(.A(G2100), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n479), .A2(G135), .ZN(new_n644));
  OR2_X1    g219(.A1(G99), .A2(G2105), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n645), .B(G2104), .C1(G111), .C2(new_n461), .ZN(new_n646));
  INV_X1    g221(.A(G123), .ZN(new_n647));
  OAI211_X1 g222(.A(new_n644), .B(new_n646), .C1(new_n647), .C2(new_n476), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2096), .Z(new_n649));
  NAND3_X1  g224(.A1(new_n642), .A2(new_n643), .A3(new_n649), .ZN(G156));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(KEYINPUT14), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT82), .Z(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n660), .B(new_n661), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n657), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(new_n666), .A3(G14), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G401));
  XNOR2_X1  g243(.A(G2072), .B(G2078), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT17), .Z(new_n670));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(new_n671), .B2(new_n669), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT83), .Z(new_n678));
  NAND3_X1  g253(.A1(new_n674), .A2(new_n671), .A3(new_n669), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT18), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n675), .A2(new_n671), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n680), .B1(new_n670), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G2096), .B(G2100), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1956), .B(G2474), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1961), .B(G1966), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NOR3_X1   g266(.A1(new_n687), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n687), .A2(new_n690), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT20), .Z(new_n694));
  AOI211_X1 g269(.A(new_n692), .B(new_n694), .C1(new_n687), .C2(new_n691), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1981), .B(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(G229));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G22), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT87), .Z(new_n704));
  OAI21_X1  g279(.A(new_n704), .B1(G166), .B2(new_n702), .ZN(new_n705));
  INV_X1    g280(.A(G1971), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n702), .A2(G6), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(new_n603), .B2(new_n702), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT32), .B(G1981), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n587), .A2(KEYINPUT86), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT86), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n583), .A2(new_n714), .A3(new_n586), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n713), .A2(G16), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G16), .B2(G23), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT33), .B(G1976), .Z(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n717), .A2(new_n719), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n720), .B(new_n721), .C1(new_n710), .C2(new_n709), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n712), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT85), .B(KEYINPUT34), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  MUX2_X1   g300(.A(G24), .B(G290), .S(G16), .Z(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(G1986), .Z(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT84), .B(G29), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(G25), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n477), .A2(G119), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n479), .A2(G131), .ZN(new_n732));
  OR2_X1    g307(.A1(G95), .A2(G2105), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n733), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n731), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n730), .B1(new_n736), .B2(new_n729), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT35), .B(G1991), .Z(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n725), .A2(new_n727), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT88), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n724), .B2(new_n723), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT36), .Z(new_n743));
  NAND2_X1  g318(.A1(new_n479), .A2(G140), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n461), .A2(G116), .ZN(new_n745));
  OAI21_X1  g320(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n746));
  INV_X1    g321(.A(G128), .ZN(new_n747));
  OAI221_X1 g322(.A(new_n744), .B1(new_n745), .B2(new_n746), .C1(new_n747), .C2(new_n476), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G29), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n728), .A2(G26), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT28), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G2067), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G171), .A2(new_n702), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G5), .B2(new_n702), .ZN(new_n756));
  INV_X1    g331(.A(G1961), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n754), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OR2_X1    g333(.A1(KEYINPUT30), .A2(G28), .ZN(new_n759));
  NAND2_X1  g334(.A1(KEYINPUT30), .A2(G28), .ZN(new_n760));
  AOI21_X1  g335(.A(G29), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT31), .B(G11), .Z(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n648), .A2(new_n728), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT24), .B(G34), .ZN(new_n765));
  AOI22_X1  g340(.A1(G160), .A2(G29), .B1(new_n728), .B2(new_n765), .ZN(new_n766));
  AOI211_X1 g341(.A(new_n763), .B(new_n764), .C1(G2084), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(G162), .A2(new_n729), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G35), .B2(new_n729), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT29), .Z(new_n770));
  OAI221_X1 g345(.A(new_n767), .B1(G2084), .B2(new_n766), .C1(new_n770), .C2(G2090), .ZN(new_n771));
  AOI211_X1 g346(.A(new_n758), .B(new_n771), .C1(new_n757), .C2(new_n756), .ZN(new_n772));
  INV_X1    g347(.A(G29), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(G32), .ZN(new_n774));
  NAND3_X1  g349(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT26), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n479), .A2(G141), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n472), .A2(G105), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AOI211_X1 g354(.A(new_n776), .B(new_n779), .C1(G129), .C2(new_n477), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n774), .B1(new_n780), .B2(new_n773), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT27), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1996), .ZN(new_n783));
  NAND2_X1  g358(.A1(G168), .A2(G16), .ZN(new_n784));
  NOR2_X1   g359(.A1(G16), .A2(G21), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(KEYINPUT92), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(KEYINPUT92), .B2(new_n784), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1966), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n772), .A2(new_n783), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n773), .A2(G33), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n469), .A2(G127), .ZN(new_n791));
  INV_X1    g366(.A(G115), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(new_n471), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n461), .B1(new_n793), .B2(KEYINPUT90), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(KEYINPUT90), .B2(new_n793), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT25), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  AOI22_X1  g374(.A1(new_n798), .A2(new_n799), .B1(new_n479), .B2(G139), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n790), .B1(new_n802), .B2(new_n773), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT91), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(G2072), .Z(new_n805));
  NOR2_X1   g380(.A1(G4), .A2(G16), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n624), .B2(G16), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT89), .B(G1348), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n789), .A2(new_n805), .A3(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(G1956), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n702), .A2(G20), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT23), .ZN(new_n813));
  INV_X1    g388(.A(G299), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(new_n702), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT93), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n811), .A2(new_n816), .B1(new_n770), .B2(G2090), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n811), .B2(new_n816), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT94), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n729), .A2(G27), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G164), .B2(new_n729), .ZN(new_n821));
  INV_X1    g396(.A(G2078), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n821), .B(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n557), .A2(new_n702), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n702), .B2(G19), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1341), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n810), .A2(new_n819), .A3(new_n823), .A4(new_n826), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n743), .A2(new_n827), .ZN(G311));
  INV_X1    g403(.A(G311), .ZN(G150));
  AND2_X1   g404(.A1(new_n537), .A2(G55), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n831));
  INV_X1    g406(.A(G93), .ZN(new_n832));
  OAI22_X1  g407(.A1(new_n831), .A2(new_n517), .B1(new_n832), .B2(new_n528), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n835), .A2(new_n555), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n555), .B(KEYINPUT71), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n836), .B1(new_n837), .B2(new_n835), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT38), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n624), .A2(G559), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n842));
  INV_X1    g417(.A(G860), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n834), .A2(new_n843), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT37), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(G145));
  XNOR2_X1  g423(.A(G160), .B(new_n483), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT95), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n648), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n499), .A2(new_n503), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n491), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n748), .B(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n780), .ZN(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT96), .Z(new_n858));
  OR3_X1    g433(.A1(new_n858), .A2(KEYINPUT97), .A3(new_n802), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n802), .ZN(new_n860));
  INV_X1    g435(.A(new_n857), .ZN(new_n861));
  OAI21_X1  g436(.A(KEYINPUT97), .B1(new_n861), .B2(new_n801), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n859), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n735), .B(new_n639), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n479), .A2(G142), .ZN(new_n865));
  OR2_X1    g440(.A1(G106), .A2(G2105), .ZN(new_n866));
  OAI211_X1 g441(.A(new_n866), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n867));
  INV_X1    g442(.A(G130), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n865), .B(new_n867), .C1(new_n868), .C2(new_n476), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n864), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT98), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n852), .B1(new_n863), .B2(new_n872), .ZN(new_n873));
  OAI211_X1 g448(.A(new_n859), .B(new_n870), .C1(new_n860), .C2(new_n862), .ZN(new_n874));
  AOI21_X1  g449(.A(G37), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n863), .B(new_n872), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n876), .A2(KEYINPUT99), .A3(new_n852), .ZN(new_n877));
  AOI21_X1  g452(.A(KEYINPUT99), .B1(new_n876), .B2(new_n852), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g455(.A1(new_n835), .A2(new_n627), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n633), .B(new_n838), .Z(new_n882));
  NAND2_X1  g457(.A1(new_n620), .A2(new_n623), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n814), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT100), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n624), .A2(G299), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n882), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT101), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n886), .B(new_n887), .Z(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT41), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT41), .B1(new_n887), .B2(new_n884), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT102), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n890), .B1(new_n882), .B2(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(G290), .B(KEYINPUT103), .Z(new_n898));
  NAND2_X1  g473(.A1(new_n713), .A2(new_n715), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n898), .B(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(G166), .B(new_n603), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n900), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(new_n903), .B2(new_n900), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n906), .A2(KEYINPUT42), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n906), .B(KEYINPUT105), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n907), .B1(new_n908), .B2(KEYINPUT42), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n897), .B(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n881), .B1(new_n910), .B2(new_n627), .ZN(G295));
  OAI21_X1  g486(.A(new_n881), .B1(new_n910), .B2(new_n627), .ZN(G331));
  NAND2_X1  g487(.A1(G286), .A2(G171), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT107), .ZN(new_n914));
  NAND2_X1  g489(.A1(G301), .A2(G168), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(KEYINPUT106), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(new_n838), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n891), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT109), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n887), .A2(new_n884), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT41), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n918), .B(new_n922), .C1(new_n888), .C2(KEYINPUT41), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n926), .B1(new_n891), .B2(new_n918), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n920), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n923), .A2(new_n924), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n908), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n919), .B1(new_n895), .B2(new_n918), .ZN(new_n931));
  INV_X1    g506(.A(new_n908), .ZN(new_n932));
  AOI21_X1  g507(.A(G37), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n930), .A2(new_n933), .A3(KEYINPUT43), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n931), .A2(new_n932), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT43), .B1(new_n935), .B2(new_n933), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT44), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n930), .A2(new_n933), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n938), .B1(new_n935), .B2(new_n933), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n937), .B1(new_n941), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g517(.A(G1384), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n855), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT110), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT45), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(G1384), .B1(new_n491), .B2(new_n854), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT110), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n467), .ZN(new_n950));
  OAI21_X1  g525(.A(G2105), .B1(new_n465), .B2(new_n950), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n951), .A2(G40), .A3(new_n473), .A4(new_n470), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n748), .B(new_n753), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n954), .B1(new_n780), .B2(new_n955), .ZN(new_n956));
  XOR2_X1   g531(.A(new_n956), .B(KEYINPUT126), .Z(new_n957));
  INV_X1    g532(.A(G1996), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n953), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT46), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT125), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n960), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n957), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT47), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n780), .B(G1996), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n954), .B1(new_n955), .B2(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n967), .B(KEYINPUT111), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n968), .A2(new_n738), .A3(new_n736), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(G2067), .B2(new_n748), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n953), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n735), .B(new_n738), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n968), .B1(new_n954), .B2(new_n972), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n954), .A2(G1986), .A3(G290), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT48), .ZN(new_n975));
  OAI211_X1 g550(.A(new_n965), .B(new_n971), .C1(new_n973), .C2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n952), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n853), .B1(new_n488), .B2(new_n490), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(G1384), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n978), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n510), .A2(KEYINPUT67), .A3(new_n491), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT67), .B1(new_n510), .B2(new_n491), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n985), .A2(new_n986), .A3(G1384), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n984), .B1(new_n987), .B2(KEYINPUT45), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n855), .A2(new_n989), .A3(new_n943), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n978), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n507), .A2(new_n943), .A3(new_n511), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n991), .B1(new_n992), .B2(KEYINPUT50), .ZN(new_n993));
  INV_X1    g568(.A(G2090), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n988), .A2(new_n706), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G8), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n532), .A2(G8), .A3(new_n533), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n997), .B(KEYINPUT55), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n995), .A2(new_n996), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1981), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n596), .A2(KEYINPUT77), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n536), .A2(new_n594), .A3(G48), .ZN(new_n1002));
  OAI22_X1  g577(.A1(new_n575), .A2(new_n589), .B1(new_n591), .B2(new_n535), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n1001), .A2(new_n1002), .B1(new_n1003), .B2(G651), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n552), .A2(G86), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1000), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1006), .B1(new_n603), .B2(new_n1000), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT49), .B1(new_n1007), .B2(KEYINPUT113), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT49), .ZN(new_n1010));
  AOI211_X1 g585(.A(G1981), .B(new_n598), .C1(new_n601), .C2(new_n602), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1009), .B(new_n1010), .C1(new_n1011), .C2(new_n1006), .ZN(new_n1012));
  NOR3_X1   g587(.A1(new_n952), .A2(new_n979), .A3(G1384), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT112), .B1(new_n1013), .B2(new_n996), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n978), .A2(new_n947), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1015), .A2(new_n1016), .A3(G8), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1008), .A2(new_n1012), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1976), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(G288), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n713), .A2(G1976), .A3(new_n715), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n1018), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1016), .B1(new_n1015), .B2(G8), .ZN(new_n1024));
  AOI211_X1 g599(.A(KEYINPUT112), .B(new_n996), .C1(new_n978), .C2(new_n947), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1022), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(KEYINPUT52), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1019), .A2(new_n1023), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n997), .B(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n983), .B1(new_n992), .B2(new_n980), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n507), .A2(new_n989), .A3(new_n943), .A4(new_n511), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n952), .B1(new_n944), .B2(KEYINPUT50), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI22_X1  g609(.A1(new_n1031), .A2(G1971), .B1(new_n1034), .B2(G2090), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1030), .B1(new_n1035), .B2(G8), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n999), .A2(new_n1028), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT51), .ZN(new_n1038));
  INV_X1    g613(.A(G2084), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n993), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n507), .A2(new_n511), .A3(new_n981), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n952), .B1(new_n944), .B2(new_n980), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1966), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1040), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1038), .B(G8), .C1(new_n1046), .C2(G286), .ZN(new_n1047));
  NOR2_X1   g622(.A1(G168), .A2(new_n996), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n993), .A2(new_n1039), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT51), .B(new_n1049), .C1(new_n1050), .C2(new_n996), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT121), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1050), .A2(KEYINPUT121), .A3(new_n1049), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1047), .B(new_n1051), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT53), .B1(new_n1031), .B2(new_n822), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n993), .A2(G1961), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT122), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1059), .B1(new_n1043), .B2(G2078), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1041), .A2(new_n1042), .A3(KEYINPUT122), .A4(new_n822), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(KEYINPUT53), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1058), .A2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(G301), .B(KEYINPUT54), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n984), .A2(KEYINPUT53), .A3(new_n822), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1064), .B1(new_n949), .B2(new_n1065), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1063), .A2(new_n1064), .B1(new_n1058), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1037), .A2(new_n1055), .A3(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT56), .B(G2072), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1031), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n1071));
  AND3_X1   g646(.A1(G299), .A2(new_n1071), .A3(KEYINPUT57), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT57), .B1(G299), .B2(new_n1071), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1034), .A2(new_n811), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1070), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT119), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1073), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n1079));
  NAND3_X1  g654(.A1(G299), .A2(new_n1071), .A3(KEYINPUT57), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT117), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1082));
  AOI21_X1  g657(.A(G1956), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1069), .ZN(new_n1084));
  AOI211_X1 g659(.A(new_n1084), .B(new_n983), .C1(new_n992), .C2(new_n980), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1081), .B(new_n1082), .C1(new_n1083), .C2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1070), .A2(new_n1074), .A3(new_n1075), .A4(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1077), .A2(new_n1086), .A3(KEYINPUT61), .A4(new_n1088), .ZN(new_n1089));
  OAI22_X1  g664(.A1(new_n1085), .A2(new_n1083), .B1(new_n1073), .B2(new_n1072), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n1076), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT61), .ZN(new_n1092));
  XNOR2_X1  g667(.A(KEYINPUT58), .B(G1341), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1013), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1094), .B1(new_n1031), .B2(new_n958), .ZN(new_n1095));
  OAI211_X1 g670(.A(KEYINPUT118), .B(KEYINPUT59), .C1(new_n1095), .C2(new_n837), .ZN(new_n1096));
  NAND2_X1  g671(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1097));
  AOI211_X1 g672(.A(G1996), .B(new_n983), .C1(new_n992), .C2(new_n980), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n557), .B(new_n1097), .C1(new_n1098), .C2(new_n1094), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1091), .A2(new_n1092), .B1(new_n1096), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1013), .A2(new_n753), .ZN(new_n1101));
  OAI211_X1 g676(.A(KEYINPUT60), .B(new_n1101), .C1(new_n993), .C2(G1348), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n624), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(new_n883), .A3(new_n1103), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1104), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OR2_X1    g683(.A1(new_n993), .A2(G1348), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT60), .B1(new_n1109), .B2(new_n1101), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1089), .B(new_n1100), .C1(new_n1108), .C2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1101), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n624), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n1086), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n1076), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1068), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1019), .A2(new_n1023), .A3(new_n1027), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1035), .A2(G8), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n998), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n993), .A2(new_n994), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1031), .A2(G1971), .ZN(new_n1121));
  OAI211_X1 g696(.A(G8), .B(new_n1030), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1050), .A2(new_n996), .A3(G286), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1117), .A2(new_n1119), .A3(new_n1122), .A4(new_n1123), .ZN(new_n1124));
  XOR2_X1   g699(.A(KEYINPUT114), .B(KEYINPUT63), .Z(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n999), .A2(new_n1028), .ZN(new_n1127));
  OAI21_X1  g702(.A(KEYINPUT115), .B1(new_n995), .B2(new_n996), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT115), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1129), .B(G8), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1128), .A2(new_n998), .A3(new_n1130), .ZN(new_n1131));
  AND4_X1   g706(.A1(KEYINPUT63), .A2(new_n1046), .A3(G8), .A4(G168), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1127), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1126), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1117), .A2(new_n999), .ZN(new_n1135));
  AOI211_X1 g710(.A(G1976), .B(G288), .C1(new_n1008), .C2(new_n1012), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1018), .B1(new_n1136), .B2(new_n1011), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1134), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT123), .B1(new_n1116), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1138), .B1(new_n1126), .B2(new_n1133), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1114), .A2(new_n1076), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1089), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1110), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1107), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n883), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1148), .B1(new_n1151), .B2(new_n1104), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1144), .B1(new_n1147), .B2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1142), .B(new_n1143), .C1(new_n1153), .C2(new_n1068), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1037), .A2(G171), .A3(new_n1063), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n1055), .A2(KEYINPUT62), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1055), .A2(KEYINPUT62), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1141), .A2(new_n1154), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n1160));
  XNOR2_X1  g735(.A(G290), .B(G1986), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n973), .B1(new_n953), .B2(new_n1161), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1159), .A2(new_n1160), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1160), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n977), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(KEYINPUT127), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1167), .B(new_n977), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1166), .A2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g744(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1171));
  OAI211_X1 g745(.A(new_n879), .B(new_n1171), .C1(new_n939), .C2(new_n940), .ZN(G225));
  INV_X1    g746(.A(G225), .ZN(G308));
endmodule


