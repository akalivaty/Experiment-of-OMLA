//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 0 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n559, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n595,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1160,
    new_n1161, new_n1162, new_n1163;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT64), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT66), .Z(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n454), .A2(new_n459), .B1(new_n448), .B2(new_n455), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT67), .Z(G319));
  INV_X1    g036(.A(KEYINPUT69), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G137), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n462), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND4_X1  g046(.A1(new_n467), .A2(KEYINPUT69), .A3(G137), .A4(new_n468), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n468), .A2(G101), .A3(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n465), .A2(new_n466), .ZN(new_n476));
  INV_X1    g051(.A(G125), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(KEYINPUT68), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT68), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n478), .A2(new_n481), .A3(G2105), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n474), .B1(new_n480), .B2(new_n482), .ZN(G160));
  NOR2_X1   g058(.A1(new_n476), .A2(new_n468), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  AND2_X1   g060(.A1(G112), .A2(G2105), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n486), .B1(G100), .B2(new_n468), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n485), .B1(new_n464), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n469), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(G136), .B2(new_n489), .ZN(G162));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n491), .B1(new_n469), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G126), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n465), .B2(new_n466), .ZN(new_n495));
  AND2_X1   g070(.A1(G114), .A2(G2104), .ZN(new_n496));
  OAI21_X1  g071(.A(G2105), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT4), .A2(G138), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n465), .B2(new_n466), .ZN(new_n499));
  AND2_X1   g074(.A1(G102), .A2(G2104), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n468), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n493), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  OAI211_X1 g080(.A(KEYINPUT70), .B(new_n504), .C1(new_n505), .C2(KEYINPUT71), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT70), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(G543), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT5), .B1(new_n505), .B2(KEYINPUT70), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT6), .B(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G88), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G50), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n516), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n514), .A2(new_n520), .ZN(G166));
  NAND2_X1  g096(.A1(new_n511), .A2(KEYINPUT72), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n523));
  OAI211_X1 g098(.A(new_n523), .B(new_n506), .C1(new_n509), .C2(new_n510), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n525), .A2(G63), .A3(G651), .ZN(new_n526));
  INV_X1    g101(.A(new_n518), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  INV_X1    g105(.A(G89), .ZN(new_n531));
  OAI211_X1 g106(.A(new_n528), .B(new_n530), .C1(new_n516), .C2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n526), .A2(new_n532), .ZN(G168));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(new_n524), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n504), .B1(new_n507), .B2(G543), .ZN(new_n536));
  OAI21_X1  g111(.A(KEYINPUT70), .B1(new_n505), .B2(KEYINPUT71), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n523), .B1(new_n538), .B2(new_n506), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G64), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n534), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G651), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n511), .A2(new_n515), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n544), .A2(G90), .B1(G52), .B2(new_n527), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n543), .A2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  INV_X1    g123(.A(G43), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n516), .A2(new_n548), .B1(new_n518), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  INV_X1    g126(.A(G68), .ZN(new_n552));
  OAI22_X1  g127(.A1(new_n540), .A2(new_n551), .B1(new_n552), .B2(new_n505), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n513), .B1(new_n553), .B2(KEYINPUT73), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n555));
  OAI221_X1 g130(.A(new_n555), .B1(new_n552), .B2(new_n505), .C1(new_n540), .C2(new_n551), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n550), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G188));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OR3_X1    g139(.A1(new_n518), .A2(KEYINPUT9), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT9), .B1(new_n518), .B2(new_n564), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n565), .A2(new_n566), .B1(new_n544), .B2(G91), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n511), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(new_n513), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(G299));
  INV_X1    g145(.A(G168), .ZN(G286));
  INV_X1    g146(.A(G166), .ZN(G303));
  OAI21_X1  g147(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n544), .A2(G87), .B1(G49), .B2(new_n527), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT74), .ZN(G288));
  AOI22_X1  g151(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(new_n513), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n544), .A2(G86), .B1(G48), .B2(new_n527), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(G305));
  AOI22_X1  g155(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n581), .A2(new_n513), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n544), .A2(G85), .B1(G47), .B2(new_n527), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(new_n544), .A2(G92), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT10), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n585), .B(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n513), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(G54), .B2(new_n527), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  MUX2_X1   g166(.A(new_n591), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g167(.A(new_n591), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g168(.A1(G286), .A2(G868), .ZN(new_n594));
  XOR2_X1   g169(.A(G299), .B(KEYINPUT75), .Z(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(G868), .ZN(G280));
  XNOR2_X1  g171(.A(G280), .B(KEYINPUT76), .ZN(G297));
  AND2_X1   g172(.A1(new_n587), .A2(new_n590), .ZN(new_n598));
  INV_X1    g173(.A(G559), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(G860), .ZN(G148));
  NAND2_X1  g175(.A1(new_n598), .A2(new_n599), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G868), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT77), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n489), .A2(G2104), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT12), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT13), .ZN(new_n608));
  INV_X1    g183(.A(G2100), .ZN(new_n609));
  OR2_X1    g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n484), .A2(G123), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT78), .ZN(new_n612));
  MUX2_X1   g187(.A(G99), .B(G111), .S(G2105), .Z(new_n613));
  AOI22_X1  g188(.A1(new_n489), .A2(G135), .B1(G2104), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT79), .B(G2096), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n608), .A2(new_n609), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n610), .A2(new_n617), .A3(new_n618), .ZN(G156));
  XOR2_X1   g194(.A(G2443), .B(G2446), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT81), .ZN(new_n621));
  XNOR2_X1  g196(.A(G2451), .B(G2454), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT14), .ZN(new_n626));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2435), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT82), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2427), .B(G2430), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n626), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n629), .B2(new_n630), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n625), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G1341), .B(G1348), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT83), .Z(new_n636));
  INV_X1    g211(.A(G14), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n633), .B2(new_n634), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(G401));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  NOR3_X1   g220(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT18), .ZN(new_n647));
  INV_X1    g222(.A(new_n643), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(KEYINPUT17), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n644), .B1(new_n650), .B2(new_n641), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n651), .B1(new_n642), .B2(new_n649), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n642), .A2(new_n645), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n648), .B1(new_n653), .B2(KEYINPUT17), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n647), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2096), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(new_n609), .ZN(G227));
  XOR2_X1   g232(.A(G1961), .B(G1966), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT84), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1956), .B(G2474), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1971), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT20), .Z(new_n666));
  NOR2_X1   g241(.A1(new_n659), .A2(new_n661), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n668), .A2(new_n664), .A3(new_n662), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n666), .B(new_n669), .C1(new_n664), .C2(new_n668), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT85), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n670), .B(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(G1991), .B(G1996), .Z(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(G229));
  MUX2_X1   g252(.A(G23), .B(new_n575), .S(G16), .Z(new_n678));
  XOR2_X1   g253(.A(KEYINPUT33), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  MUX2_X1   g255(.A(G6), .B(G305), .S(G16), .Z(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT32), .B(G1981), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(G16), .A2(G22), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(G166), .B2(G16), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT87), .B(G1971), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n680), .A2(new_n683), .A3(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(KEYINPUT34), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(G25), .A2(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n484), .A2(G119), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n489), .A2(G131), .ZN(new_n693));
  MUX2_X1   g268(.A(G95), .B(G107), .S(G2105), .Z(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G2104), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n691), .B1(new_n697), .B2(G29), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT35), .B(G1991), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(G16), .A2(G24), .ZN(new_n701));
  INV_X1    g276(.A(G290), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(G16), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT86), .B(G1986), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n690), .A2(new_n700), .A3(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n688), .A2(new_n689), .ZN(new_n707));
  OAI22_X1  g282(.A1(new_n706), .A2(new_n707), .B1(KEYINPUT88), .B2(KEYINPUT36), .ZN(new_n708));
  NAND2_X1  g283(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n708), .B(new_n709), .Z(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT31), .B(G11), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT94), .B(G28), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n712), .A2(KEYINPUT30), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(KEYINPUT30), .ZN(new_n714));
  INV_X1    g289(.A(G29), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OAI221_X1 g291(.A(new_n711), .B1(new_n713), .B2(new_n716), .C1(new_n615), .C2(new_n715), .ZN(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NOR2_X1   g293(.A1(G168), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n718), .B2(G21), .ZN(new_n720));
  INV_X1    g295(.A(G1966), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(G29), .A2(G35), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G162), .B2(G29), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT29), .Z(new_n725));
  INV_X1    g300(.A(G2090), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT98), .ZN(new_n728));
  AOI211_X1 g303(.A(new_n717), .B(new_n722), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT24), .B(G34), .Z(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(G29), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G160), .B2(G29), .ZN(new_n732));
  AOI21_X1  g307(.A(KEYINPUT92), .B1(new_n732), .B2(G2084), .ZN(new_n733));
  INV_X1    g308(.A(new_n727), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(KEYINPUT98), .ZN(new_n735));
  NAND3_X1  g310(.A1(new_n732), .A2(KEYINPUT92), .A3(G2084), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n484), .A2(G129), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n489), .A2(G141), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT26), .Z(new_n741));
  NAND4_X1  g316(.A1(new_n737), .A2(new_n738), .A3(new_n739), .A4(new_n741), .ZN(new_n742));
  MUX2_X1   g317(.A(G32), .B(new_n742), .S(G29), .Z(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT93), .Z(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT27), .B(G1996), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OAI22_X1  g321(.A1(new_n725), .A2(new_n726), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n718), .A2(G20), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT99), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT23), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G299), .B2(G16), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT100), .B(G1956), .Z(new_n752));
  OAI22_X1  g327(.A1(new_n720), .A2(new_n721), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n747), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n729), .A2(new_n735), .A3(new_n736), .A4(new_n754), .ZN(new_n755));
  NOR2_X1   g330(.A1(G27), .A2(G29), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G164), .B2(G29), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT97), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT96), .B(G2078), .Z(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n715), .A2(G33), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(KEYINPUT25), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(KEYINPUT25), .ZN(new_n764));
  INV_X1    g339(.A(G139), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n763), .B(new_n764), .C1(new_n469), .C2(new_n765), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT91), .Z(new_n767));
  AOI22_X1  g342(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n767), .B1(G2105), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n761), .B1(new_n770), .B2(new_n715), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n771), .A2(G2072), .B1(new_n751), .B2(new_n752), .ZN(new_n772));
  INV_X1    g347(.A(G1961), .ZN(new_n773));
  NOR2_X1   g348(.A1(G171), .A2(new_n718), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G5), .B2(new_n718), .ZN(new_n775));
  OAI221_X1 g350(.A(new_n772), .B1(G2072), .B2(new_n771), .C1(new_n773), .C2(new_n775), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n755), .A2(new_n760), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n715), .A2(G26), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT28), .Z(new_n779));
  MUX2_X1   g354(.A(G104), .B(G116), .S(G2105), .Z(new_n780));
  AOI22_X1  g355(.A1(new_n484), .A2(G128), .B1(G2104), .B2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(G140), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(new_n469), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n779), .B1(new_n783), .B2(G29), .ZN(new_n784));
  XOR2_X1   g359(.A(KEYINPUT89), .B(G2067), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(G4), .A2(G16), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n598), .B2(G16), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G1348), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n786), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(G16), .A2(G19), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n557), .B2(G16), .ZN(new_n793));
  INV_X1    g368(.A(G1341), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  OAI221_X1 g371(.A(new_n791), .B1(new_n790), .B2(new_n789), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT90), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n744), .A2(new_n746), .ZN(new_n801));
  INV_X1    g376(.A(new_n775), .ZN(new_n802));
  OAI221_X1 g377(.A(new_n801), .B1(G2084), .B2(new_n732), .C1(new_n802), .C2(G1961), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT95), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n777), .A2(new_n799), .A3(new_n800), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n710), .A2(new_n805), .ZN(G311));
  INV_X1    g381(.A(G311), .ZN(G150));
  NAND2_X1  g382(.A1(new_n598), .A2(G559), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT38), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n544), .A2(G93), .B1(G55), .B2(new_n527), .ZN(new_n810));
  OAI21_X1  g385(.A(G67), .B1(new_n535), .B2(new_n539), .ZN(new_n811));
  NAND2_X1  g386(.A1(G80), .A2(G543), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(KEYINPUT101), .B1(new_n813), .B2(G651), .ZN(new_n814));
  INV_X1    g389(.A(G67), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n522), .B2(new_n524), .ZN(new_n816));
  INV_X1    g391(.A(new_n812), .ZN(new_n817));
  OAI211_X1 g392(.A(KEYINPUT101), .B(G651), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n810), .B1(new_n814), .B2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT102), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n554), .A2(new_n556), .ZN(new_n823));
  INV_X1    g398(.A(new_n550), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n810), .ZN(new_n826));
  OAI21_X1  g401(.A(G651), .B1(new_n816), .B2(new_n817), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT101), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n826), .B1(new_n829), .B2(new_n818), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT102), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n822), .A2(new_n825), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n557), .A2(new_n820), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n809), .B(new_n834), .Z(new_n835));
  INV_X1    g410(.A(KEYINPUT39), .ZN(new_n836));
  AOI21_X1  g411(.A(G860), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n836), .B2(new_n835), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n822), .A2(new_n831), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G860), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT103), .B(KEYINPUT37), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n838), .A2(new_n842), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT104), .Z(G145));
  XNOR2_X1  g419(.A(new_n607), .B(new_n696), .ZN(new_n845));
  MUX2_X1   g420(.A(G106), .B(G118), .S(G2105), .Z(new_n846));
  AOI22_X1  g421(.A1(new_n484), .A2(G130), .B1(G2104), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(G142), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(new_n848), .B2(new_n469), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n845), .B(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n850), .A2(KEYINPUT107), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n783), .B(new_n502), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n742), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT105), .Z(new_n854));
  NAND3_X1  g429(.A1(new_n854), .A2(KEYINPUT106), .A3(new_n770), .ZN(new_n855));
  INV_X1    g430(.A(new_n770), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n850), .A2(KEYINPUT107), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(KEYINPUT106), .B1(new_n854), .B2(new_n770), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n851), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n859), .ZN(new_n861));
  INV_X1    g436(.A(new_n851), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n861), .A2(new_n855), .A3(new_n857), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(G162), .B(G160), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n615), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(G37), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n860), .A2(new_n863), .A3(new_n866), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n868), .A2(KEYINPUT40), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT40), .B1(new_n868), .B2(new_n869), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(G395));
  NOR2_X1   g447(.A1(new_n839), .A2(G868), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n834), .B(new_n601), .ZN(new_n874));
  INV_X1    g449(.A(G299), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n598), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n591), .A2(G299), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n876), .A2(KEYINPUT41), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT41), .B1(new_n876), .B2(new_n877), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n874), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n876), .A2(new_n877), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n882), .B1(new_n874), .B2(new_n883), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n884), .A2(KEYINPUT42), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(KEYINPUT42), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(G290), .B(new_n575), .ZN(new_n888));
  XNOR2_X1  g463(.A(G303), .B(G305), .ZN(new_n889));
  XOR2_X1   g464(.A(new_n888), .B(new_n889), .Z(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n885), .A2(new_n890), .A3(new_n886), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n873), .B1(new_n894), .B2(G868), .ZN(G295));
  AOI21_X1  g470(.A(new_n873), .B1(new_n894), .B2(G868), .ZN(G331));
  XNOR2_X1  g471(.A(G301), .B(G286), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n832), .A2(new_n833), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n897), .B1(new_n832), .B2(new_n833), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n881), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT108), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n897), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n830), .A2(KEYINPUT102), .ZN(new_n904));
  AOI211_X1 g479(.A(new_n821), .B(new_n826), .C1(new_n829), .C2(new_n818), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n904), .A2(new_n905), .A3(new_n557), .ZN(new_n906));
  INV_X1    g481(.A(new_n833), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n832), .A2(new_n897), .A3(new_n833), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n908), .A2(new_n877), .A3(new_n876), .A4(new_n909), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n881), .B(KEYINPUT108), .C1(new_n898), .C2(new_n899), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n902), .A2(new_n891), .A3(new_n910), .A4(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(G37), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n900), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(new_n890), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n912), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT41), .ZN(new_n918));
  INV_X1    g493(.A(new_n877), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n591), .A2(G299), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n878), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n922), .B1(new_n908), .B2(new_n909), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n910), .B1(new_n923), .B2(KEYINPUT108), .ZN(new_n924));
  INV_X1    g499(.A(new_n911), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n890), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n926), .A2(new_n927), .A3(new_n913), .A4(new_n912), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n917), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT44), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n916), .A2(new_n927), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n926), .A2(KEYINPUT43), .A3(new_n913), .A4(new_n912), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT44), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n930), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n934), .B1(new_n917), .B2(new_n928), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT44), .B1(new_n931), .B2(new_n932), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT109), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(G397));
  INV_X1    g516(.A(KEYINPUT120), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT113), .ZN(new_n943));
  INV_X1    g518(.A(G8), .ZN(new_n944));
  NOR2_X1   g519(.A1(G166), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT55), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n945), .A2(KEYINPUT55), .ZN(new_n949));
  MUX2_X1   g524(.A(new_n943), .B(new_n948), .S(new_n949), .Z(new_n950));
  INV_X1    g525(.A(G1384), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n502), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n502), .A2(KEYINPUT45), .A3(new_n951), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AND2_X1   g531(.A1(G160), .A2(G40), .ZN(new_n957));
  AOI21_X1  g532(.A(G1971), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(G160), .A2(G40), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n952), .A2(KEYINPUT112), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n502), .A2(new_n961), .A3(new_n951), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(KEYINPUT50), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT50), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n952), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n959), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n958), .B1(new_n726), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n950), .B1(new_n967), .B2(new_n944), .ZN(new_n968));
  INV_X1    g543(.A(new_n958), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n502), .A2(new_n961), .A3(new_n951), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n961), .B1(new_n502), .B2(new_n951), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n964), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n502), .A2(KEYINPUT50), .A3(new_n951), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n959), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(new_n726), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n944), .B1(new_n969), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n949), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT113), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n978), .B1(new_n948), .B2(new_n977), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n976), .A2(new_n979), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n960), .A2(G160), .A3(G40), .A4(new_n962), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n982));
  INV_X1    g557(.A(G1976), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n982), .B1(new_n575), .B2(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n573), .A2(KEYINPUT114), .A3(new_n574), .A4(G1976), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n981), .A2(new_n984), .A3(G8), .A4(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT115), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n986), .A2(new_n990), .A3(KEYINPUT52), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT52), .B1(G288), .B2(new_n983), .ZN(new_n993));
  INV_X1    g568(.A(G1981), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n994), .B1(new_n578), .B2(new_n579), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n578), .A2(new_n579), .A3(new_n994), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT49), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n997), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT49), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n999), .A2(new_n1000), .A3(new_n995), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n981), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1003), .A2(new_n944), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n987), .A2(new_n993), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1005));
  AND4_X1   g580(.A1(new_n968), .A2(new_n980), .A3(new_n992), .A4(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT117), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT45), .B1(new_n960), .B2(new_n962), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1007), .B1(new_n1008), .B2(new_n959), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n953), .B1(new_n970), .B2(new_n971), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n957), .A2(new_n1010), .A3(KEYINPUT117), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1009), .A2(new_n955), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(new_n721), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT118), .ZN(new_n1014));
  INV_X1    g589(.A(new_n974), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1014), .B1(new_n1015), .B2(G2084), .ZN(new_n1016));
  INV_X1    g591(.A(G2084), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n974), .A2(KEYINPUT118), .A3(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1013), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(G286), .A2(new_n944), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(KEYINPUT119), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT119), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1006), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT63), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n992), .A2(new_n1005), .ZN(new_n1026));
  INV_X1    g601(.A(new_n976), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1025), .B1(new_n1027), .B2(new_n950), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1026), .A2(new_n1028), .A3(new_n980), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT119), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n1021), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n1024), .A2(new_n1025), .B1(new_n1029), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1004), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1036));
  OR3_X1    g611(.A1(new_n1036), .A2(G1976), .A3(G288), .ZN(new_n1037));
  XOR2_X1   g612(.A(new_n997), .B(KEYINPUT116), .Z(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1035), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  AND4_X1   g615(.A1(new_n979), .A2(new_n992), .A3(new_n976), .A4(new_n1005), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n942), .B1(new_n1034), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT54), .ZN(new_n1045));
  INV_X1    g620(.A(G2078), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n956), .A2(new_n957), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1048), .A2(G2078), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n479), .A2(G40), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n474), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1051), .B1(KEYINPUT125), .B2(new_n1052), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n956), .B(new_n1053), .C1(KEYINPUT125), .C2(new_n1052), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1049), .B(new_n1054), .C1(G1961), .C2(new_n974), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1055), .A2(G171), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1015), .A2(new_n773), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1009), .A2(new_n1011), .A3(new_n955), .A4(new_n1050), .ZN(new_n1058));
  AOI21_X1  g633(.A(G301), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1045), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1045), .B1(new_n1055), .B2(G171), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT126), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1057), .A2(new_n1058), .A3(G301), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1062), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1006), .B(new_n1060), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1013), .A2(new_n1016), .A3(G168), .A4(new_n1018), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1067), .B1(new_n1068), .B2(G8), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1019), .A2(G286), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(KEYINPUT51), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1068), .A2(G8), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1069), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1066), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n956), .A2(new_n957), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT58), .B(G1341), .ZN(new_n1077));
  OAI22_X1  g652(.A1(new_n1076), .A2(G1996), .B1(new_n1003), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n557), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1080));
  XNOR2_X1  g655(.A(new_n1079), .B(new_n1080), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT56), .B(G2072), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n956), .A2(new_n957), .A3(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1083), .B1(new_n966), .B2(G1956), .ZN(new_n1084));
  XNOR2_X1  g659(.A(G299), .B(KEYINPUT57), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1085), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1087), .B(new_n1083), .C1(G1956), .C2(new_n966), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT61), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n1088), .B(KEYINPUT122), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1086), .A2(KEYINPUT61), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1081), .B(new_n1091), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(G2067), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1003), .A2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(new_n1096), .B(KEYINPUT60), .C1(G1348), .C2(new_n974), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1097), .A2(KEYINPUT123), .A3(new_n598), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT123), .B1(new_n1097), .B2(new_n598), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1097), .A2(new_n598), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1096), .B1(new_n974), .B2(G1348), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(KEYINPUT60), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT124), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1104), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1106), .B(new_n1107), .C1(new_n1108), .C2(new_n1098), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1094), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1088), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1102), .A2(new_n598), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1111), .B1(new_n1112), .B2(new_n1086), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1075), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT63), .B1(new_n1033), .B2(new_n1006), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1026), .A2(new_n1028), .A3(new_n980), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1116), .B1(new_n1021), .B2(new_n1032), .ZN(new_n1117));
  OAI211_X1 g692(.A(KEYINPUT120), .B(new_n1042), .C1(new_n1115), .C2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1074), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1072), .B1(KEYINPUT51), .B2(new_n1070), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT62), .B1(new_n1121), .B2(new_n1069), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1120), .A2(new_n1122), .A3(new_n1006), .A4(new_n1059), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1044), .A2(new_n1114), .A3(new_n1118), .A4(new_n1123), .ZN(new_n1124));
  OR3_X1    g699(.A1(new_n959), .A2(KEYINPUT110), .A3(new_n954), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT110), .B1(new_n959), .B2(new_n954), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n783), .B(new_n1095), .ZN(new_n1129));
  INV_X1    g704(.A(G1996), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n742), .B(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(new_n696), .B(new_n699), .Z(new_n1133));
  NOR2_X1   g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(G1986), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n702), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1134), .B1(new_n1137), .B2(KEYINPUT111), .ZN(new_n1138));
  NOR2_X1   g713(.A1(G290), .A2(G1986), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1139), .A2(KEYINPUT111), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1140), .A2(new_n1136), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1128), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1124), .A2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1128), .A2(KEYINPUT48), .A3(new_n1139), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(new_n1127), .B2(new_n1134), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT48), .B1(new_n1128), .B2(new_n1139), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT46), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1129), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1128), .B1(new_n742), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g727(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1152), .B(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n697), .A2(new_n699), .ZN(new_n1155));
  OAI22_X1  g730(.A1(new_n1132), .A2(new_n1155), .B1(G2067), .B2(new_n783), .ZN(new_n1156));
  AOI211_X1 g731(.A(new_n1147), .B(new_n1154), .C1(new_n1128), .C2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1143), .A2(new_n1157), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g733(.A1(G229), .A2(new_n460), .A3(G227), .ZN(new_n1160));
  NAND2_X1  g734(.A1(new_n1160), .A2(new_n639), .ZN(new_n1161));
  AOI21_X1  g735(.A(new_n1161), .B1(new_n868), .B2(new_n869), .ZN(new_n1162));
  INV_X1    g736(.A(new_n933), .ZN(new_n1163));
  AND2_X1   g737(.A1(new_n1162), .A2(new_n1163), .ZN(G308));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(G225));
endmodule


