//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n833, new_n834, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958;
  XOR2_X1   g000(.A(KEYINPUT93), .B(G36gat), .Z(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G29gat), .ZN(new_n203));
  OAI211_X1 g002(.A(KEYINPUT92), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(G29gat), .A2(G36gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT14), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n203), .B(new_n204), .C1(new_n207), .C2(KEYINPUT92), .ZN(new_n208));
  XNOR2_X1  g007(.A(G43gat), .B(G50gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(KEYINPUT15), .A3(new_n209), .ZN(new_n210));
  OR3_X1    g009(.A1(new_n209), .A2(KEYINPUT94), .A3(KEYINPUT15), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT15), .B1(new_n209), .B2(KEYINPUT94), .ZN(new_n212));
  NAND4_X1  g011(.A1(new_n211), .A2(new_n207), .A3(new_n212), .A4(new_n203), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n214), .B(KEYINPUT17), .ZN(new_n215));
  XNOR2_X1  g014(.A(KEYINPUT102), .B(KEYINPUT7), .ZN(new_n216));
  NAND3_X1  g015(.A1(KEYINPUT101), .A2(G85gat), .A3(G92gat), .ZN(new_n217));
  OR2_X1    g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G99gat), .A2(G106gat), .ZN(new_n219));
  INV_X1    g018(.A(G85gat), .ZN(new_n220));
  INV_X1    g019(.A(G92gat), .ZN(new_n221));
  AOI22_X1  g020(.A1(KEYINPUT8), .A2(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n216), .A2(new_n217), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n218), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G99gat), .B(G106gat), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n218), .A2(new_n225), .A3(new_n222), .A4(new_n223), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n215), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n229), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(new_n214), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G134gat), .B(G162gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n235), .B(KEYINPUT103), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n234), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(G190gat), .B(G218gat), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n237), .A2(new_n240), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G231gat), .A2(G233gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(KEYINPUT99), .ZN(new_n245));
  XOR2_X1   g044(.A(KEYINPUT100), .B(G211gat), .Z(new_n246));
  XOR2_X1   g045(.A(new_n245), .B(new_n246), .Z(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(G127gat), .B(G155gat), .Z(new_n249));
  XOR2_X1   g048(.A(G57gat), .B(G64gat), .Z(new_n250));
  NAND2_X1  g049(.A1(G71gat), .A2(G78gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT9), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G71gat), .ZN(new_n254));
  INV_X1    g053(.A(G78gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(new_n251), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n250), .A2(new_n253), .A3(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT98), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n250), .A2(new_n253), .ZN(new_n260));
  INV_X1    g059(.A(new_n251), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT97), .ZN(new_n262));
  OR2_X1    g061(.A1(new_n261), .A2(KEYINPUT97), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n260), .A2(new_n262), .A3(new_n263), .A4(new_n256), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT21), .ZN(new_n266));
  INV_X1    g065(.A(G183gat), .ZN(new_n267));
  XOR2_X1   g066(.A(G15gat), .B(G22gat), .Z(new_n268));
  INV_X1    g067(.A(G1gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT95), .ZN(new_n271));
  AOI21_X1  g070(.A(G8gat), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT16), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n273), .A2(G1gat), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n270), .B1(new_n274), .B2(new_n268), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n272), .B(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n266), .A2(new_n267), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n267), .B1(new_n266), .B2(new_n276), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n249), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n279), .ZN(new_n281));
  INV_X1    g080(.A(new_n249), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n281), .A2(new_n282), .A3(new_n277), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n248), .B1(new_n280), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  OR2_X1    g084(.A1(new_n265), .A2(KEYINPUT21), .ZN(new_n286));
  XNOR2_X1  g085(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n287));
  XOR2_X1   g086(.A(new_n286), .B(new_n287), .Z(new_n288));
  NAND3_X1  g087(.A1(new_n280), .A2(new_n283), .A3(new_n248), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n285), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n288), .ZN(new_n291));
  INV_X1    g090(.A(new_n289), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n291), .B1(new_n292), .B2(new_n284), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G120gat), .B(G148gat), .ZN(new_n295));
  INV_X1    g094(.A(G176gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G204gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n259), .A2(new_n264), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(new_n229), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n259), .A2(new_n264), .A3(new_n227), .A4(new_n228), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G230gat), .A2(G233gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT10), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n301), .A2(new_n306), .A3(new_n302), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n265), .A2(new_n232), .A3(KEYINPUT10), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AOI211_X1 g108(.A(new_n299), .B(new_n305), .C1(new_n304), .C2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT104), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n312), .B1(new_n309), .B2(new_n304), .ZN(new_n313));
  INV_X1    g112(.A(new_n304), .ZN(new_n314));
  AOI211_X1 g113(.A(KEYINPUT104), .B(new_n314), .C1(new_n307), .C2(new_n308), .ZN(new_n315));
  OR2_X1    g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n316), .A2(new_n305), .ZN(new_n317));
  INV_X1    g116(.A(new_n299), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n311), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n243), .A2(new_n294), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT96), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT66), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT25), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT23), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n325), .B1(G169gat), .B2(G176gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(KEYINPUT65), .ZN(new_n327));
  INV_X1    g126(.A(G190gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n267), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n329), .A2(KEYINPUT24), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G169gat), .A2(G176gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(G169gat), .A2(G176gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT23), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT24), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(G183gat), .A3(G190gat), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n331), .A2(new_n332), .A3(new_n334), .A4(new_n336), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n323), .B(new_n324), .C1(new_n327), .C2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT65), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n326), .B(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n330), .A2(KEYINPUT24), .ZN(new_n341));
  NOR2_X1   g140(.A1(G183gat), .A2(G190gat), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n332), .B(new_n336), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n323), .A2(new_n324), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n340), .A2(new_n344), .A3(new_n345), .A4(new_n334), .ZN(new_n346));
  NAND2_X1  g145(.A1(KEYINPUT66), .A2(KEYINPUT25), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n338), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT26), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(new_n332), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT27), .B(G183gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n353), .A2(KEYINPUT28), .A3(new_n328), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT68), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n353), .A2(KEYINPUT68), .A3(KEYINPUT28), .A4(new_n328), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  XOR2_X1   g157(.A(KEYINPUT27), .B(G183gat), .Z(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT67), .ZN(new_n360));
  OR2_X1    g159(.A1(new_n267), .A2(KEYINPUT27), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT67), .ZN(new_n362));
  AOI21_X1  g161(.A(G190gat), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT28), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n330), .B(new_n352), .C1(new_n358), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT1), .ZN(new_n367));
  INV_X1    g166(.A(G113gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(G120gat), .ZN(new_n369));
  INV_X1    g168(.A(G120gat), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n370), .A2(G113gat), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n367), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G134gat), .ZN(new_n373));
  OR2_X1    g172(.A1(KEYINPUT70), .A2(G127gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(KEYINPUT70), .A2(G127gat), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT69), .ZN(new_n377));
  INV_X1    g176(.A(G127gat), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n377), .B1(new_n378), .B2(G134gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n373), .A2(KEYINPUT69), .A3(G127gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n372), .B1(new_n376), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT71), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT71), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n372), .B(new_n384), .C1(new_n376), .C2(new_n381), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n370), .A2(G113gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n368), .A2(G120gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G127gat), .B(G134gat), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n388), .A2(new_n389), .A3(new_n367), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT72), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n388), .A2(new_n389), .A3(KEYINPUT72), .A4(new_n367), .ZN(new_n393));
  AOI22_X1  g192(.A1(new_n383), .A2(new_n385), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n366), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n348), .A2(new_n365), .A3(new_n394), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n399), .B(KEYINPUT64), .Z(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT33), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G15gat), .B(G43gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(G71gat), .B(G99gat), .ZN(new_n404));
  XOR2_X1   g203(.A(new_n403), .B(new_n404), .Z(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n348), .A2(new_n365), .A3(new_n394), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n394), .B1(new_n348), .B2(new_n365), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(KEYINPUT32), .B1(new_n411), .B2(new_n400), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(new_n399), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT34), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n401), .A2(KEYINPUT34), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n412), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n412), .B1(new_n414), .B2(new_n416), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n408), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n414), .A2(new_n416), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT32), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n422), .B1(new_n398), .B2(new_n401), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(new_n407), .A3(new_n417), .ZN(new_n425));
  XOR2_X1   g224(.A(G141gat), .B(G148gat), .Z(new_n426));
  OR2_X1    g225(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n427));
  NAND2_X1  g226(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(G155gat), .ZN(new_n430));
  INV_X1    g229(.A(G162gat), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n431), .A3(KEYINPUT76), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT76), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n433), .B1(G155gat), .B2(G162gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(G155gat), .A2(G162gat), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n429), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(G141gat), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n439), .A2(G148gat), .ZN(new_n440));
  INV_X1    g239(.A(G148gat), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n441), .A2(G141gat), .ZN(new_n442));
  NOR3_X1   g241(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n443));
  INV_X1    g242(.A(new_n435), .ZN(new_n444));
  OAI22_X1  g243(.A1(new_n440), .A2(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n438), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(G197gat), .B(G204gat), .ZN(new_n447));
  INV_X1    g246(.A(G211gat), .ZN(new_n448));
  INV_X1    g247(.A(G218gat), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n447), .B1(KEYINPUT22), .B2(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G211gat), .B(G218gat), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n452), .B(new_n447), .C1(KEYINPUT22), .C2(new_n450), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT29), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n446), .B1(new_n456), .B2(KEYINPUT3), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT81), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n457), .B(new_n458), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n443), .A2(new_n444), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n429), .A2(new_n437), .B1(new_n460), .B2(new_n426), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT78), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT3), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n427), .A2(new_n428), .ZN(new_n465));
  XNOR2_X1  g264(.A(G141gat), .B(G148gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n463), .B(new_n445), .C1(new_n467), .C2(new_n436), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT78), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT29), .B1(new_n464), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(G228gat), .ZN(new_n473));
  INV_X1    g272(.A(G233gat), .ZN(new_n474));
  OAI22_X1  g273(.A1(new_n459), .A2(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n473), .A2(new_n474), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n476), .B(new_n457), .C1(new_n470), .C2(new_n471), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n477), .A2(KEYINPUT82), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(KEYINPUT82), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(G78gat), .B(G106gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(KEYINPUT31), .B(G50gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n483), .A2(G22gat), .ZN(new_n484));
  INV_X1    g283(.A(G22gat), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n485), .A2(KEYINPUT83), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n484), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n480), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n487), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n475), .B(new_n489), .C1(new_n478), .C2(new_n479), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n420), .A2(new_n425), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT89), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n420), .A2(new_n491), .A3(KEYINPUT89), .A4(new_n425), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(G226gat), .A2(G233gat), .ZN(new_n497));
  XOR2_X1   g296(.A(new_n497), .B(KEYINPUT73), .Z(new_n498));
  AND3_X1   g297(.A1(new_n348), .A2(new_n365), .A3(new_n498), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n498), .A2(KEYINPUT29), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n500), .B1(new_n348), .B2(new_n365), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n471), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n471), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n348), .A2(new_n365), .A3(new_n498), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n348), .A2(new_n365), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n503), .B(new_n504), .C1(new_n505), .C2(new_n500), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n502), .A2(new_n506), .A3(KEYINPUT74), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT74), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n508), .B(new_n471), .C1(new_n499), .C2(new_n501), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  XOR2_X1   g309(.A(G8gat), .B(G36gat), .Z(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(G64gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n512), .B(new_n221), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT75), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT30), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n507), .A2(new_n509), .A3(new_n513), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n513), .B1(new_n507), .B2(new_n509), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT30), .B1(new_n520), .B2(KEYINPUT75), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT0), .B(G57gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(G85gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(G1gat), .B(G29gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n392), .A2(new_n393), .ZN(new_n527));
  INV_X1    g326(.A(new_n385), .ZN(new_n528));
  AND2_X1   g327(.A1(KEYINPUT70), .A2(G127gat), .ZN(new_n529));
  NOR2_X1   g328(.A1(KEYINPUT70), .A2(G127gat), .ZN(new_n530));
  OAI21_X1  g329(.A(G134gat), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n531), .A2(new_n379), .A3(new_n380), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n384), .B1(new_n532), .B2(new_n372), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n461), .B(new_n527), .C1(new_n528), .C2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT79), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n383), .A2(new_n385), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n537), .A2(KEYINPUT79), .A3(new_n461), .A4(new_n527), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n536), .B(new_n538), .C1(new_n461), .C2(new_n394), .ZN(new_n539));
  NAND2_X1  g338(.A1(G225gat), .A2(G233gat), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT5), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT4), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT79), .B1(new_n394), .B2(new_n461), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n534), .A2(new_n535), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT80), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n534), .A2(KEYINPUT4), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n536), .A2(new_n538), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT80), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(new_n551), .A3(new_n544), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n548), .A2(new_n549), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n464), .A2(new_n469), .ZN(new_n554));
  OAI211_X1 g353(.A(new_n554), .B(new_n395), .C1(new_n463), .C2(new_n461), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n540), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n543), .B1(new_n553), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n550), .A2(KEYINPUT4), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n534), .A2(new_n544), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n559), .A2(new_n555), .A3(new_n560), .ZN(new_n561));
  OR2_X1    g360(.A1(new_n541), .A2(KEYINPUT5), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n526), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n526), .ZN(new_n565));
  INV_X1    g364(.A(new_n563), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n551), .B1(new_n550), .B2(new_n544), .ZN(new_n567));
  AOI211_X1 g366(.A(KEYINPUT80), .B(KEYINPUT4), .C1(new_n536), .C2(new_n538), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n556), .B1(new_n569), .B2(new_n549), .ZN(new_n570));
  OAI211_X1 g369(.A(new_n565), .B(new_n566), .C1(new_n570), .C2(new_n543), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT6), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n564), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  OAI211_X1 g372(.A(KEYINPUT6), .B(new_n526), .C1(new_n558), .C2(new_n563), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n522), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n496), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(KEYINPUT88), .A2(KEYINPUT35), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n420), .A2(new_n491), .A3(new_n425), .A4(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n526), .B(KEYINPUT84), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(new_n558), .B2(new_n563), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n581), .A2(new_n571), .A3(new_n572), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n578), .B1(new_n574), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(KEYINPUT88), .A2(KEYINPUT35), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n522), .A2(new_n584), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n576), .A2(KEYINPUT35), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT37), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n587), .B1(new_n502), .B2(new_n506), .ZN(new_n588));
  NOR3_X1   g387(.A1(new_n588), .A2(KEYINPUT38), .A3(new_n514), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT86), .B1(new_n510), .B2(new_n587), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT86), .ZN(new_n591));
  AOI211_X1 g390(.A(new_n591), .B(KEYINPUT37), .C1(new_n507), .C2(new_n509), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n589), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n582), .A2(new_n574), .A3(new_n515), .A4(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT87), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n510), .A2(new_n587), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n591), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n510), .A2(KEYINPUT86), .A3(new_n587), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n600), .B1(new_n587), .B2(new_n510), .ZN(new_n601));
  OAI21_X1  g400(.A(KEYINPUT38), .B1(new_n601), .B2(new_n514), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n520), .B1(new_n600), .B2(new_n589), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n603), .A2(KEYINPUT87), .A3(new_n574), .A4(new_n582), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n596), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n491), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n561), .A2(new_n607), .A3(new_n541), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n561), .A2(new_n541), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n539), .A2(new_n541), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n579), .B(new_n608), .C1(new_n611), .C2(new_n607), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT40), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n612), .A2(KEYINPUT85), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n613), .B1(new_n612), .B2(KEYINPUT85), .ZN(new_n615));
  INV_X1    g414(.A(new_n581), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n606), .B1(new_n617), .B2(new_n522), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n605), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT36), .ZN(new_n620));
  INV_X1    g419(.A(new_n420), .ZN(new_n621));
  INV_X1    g420(.A(new_n425), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n620), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n420), .A2(new_n425), .A3(KEYINPUT36), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n625), .B1(new_n575), .B2(new_n491), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n586), .B1(new_n619), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n215), .A2(new_n276), .ZN(new_n629));
  INV_X1    g428(.A(new_n214), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n630), .A2(new_n276), .ZN(new_n631));
  NAND2_X1  g430(.A1(G229gat), .A2(G233gat), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT18), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n630), .B(new_n276), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n632), .B(KEYINPUT13), .Z(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n629), .A2(KEYINPUT18), .A3(new_n631), .A4(new_n632), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n635), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G113gat), .B(G141gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(G169gat), .B(G197gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g442(.A(KEYINPUT90), .B(KEYINPUT11), .Z(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT91), .B(KEYINPUT12), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n640), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n647), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n635), .A2(new_n649), .A3(new_n638), .A4(new_n639), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n322), .B1(new_n628), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n626), .B1(new_n605), .B2(new_n618), .ZN(new_n654));
  OAI211_X1 g453(.A(KEYINPUT96), .B(new_n651), .C1(new_n654), .C2(new_n586), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n321), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n573), .A2(new_n574), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n522), .ZN(new_n660));
  XNOR2_X1  g459(.A(KEYINPUT105), .B(G8gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(new_n273), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n660), .A2(KEYINPUT42), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT42), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n664), .B1(new_n660), .B2(G8gat), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n660), .A2(new_n662), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(G1325gat));
  NOR2_X1   g466(.A1(new_n621), .A2(new_n622), .ZN(new_n668));
  AOI21_X1  g467(.A(G15gat), .B1(new_n656), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n625), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n656), .A2(G15gat), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(G1326gat));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n606), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT43), .B(G22gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n676), .B1(new_n628), .B2(new_n243), .ZN(new_n677));
  INV_X1    g476(.A(new_n243), .ZN(new_n678));
  OAI211_X1 g477(.A(KEYINPUT44), .B(new_n678), .C1(new_n654), .C2(new_n586), .ZN(new_n679));
  INV_X1    g478(.A(new_n294), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n320), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(new_n652), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT106), .ZN(new_n683));
  AND4_X1   g482(.A1(new_n657), .A2(new_n677), .A3(new_n679), .A4(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(G29gat), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT45), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n681), .A2(new_n243), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n688), .B1(new_n653), .B2(new_n655), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(new_n685), .A3(new_n657), .ZN(new_n690));
  MUX2_X1   g489(.A(KEYINPUT45), .B(new_n686), .S(new_n690), .Z(G1328gat));
  INV_X1    g490(.A(KEYINPUT46), .ZN(new_n692));
  INV_X1    g491(.A(new_n202), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n689), .A2(new_n692), .A3(new_n693), .A4(new_n522), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n689), .A2(new_n693), .A3(new_n522), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n677), .A2(new_n522), .A3(new_n679), .A4(new_n683), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n697), .A2(KEYINPUT46), .B1(new_n202), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n694), .A2(new_n695), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n696), .A2(new_n699), .A3(new_n700), .ZN(G1329gat));
  INV_X1    g500(.A(KEYINPUT47), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n677), .A2(new_n670), .A3(new_n679), .A4(new_n683), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(G43gat), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n653), .A2(new_n655), .ZN(new_n705));
  INV_X1    g504(.A(G43gat), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n705), .A2(new_n706), .A3(new_n668), .A4(new_n687), .ZN(new_n707));
  AOI211_X1 g506(.A(KEYINPUT108), .B(new_n702), .C1(new_n704), .C2(new_n707), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n702), .A2(KEYINPUT108), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n702), .A2(KEYINPUT108), .ZN(new_n710));
  AND4_X1   g509(.A1(new_n709), .A2(new_n704), .A3(new_n707), .A4(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n708), .A2(new_n711), .ZN(G1330gat));
  INV_X1    g511(.A(G50gat), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n689), .A2(new_n713), .A3(new_n606), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n677), .A2(new_n606), .A3(new_n679), .A4(new_n683), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(G50gat), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT48), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n715), .A2(KEYINPUT109), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n715), .A2(KEYINPUT109), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n720), .A2(new_n721), .A3(new_n713), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n714), .A2(KEYINPUT48), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n719), .B1(new_n722), .B2(new_n723), .ZN(G1331gat));
  AOI22_X1  g523(.A1(new_n241), .A2(new_n242), .B1(new_n290), .B2(new_n293), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n725), .A2(new_n652), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n319), .B(new_n726), .C1(new_n654), .C2(new_n586), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n657), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(G57gat), .ZN(G1332gat));
  INV_X1    g529(.A(new_n522), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n619), .A2(new_n627), .ZN(new_n732));
  INV_X1    g531(.A(new_n586), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n734), .A2(new_n735), .A3(new_n319), .A4(new_n726), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n727), .A2(KEYINPUT110), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n731), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g539(.A(KEYINPUT49), .B(G64gat), .Z(new_n741));
  AOI211_X1 g540(.A(new_n731), .B(new_n741), .C1(new_n736), .C2(new_n737), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT111), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n741), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n738), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n746));
  OAI211_X1 g545(.A(new_n745), .B(new_n746), .C1(new_n738), .C2(new_n739), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n743), .A2(new_n747), .ZN(G1333gat));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n736), .A2(new_n737), .ZN(new_n750));
  OAI21_X1  g549(.A(G71gat), .B1(new_n750), .B2(new_n625), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n728), .A2(new_n254), .A3(new_n668), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n749), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n625), .B1(new_n736), .B2(new_n737), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n749), .B(new_n752), .C1(new_n754), .C2(new_n254), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n753), .A2(new_n756), .ZN(G1334gat));
  NOR2_X1   g556(.A1(new_n750), .A2(new_n491), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(new_n255), .ZN(G1335gat));
  NOR2_X1   g558(.A1(new_n294), .A2(new_n651), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n734), .A2(KEYINPUT51), .A3(new_n678), .A4(new_n760), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n678), .B(new_n760), .C1(new_n654), .C2(new_n586), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n320), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(G85gat), .B1(new_n765), .B2(new_n657), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n677), .A2(new_n319), .A3(new_n679), .A4(new_n760), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(new_n220), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n766), .B1(new_n657), .B2(new_n768), .ZN(G1336gat));
  OAI21_X1  g568(.A(G92gat), .B1(new_n767), .B2(new_n731), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n761), .A2(new_n764), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n320), .A2(new_n731), .A3(G92gat), .ZN(new_n772));
  OR2_X1    g571(.A1(new_n772), .A2(KEYINPUT112), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(KEYINPUT112), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT52), .ZN(new_n777));
  AOI21_X1  g576(.A(KEYINPUT52), .B1(new_n771), .B2(new_n772), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n770), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1337gat));
  AOI21_X1  g579(.A(G99gat), .B1(new_n765), .B2(new_n668), .ZN(new_n781));
  INV_X1    g580(.A(G99gat), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n767), .A2(new_n782), .A3(new_n625), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n781), .A2(new_n783), .ZN(G1338gat));
  NAND2_X1  g583(.A1(new_n765), .A2(new_n606), .ZN(new_n785));
  INV_X1    g584(.A(G106gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OR3_X1    g586(.A1(new_n767), .A2(new_n786), .A3(new_n491), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(new_n788), .A3(KEYINPUT53), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790));
  AOI21_X1  g589(.A(G106gat), .B1(new_n765), .B2(new_n606), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n767), .A2(new_n786), .A3(new_n491), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n789), .A2(new_n793), .ZN(G1339gat));
  NAND2_X1  g593(.A1(new_n657), .A2(new_n731), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(new_n313), .B2(new_n315), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n309), .A2(new_n304), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n307), .A2(new_n314), .A3(new_n308), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(KEYINPUT54), .A3(new_n799), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n797), .A2(KEYINPUT55), .A3(new_n299), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n311), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT114), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n801), .A2(new_n804), .A3(new_n311), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n797), .A2(new_n299), .A3(new_n800), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n803), .A2(new_n651), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n632), .B1(new_n629), .B2(new_n631), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n636), .A2(new_n637), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n645), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n650), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n319), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n678), .B1(new_n809), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n803), .A2(new_n813), .A3(new_n805), .A4(new_n808), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n243), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n680), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT113), .B1(new_n321), .B2(new_n651), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n725), .A2(new_n820), .A3(new_n652), .A4(new_n320), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n795), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n823), .A2(new_n496), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n824), .A2(new_n368), .A3(new_n651), .ZN(new_n825));
  INV_X1    g624(.A(new_n492), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(G113gat), .B1(new_n827), .B2(new_n652), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n828), .ZN(G1340gat));
  NAND3_X1  g628(.A1(new_n824), .A2(new_n370), .A3(new_n319), .ZN(new_n830));
  OAI21_X1  g629(.A(G120gat), .B1(new_n827), .B2(new_n320), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(G1341gat));
  NAND2_X1  g631(.A1(new_n374), .A2(new_n375), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n827), .A2(new_n833), .A3(new_n680), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n824), .A2(new_n294), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT115), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n834), .B1(new_n836), .B2(new_n833), .ZN(G1342gat));
  NAND3_X1  g636(.A1(new_n824), .A2(new_n373), .A3(new_n678), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT56), .ZN(new_n839));
  OAI21_X1  g638(.A(G134gat), .B1(new_n827), .B2(new_n243), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT56), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n824), .A2(new_n841), .A3(new_n373), .A4(new_n678), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n839), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT116), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n839), .A2(new_n845), .A3(new_n840), .A4(new_n842), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(new_n846), .ZN(G1343gat));
  NOR3_X1   g646(.A1(new_n670), .A2(new_n652), .A3(new_n491), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n823), .A2(new_n439), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n625), .A2(new_n657), .A3(new_n731), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n819), .A2(new_n821), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n651), .A2(new_n808), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n814), .B1(new_n852), .B2(new_n802), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n243), .ZN(new_n854));
  AOI22_X1  g653(.A1(new_n802), .A2(KEYINPUT114), .B1(new_n807), .B2(new_n806), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n678), .A2(new_n855), .A3(new_n813), .A4(new_n805), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n294), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n606), .B1(new_n851), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n850), .B1(new_n858), .B2(KEYINPUT57), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n491), .B1(new_n818), .B2(new_n822), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n859), .A2(new_n651), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n849), .B1(new_n863), .B2(new_n439), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(KEYINPUT58), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(KEYINPUT58), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n849), .B(new_n868), .C1(new_n863), .C2(new_n439), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n867), .A2(new_n869), .ZN(G1344gat));
  INV_X1    g669(.A(new_n850), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n860), .A2(new_n441), .A3(new_n319), .A4(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n818), .A2(new_n822), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n606), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT57), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n321), .B2(new_n651), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n725), .A2(KEYINPUT118), .A3(new_n652), .A4(new_n320), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n861), .B(new_n606), .C1(new_n857), .C2(new_n880), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n876), .A2(new_n319), .A3(new_n871), .A4(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n441), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n881), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n885), .B1(KEYINPUT57), .B2(new_n875), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n886), .A2(KEYINPUT119), .A3(new_n319), .A4(new_n871), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n873), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n859), .A2(new_n862), .ZN(new_n889));
  AOI211_X1 g688(.A(KEYINPUT59), .B(new_n441), .C1(new_n889), .C2(new_n319), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n872), .B1(new_n888), .B2(new_n890), .ZN(G1345gat));
  NAND3_X1  g690(.A1(new_n889), .A2(G155gat), .A3(new_n294), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n860), .A2(new_n871), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n430), .B1(new_n893), .B2(new_n680), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n892), .A2(new_n894), .ZN(G1346gat));
  NAND3_X1  g694(.A1(new_n889), .A2(G162gat), .A3(new_n678), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n431), .B1(new_n893), .B2(new_n243), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(G1347gat));
  NOR2_X1   g697(.A1(new_n657), .A2(new_n731), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n874), .A2(new_n496), .A3(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(G169gat), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(new_n901), .A3(new_n651), .ZN(new_n902));
  INV_X1    g701(.A(new_n899), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n903), .B1(new_n818), .B2(new_n822), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n651), .A3(new_n826), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n905), .A2(KEYINPUT120), .A3(G169gat), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT120), .B1(new_n905), .B2(G169gat), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n902), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT121), .ZN(G1348gat));
  AOI21_X1  g708(.A(G176gat), .B1(new_n900), .B2(new_n319), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n874), .A2(new_n826), .A3(new_n899), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n911), .A2(new_n296), .A3(new_n320), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n910), .A2(new_n912), .ZN(G1349gat));
  INV_X1    g712(.A(KEYINPUT122), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n900), .A2(new_n914), .A3(new_n353), .A4(new_n294), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n904), .A2(new_n353), .A3(new_n496), .A4(new_n294), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT122), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n919), .B1(new_n911), .B2(new_n680), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n904), .A2(KEYINPUT123), .A3(new_n826), .A4(new_n294), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n920), .A2(G183gat), .A3(new_n921), .ZN(new_n922));
  AOI211_X1 g721(.A(KEYINPUT124), .B(KEYINPUT60), .C1(new_n918), .C2(new_n922), .ZN(new_n923));
  OR2_X1    g722(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n924));
  NAND2_X1  g723(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n925));
  AND4_X1   g724(.A1(new_n924), .A2(new_n918), .A3(new_n922), .A4(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n923), .A2(new_n926), .ZN(G1350gat));
  OAI21_X1  g726(.A(G190gat), .B1(new_n911), .B2(new_n243), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n928), .B(KEYINPUT61), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n900), .A2(new_n328), .A3(new_n678), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1351gat));
  NOR2_X1   g730(.A1(new_n903), .A2(new_n670), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n876), .A2(new_n881), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(G197gat), .B1(new_n933), .B2(new_n652), .ZN(new_n934));
  INV_X1    g733(.A(G197gat), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n904), .A2(new_n935), .A3(new_n848), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT125), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(new_n937), .ZN(G1352gat));
  NAND2_X1  g737(.A1(new_n860), .A2(new_n932), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n939), .A2(G204gat), .A3(new_n320), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT62), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n886), .A2(new_n319), .A3(new_n932), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n298), .B2(new_n942), .ZN(G1353gat));
  NAND3_X1  g742(.A1(new_n886), .A2(new_n294), .A3(new_n932), .ZN(new_n944));
  AOI21_X1  g743(.A(KEYINPUT63), .B1(new_n944), .B2(G211gat), .ZN(new_n945));
  OAI211_X1 g744(.A(KEYINPUT63), .B(G211gat), .C1(new_n933), .C2(new_n680), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n294), .A2(new_n448), .ZN(new_n948));
  OAI22_X1  g747(.A1(new_n945), .A2(new_n947), .B1(new_n939), .B2(new_n948), .ZN(G1354gat));
  NAND4_X1  g748(.A1(new_n886), .A2(G218gat), .A3(new_n678), .A4(new_n932), .ZN(new_n950));
  OAI211_X1 g749(.A(KEYINPUT126), .B(new_n449), .C1(new_n939), .C2(new_n243), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n449), .B1(new_n939), .B2(new_n243), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT126), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n950), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT127), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n950), .A2(new_n951), .A3(KEYINPUT127), .A4(new_n954), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1355gat));
endmodule


