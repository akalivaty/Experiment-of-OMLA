//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n938,
    new_n939, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995,
    new_n996;
  AND2_X1   g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G141gat), .B(G148gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT2), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n206), .B1(G155gat), .B2(G162gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G141gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G148gat), .ZN(new_n210));
  INV_X1    g009(.A(G148gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G141gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G155gat), .B(G162gat), .ZN(new_n214));
  INV_X1    g013(.A(G155gat), .ZN(new_n215));
  INV_X1    g014(.A(G162gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT2), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n213), .A2(new_n214), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n208), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT29), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G197gat), .B(G204gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT22), .ZN(new_n224));
  INV_X1    g023(.A(G211gat), .ZN(new_n225));
  INV_X1    g024(.A(G218gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G211gat), .B(G218gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n228), .B(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n230), .A2(KEYINPUT75), .ZN(new_n231));
  INV_X1    g030(.A(new_n229), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n228), .B(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT75), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n222), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(G228gat), .A2(G233gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n219), .B1(new_n230), .B2(KEYINPUT29), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n208), .A2(new_n218), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n236), .A2(new_n237), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT78), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n208), .A2(new_n218), .A3(KEYINPUT78), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n238), .A2(new_n245), .B1(new_n230), .B2(new_n222), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n241), .B1(new_n246), .B2(new_n237), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(G22gat), .ZN(new_n248));
  INV_X1    g047(.A(G22gat), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n241), .B(new_n249), .C1(new_n246), .C2(new_n237), .ZN(new_n250));
  XNOR2_X1  g049(.A(G78gat), .B(G106gat), .ZN(new_n251));
  INV_X1    g050(.A(G50gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n248), .A2(new_n250), .A3(KEYINPUT84), .A4(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n248), .A2(KEYINPUT84), .A3(new_n250), .ZN(new_n257));
  INV_X1    g056(.A(new_n255), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT84), .B1(new_n248), .B2(new_n250), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n235), .A2(new_n231), .ZN(new_n262));
  NAND2_X1  g061(.A1(G226gat), .A2(G233gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(new_n267), .A3(KEYINPUT26), .ZN(new_n268));
  INV_X1    g067(.A(new_n266), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n269), .A2(KEYINPUT69), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT26), .ZN(new_n271));
  INV_X1    g070(.A(G169gat), .ZN(new_n272));
  INV_X1    g071(.A(G176gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n265), .B(new_n268), .C1(new_n270), .C2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT27), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n277), .A2(G183gat), .ZN(new_n278));
  INV_X1    g077(.A(G183gat), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n279), .A2(KEYINPUT27), .ZN(new_n280));
  NOR4_X1   g079(.A1(new_n278), .A2(new_n280), .A3(KEYINPUT28), .A4(G190gat), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT67), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(new_n278), .B2(new_n280), .ZN(new_n283));
  INV_X1    g082(.A(G190gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n279), .A2(KEYINPUT27), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n277), .A2(G183gat), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n285), .A2(new_n286), .A3(KEYINPUT67), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n283), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n281), .B1(new_n288), .B2(KEYINPUT28), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT68), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n276), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  AOI211_X1 g090(.A(KEYINPUT68), .B(new_n281), .C1(new_n288), .C2(KEYINPUT28), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(new_n265), .ZN(new_n294));
  NAND3_X1  g093(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n272), .A2(new_n273), .A3(KEYINPUT23), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT64), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT64), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n266), .A2(new_n300), .A3(KEYINPUT23), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT23), .B1(new_n272), .B2(new_n273), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n299), .A2(new_n301), .B1(new_n269), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT65), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n297), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n269), .ZN(new_n306));
  INV_X1    g105(.A(new_n301), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n300), .B1(new_n266), .B2(KEYINPUT23), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT65), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT25), .B1(new_n305), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n306), .A2(KEYINPUT25), .A3(new_n298), .ZN(new_n312));
  XOR2_X1   g111(.A(new_n295), .B(KEYINPUT66), .Z(new_n313));
  AOI21_X1  g112(.A(new_n312), .B1(new_n313), .B2(new_n294), .ZN(new_n314));
  OAI22_X1  g113(.A1(new_n291), .A2(new_n292), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n264), .B1(new_n315), .B2(new_n221), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n288), .A2(KEYINPUT28), .ZN(new_n317));
  INV_X1    g116(.A(new_n281), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT68), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n289), .A2(new_n290), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(new_n321), .A3(new_n276), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT25), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n296), .B1(new_n309), .B2(KEYINPUT65), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n303), .A2(new_n304), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n314), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n263), .B1(new_n322), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n262), .B1(new_n316), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G8gat), .B(G36gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(G64gat), .B(G92gat), .ZN(new_n332));
  XOR2_X1   g131(.A(new_n331), .B(new_n332), .Z(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n315), .A2(new_n264), .ZN(new_n335));
  AOI21_X1  g134(.A(KEYINPUT29), .B1(new_n322), .B2(new_n328), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n230), .B(new_n335), .C1(new_n336), .C2(new_n264), .ZN(new_n337));
  AND3_X1   g136(.A1(new_n330), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n334), .B1(new_n330), .B2(new_n337), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n338), .B1(KEYINPUT30), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n330), .A2(new_n337), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(new_n333), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT30), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n342), .A2(KEYINPUT76), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n345), .B1(new_n339), .B2(KEYINPUT30), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n340), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n239), .A2(KEYINPUT3), .ZN(new_n348));
  INV_X1    g147(.A(G113gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G120gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT71), .B(G120gat), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n351), .B1(new_n352), .B2(G113gat), .ZN(new_n353));
  INV_X1    g152(.A(G127gat), .ZN(new_n354));
  INV_X1    g153(.A(G134gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G127gat), .A2(G134gat), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT1), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT70), .B(G127gat), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n356), .B1(new_n360), .B2(new_n355), .ZN(new_n361));
  INV_X1    g160(.A(G120gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(G113gat), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT1), .B1(new_n350), .B2(new_n363), .ZN(new_n364));
  OAI22_X1  g163(.A1(new_n353), .A2(new_n359), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n348), .A2(new_n365), .A3(new_n220), .ZN(new_n366));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n367), .B(KEYINPUT77), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  AND2_X1   g168(.A1(new_n366), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT79), .B1(new_n365), .B2(new_n239), .ZN(new_n371));
  INV_X1    g170(.A(new_n364), .ZN(new_n372));
  INV_X1    g171(.A(new_n356), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n354), .A2(KEYINPUT70), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT70), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(G127gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n373), .B1(new_n377), .B2(G134gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n362), .A2(KEYINPUT71), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT71), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G120gat), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n379), .A2(new_n381), .A3(G113gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(new_n350), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n372), .A2(new_n378), .B1(new_n383), .B2(new_n358), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT79), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n208), .A2(new_n218), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n371), .A2(KEYINPUT4), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT4), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n389), .B1(new_n245), .B2(new_n365), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT5), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n370), .A2(new_n388), .A3(new_n390), .A4(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(KEYINPUT4), .B1(new_n371), .B2(new_n387), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n243), .A2(new_n384), .A3(KEYINPUT4), .A4(new_n244), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(new_n369), .A3(new_n366), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT5), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n371), .A2(new_n387), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n365), .A2(new_n239), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n369), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n392), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  XOR2_X1   g199(.A(G1gat), .B(G29gat), .Z(new_n401));
  XNOR2_X1  g200(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G57gat), .B(G85gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n403), .B(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n394), .A2(new_n369), .A3(new_n366), .ZN(new_n407));
  NOR3_X1   g206(.A1(new_n365), .A2(KEYINPUT79), .A3(new_n239), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n385), .B1(new_n384), .B2(new_n386), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n389), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n398), .B1(new_n408), .B2(new_n409), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n368), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(KEYINPUT5), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n405), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n415), .A3(new_n392), .ZN(new_n416));
  XOR2_X1   g215(.A(KEYINPUT81), .B(KEYINPUT6), .Z(new_n417));
  NAND3_X1  g216(.A1(new_n406), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT82), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n415), .B1(new_n414), .B2(new_n392), .ZN(new_n420));
  INV_X1    g219(.A(new_n417), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AND4_X1   g221(.A1(new_n419), .A2(new_n400), .A3(new_n405), .A4(new_n421), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n418), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n261), .B1(new_n347), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n261), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n339), .A2(KEYINPUT30), .ZN(new_n428));
  INV_X1    g227(.A(new_n338), .ZN(new_n429));
  AND4_X1   g228(.A1(new_n344), .A2(new_n346), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n388), .A2(new_n390), .A3(new_n366), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n368), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n432), .B(KEYINPUT39), .C1(new_n368), .C2(new_n412), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT39), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n431), .A2(new_n434), .A3(new_n368), .ZN(new_n435));
  AND3_X1   g234(.A1(new_n435), .A2(KEYINPUT85), .A3(new_n415), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT85), .B1(new_n435), .B2(new_n415), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n433), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT40), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(KEYINPUT40), .B(new_n433), .C1(new_n436), .C2(new_n437), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(new_n406), .A3(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n427), .B1(new_n430), .B2(new_n442), .ZN(new_n443));
  OAI211_X1 g242(.A(new_n418), .B(new_n342), .C1(new_n422), .C2(new_n423), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT37), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n316), .A2(new_n329), .ZN(new_n446));
  INV_X1    g245(.A(new_n262), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n233), .B1(new_n316), .B2(new_n329), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n333), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT86), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(new_n341), .B2(new_n445), .ZN(new_n452));
  AOI211_X1 g251(.A(KEYINPUT86), .B(KEYINPUT37), .C1(new_n330), .C2(new_n337), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT38), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n330), .A2(new_n337), .A3(KEYINPUT37), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n333), .A2(new_n455), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n457), .B(new_n458), .C1(new_n452), .C2(new_n453), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n444), .B1(new_n456), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n426), .B1(new_n443), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n315), .A2(new_n384), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n322), .A2(new_n365), .A3(new_n328), .ZN(new_n463));
  INV_X1    g262(.A(G227gat), .ZN(new_n464));
  INV_X1    g263(.A(G233gat), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n462), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT32), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT33), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  XOR2_X1   g269(.A(G15gat), .B(G43gat), .Z(new_n471));
  XNOR2_X1  g270(.A(G71gat), .B(G99gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n471), .B(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n468), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n473), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n467), .B(KEYINPUT32), .C1(new_n469), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n463), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n478), .B1(new_n464), .B2(new_n465), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT34), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT34), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n478), .B(new_n481), .C1(new_n464), .C2(new_n465), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n474), .A2(new_n480), .A3(new_n482), .A4(new_n476), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(KEYINPUT72), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT72), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n477), .A2(new_n487), .A3(new_n483), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT74), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n477), .A2(KEYINPUT74), .A3(new_n483), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n485), .A3(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n494));
  AOI22_X1  g293(.A1(KEYINPUT36), .A2(new_n489), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT35), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n261), .B1(new_n486), .B2(new_n488), .ZN(new_n497));
  AND4_X1   g296(.A1(new_n424), .A2(new_n340), .A3(new_n344), .A4(new_n346), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n496), .B(new_n256), .C1(new_n259), .C2(new_n260), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n430), .A2(new_n424), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n502), .A2(new_n493), .ZN(new_n503));
  OAI22_X1  g302(.A1(new_n461), .A2(new_n495), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  XOR2_X1   g303(.A(G71gat), .B(G78gat), .Z(new_n505));
  INV_X1    g304(.A(KEYINPUT9), .ZN(new_n506));
  XNOR2_X1  g305(.A(G57gat), .B(G64gat), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n505), .B(KEYINPUT91), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT91), .ZN(new_n509));
  INV_X1    g308(.A(G57gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(G64gat), .ZN(new_n511));
  INV_X1    g310(.A(G64gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(G57gat), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n506), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g313(.A1(G71gat), .A2(G78gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(G71gat), .A2(G78gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n509), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n508), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT92), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(new_n512), .B2(G57gat), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT93), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(new_n510), .B2(G64gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n510), .A2(KEYINPUT92), .A3(G64gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n512), .A2(KEYINPUT93), .A3(G57gat), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n521), .A2(new_n523), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT94), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n516), .B1(new_n515), .B2(new_n506), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n527), .B1(new_n526), .B2(new_n528), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n519), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT21), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G231gat), .A2(G233gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(G127gat), .B(G155gat), .Z(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT20), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n535), .B(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G183gat), .B(G211gat), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n538), .B(new_n539), .Z(new_n540));
  XNOR2_X1  g339(.A(G15gat), .B(G22gat), .ZN(new_n541));
  INV_X1    g340(.A(G1gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT16), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT88), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n546), .B1(new_n541), .B2(G1gat), .ZN(new_n547));
  OAI21_X1  g346(.A(G8gat), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  OR2_X1    g347(.A1(new_n541), .A2(G1gat), .ZN(new_n549));
  INV_X1    g348(.A(G8gat), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n549), .A2(new_n544), .A3(new_n546), .A4(new_n550), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(new_n531), .B2(new_n532), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT95), .B(KEYINPUT19), .Z(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n538), .B(new_n539), .ZN(new_n557));
  INV_X1    g356(.A(new_n555), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G113gat), .B(G141gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(G197gat), .ZN(new_n563));
  XOR2_X1   g362(.A(KEYINPUT11), .B(G169gat), .Z(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n565), .B(KEYINPUT12), .Z(new_n566));
  NAND2_X1  g365(.A1(new_n548), .A2(new_n551), .ZN(new_n567));
  INV_X1    g366(.A(G29gat), .ZN(new_n568));
  INV_X1    g367(.A(G36gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT14), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT14), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n571), .B1(G29gat), .B2(G36gat), .ZN(new_n572));
  AND2_X1   g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G43gat), .B(G50gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT15), .ZN(new_n575));
  NAND2_X1  g374(.A1(G29gat), .A2(G36gat), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT87), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(G43gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n252), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT15), .ZN(new_n581));
  NAND2_X1  g380(.A1(G43gat), .A2(G50gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n573), .A2(new_n575), .A3(new_n578), .A4(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n570), .A2(new_n572), .A3(new_n576), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(KEYINPUT15), .A3(new_n574), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n567), .B(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G229gat), .A2(G233gat), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n589), .B(KEYINPUT13), .Z(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n589), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT17), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n584), .A2(new_n593), .A3(new_n586), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n593), .B1(new_n584), .B2(new_n586), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n552), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n567), .A2(new_n587), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(KEYINPUT89), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT89), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n552), .B(new_n600), .C1(new_n595), .C2(new_n596), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n592), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n591), .B1(new_n602), .B2(KEYINPUT18), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n598), .A2(KEYINPUT89), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n587), .A2(KEYINPUT17), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n567), .B1(new_n605), .B2(new_n594), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n601), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n607), .A2(KEYINPUT18), .A3(new_n589), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n566), .B1(new_n603), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT90), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n607), .A2(new_n589), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT18), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n566), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n614), .A2(new_n615), .A3(new_n608), .A4(new_n591), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n610), .A2(new_n611), .A3(new_n616), .ZN(new_n617));
  OAI211_X1 g416(.A(KEYINPUT90), .B(new_n566), .C1(new_n603), .C2(new_n609), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(G85gat), .ZN(new_n620));
  INV_X1    g419(.A(G92gat), .ZN(new_n621));
  OAI21_X1  g420(.A(KEYINPUT7), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT7), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n623), .A2(G85gat), .A3(G92gat), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G99gat), .A2(G106gat), .ZN(new_n626));
  AOI22_X1  g425(.A1(KEYINPUT8), .A2(new_n626), .B1(new_n620), .B2(new_n621), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G99gat), .B(G106gat), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n625), .A2(new_n629), .A3(new_n627), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n531), .A2(new_n633), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n625), .A2(new_n629), .A3(new_n627), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n629), .B1(new_n625), .B2(new_n627), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n637), .B(new_n519), .C1(new_n530), .C2(new_n529), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT10), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n634), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n531), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n642), .B1(new_n635), .B2(new_n636), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n631), .A2(KEYINPUT97), .A3(new_n632), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n641), .A2(KEYINPUT10), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(G230gat), .A2(G233gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n648), .B1(new_n634), .B2(new_n638), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G120gat), .B(G148gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(G176gat), .B(G204gat), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n652), .B(new_n653), .Z(new_n654));
  NAND3_X1  g453(.A1(new_n649), .A2(new_n651), .A3(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(KEYINPUT99), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n657));
  INV_X1    g456(.A(new_n648), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n658), .B1(new_n640), .B2(new_n646), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n659), .A2(new_n650), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n657), .B1(new_n660), .B2(new_n654), .ZN(new_n661));
  OAI22_X1  g460(.A1(new_n656), .A2(new_n661), .B1(new_n660), .B2(new_n654), .ZN(new_n662));
  XNOR2_X1  g461(.A(G190gat), .B(G218gat), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT98), .ZN(new_n665));
  NAND3_X1  g464(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n666), .B1(new_n664), .B2(KEYINPUT98), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n667), .B1(new_n645), .B2(new_n587), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n644), .B(new_n643), .C1(new_n595), .C2(new_n596), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n665), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n672));
  XOR2_X1   g471(.A(new_n672), .B(KEYINPUT96), .Z(new_n673));
  XNOR2_X1  g472(.A(G134gat), .B(G162gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n668), .A2(new_n669), .A3(new_n665), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n671), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n675), .ZN(new_n678));
  INV_X1    g477(.A(new_n676), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n679), .B2(new_n670), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NOR4_X1   g480(.A1(new_n561), .A2(new_n619), .A3(new_n662), .A4(new_n681), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n504), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n425), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g484(.A(KEYINPUT100), .B(KEYINPUT16), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(new_n550), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n683), .A2(new_n347), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n683), .ZN(new_n691));
  OAI21_X1  g490(.A(G8gat), .B1(new_n691), .B2(new_n430), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n688), .A2(new_n689), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(G1325gat));
  NAND2_X1  g493(.A1(new_n489), .A2(KEYINPUT36), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n493), .A2(new_n494), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G15gat), .B1(new_n691), .B2(new_n697), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n493), .A2(G15gat), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n698), .B1(new_n691), .B2(new_n699), .ZN(G1326gat));
  NAND2_X1  g499(.A1(new_n683), .A2(new_n261), .ZN(new_n701));
  XNOR2_X1  g500(.A(KEYINPUT43), .B(G22gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1327gat));
  INV_X1    g502(.A(new_n681), .ZN(new_n704));
  INV_X1    g503(.A(new_n442), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n261), .B1(new_n705), .B2(new_n347), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n457), .A2(new_n458), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n341), .A2(new_n445), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT86), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n341), .A2(new_n451), .A3(new_n445), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n707), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n455), .B2(new_n454), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n706), .B1(new_n712), .B2(new_n444), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n713), .A3(new_n426), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n489), .A2(new_n498), .A3(new_n427), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(KEYINPUT35), .ZN(new_n716));
  INV_X1    g515(.A(new_n493), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n717), .A2(new_n498), .A3(new_n501), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n704), .B1(new_n714), .B2(new_n719), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n560), .A2(new_n619), .A3(new_n662), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n722), .A2(new_n568), .A3(new_n425), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT45), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n427), .B1(new_n430), .B2(new_n424), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n456), .A2(new_n459), .ZN(new_n727));
  INV_X1    g526(.A(new_n444), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n726), .B1(new_n729), .B2(new_n706), .ZN(new_n730));
  AOI22_X1  g529(.A1(new_n730), .A2(new_n697), .B1(new_n716), .B2(new_n718), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n725), .B1(new_n731), .B2(new_n704), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n504), .A2(KEYINPUT44), .A3(new_n681), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n721), .B(KEYINPUT101), .Z(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(G29gat), .B1(new_n736), .B2(new_n424), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n724), .A2(new_n737), .ZN(G1328gat));
  NAND3_X1  g537(.A1(new_n722), .A2(new_n569), .A3(new_n347), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(KEYINPUT46), .Z(new_n740));
  OAI21_X1  g539(.A(G36gat), .B1(new_n736), .B2(new_n430), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(G1329gat));
  NAND4_X1  g541(.A1(new_n732), .A2(new_n495), .A3(new_n733), .A4(new_n735), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(G43gat), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n722), .A2(new_n579), .A3(new_n717), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT47), .B1(new_n745), .B2(KEYINPUT102), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1330gat));
  NAND4_X1  g547(.A1(new_n732), .A2(new_n261), .A3(new_n733), .A4(new_n735), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G50gat), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT103), .ZN(new_n751));
  AOI21_X1  g550(.A(KEYINPUT48), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n722), .A2(new_n252), .A3(new_n261), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n750), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n752), .B(new_n754), .ZN(G1331gat));
  NAND3_X1  g554(.A1(new_n560), .A2(new_n619), .A3(new_n704), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n660), .A2(new_n654), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n655), .A2(KEYINPUT99), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n660), .A2(new_n657), .A3(new_n654), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n756), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n504), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT104), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n504), .A2(KEYINPUT104), .A3(new_n761), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n766), .A2(new_n424), .ZN(new_n767));
  XOR2_X1   g566(.A(KEYINPUT105), .B(G57gat), .Z(new_n768));
  XNOR2_X1  g567(.A(new_n767), .B(new_n768), .ZN(G1332gat));
  NOR2_X1   g568(.A1(new_n766), .A2(new_n430), .ZN(new_n770));
  NOR2_X1   g569(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n771));
  AND2_X1   g570(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n770), .B2(new_n771), .ZN(G1333gat));
  OR3_X1    g573(.A1(new_n766), .A2(G71gat), .A3(new_n493), .ZN(new_n775));
  OAI21_X1  g574(.A(G71gat), .B1(new_n766), .B2(new_n697), .ZN(new_n776));
  XNOR2_X1  g575(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n775), .B2(new_n776), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n778), .A2(new_n779), .ZN(G1334gat));
  NOR2_X1   g579(.A1(new_n766), .A2(new_n427), .ZN(new_n781));
  XOR2_X1   g580(.A(new_n781), .B(G78gat), .Z(G1335gat));
  INV_X1    g581(.A(new_n619), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n560), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT51), .B1(new_n720), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n785), .A2(KEYINPUT107), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n504), .A2(new_n681), .ZN(new_n788));
  INV_X1    g587(.A(new_n784), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n720), .A2(KEYINPUT51), .A3(new_n784), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n786), .B1(KEYINPUT107), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n425), .A2(new_n620), .A3(new_n662), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n789), .A2(new_n760), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n734), .A2(new_n425), .A3(new_n795), .ZN(new_n796));
  OAI22_X1  g595(.A1(new_n793), .A2(new_n794), .B1(new_n796), .B2(new_n620), .ZN(G1336gat));
  NOR3_X1   g596(.A1(new_n430), .A2(G92gat), .A3(new_n760), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n793), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n732), .A2(new_n347), .A3(new_n733), .A4(new_n795), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G92gat), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n792), .A2(new_n798), .B1(new_n801), .B2(G92gat), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n800), .A2(new_n804), .B1(new_n803), .B2(new_n805), .ZN(G1337gat));
  NAND3_X1  g605(.A1(new_n734), .A2(new_n495), .A3(new_n795), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT108), .ZN(new_n808));
  XNOR2_X1  g607(.A(KEYINPUT109), .B(G99gat), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n807), .A2(KEYINPUT108), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n717), .A2(new_n662), .A3(new_n809), .ZN(new_n813));
  OAI22_X1  g612(.A1(new_n811), .A2(new_n812), .B1(new_n793), .B2(new_n813), .ZN(G1338gat));
  NAND4_X1  g613(.A1(new_n732), .A2(new_n261), .A3(new_n733), .A4(new_n795), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT53), .B1(new_n815), .B2(G106gat), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n427), .A2(G106gat), .A3(new_n760), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n816), .B1(new_n793), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT110), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n815), .A2(G106gat), .ZN(new_n821));
  AND4_X1   g620(.A1(KEYINPUT51), .A2(new_n504), .A3(new_n681), .A4(new_n784), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n817), .B1(new_n785), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n820), .B1(new_n824), .B2(KEYINPUT53), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n826));
  AOI211_X1 g625(.A(KEYINPUT110), .B(new_n826), .C1(new_n821), .C2(new_n823), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n819), .B1(new_n825), .B2(new_n827), .ZN(G1339gat));
  NAND4_X1  g627(.A1(new_n560), .A2(new_n619), .A3(new_n760), .A4(new_n704), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n640), .A2(new_n646), .A3(new_n658), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n649), .A2(KEYINPUT54), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT111), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n834), .B1(new_n647), .B2(new_n648), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(KEYINPUT111), .A3(new_n830), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n654), .B1(new_n659), .B2(new_n834), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n838), .A2(KEYINPUT55), .ZN(new_n839));
  AOI22_X1  g638(.A1(new_n837), .A2(new_n839), .B1(new_n758), .B2(new_n759), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n835), .A2(KEYINPUT111), .A3(new_n830), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT111), .B1(new_n835), .B2(new_n830), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n838), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI22_X1  g644(.A1(new_n607), .A2(new_n589), .B1(new_n588), .B2(new_n590), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n565), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n616), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n704), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n840), .A2(new_n845), .A3(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n839), .B1(new_n841), .B2(new_n842), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n758), .A2(new_n759), .ZN(new_n853));
  INV_X1    g652(.A(new_n838), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n854), .B1(new_n833), .B2(new_n836), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n852), .B(new_n853), .C1(new_n855), .C2(KEYINPUT55), .ZN(new_n856));
  OAI22_X1  g655(.A1(new_n856), .A2(new_n619), .B1(new_n760), .B2(new_n848), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n851), .B1(new_n857), .B2(new_n704), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n829), .B1(new_n858), .B2(new_n560), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n859), .A2(new_n427), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n347), .A2(new_n424), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(new_n493), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n349), .B1(new_n864), .B2(new_n783), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(KEYINPUT112), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n859), .A2(new_n425), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n497), .A2(new_n430), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n783), .A2(new_n349), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT113), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n866), .B1(new_n869), .B2(new_n871), .ZN(G1340gat));
  INV_X1    g671(.A(new_n864), .ZN(new_n873));
  OAI21_X1  g672(.A(G120gat), .B1(new_n873), .B2(new_n760), .ZN(new_n874));
  INV_X1    g673(.A(new_n869), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n352), .A3(new_n662), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(G1341gat));
  OAI21_X1  g676(.A(new_n377), .B1(new_n873), .B2(new_n561), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n875), .A2(new_n360), .A3(new_n560), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1342gat));
  NAND3_X1  g679(.A1(new_n875), .A2(new_n355), .A3(new_n681), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n881), .A2(KEYINPUT56), .ZN(new_n882));
  OAI21_X1  g681(.A(G134gat), .B1(new_n873), .B2(new_n704), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(KEYINPUT56), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(G1343gat));
  NOR3_X1   g684(.A1(new_n495), .A2(new_n347), .A3(new_n427), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n619), .A2(G141gat), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT115), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n867), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT116), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT58), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT116), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n867), .A2(new_n892), .A3(new_n886), .A4(new_n888), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n859), .A2(new_n895), .A3(new_n261), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n495), .A2(new_n862), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n856), .A2(new_n619), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT114), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n662), .A2(new_n899), .A3(new_n616), .A4(new_n847), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT114), .B1(new_n760), .B2(new_n848), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n704), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n560), .B1(new_n903), .B2(new_n850), .ZN(new_n904));
  INV_X1    g703(.A(new_n829), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(new_n427), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n896), .B(new_n897), .C1(new_n907), .C2(new_n895), .ZN(new_n908));
  OAI21_X1  g707(.A(G141gat), .B1(new_n908), .B2(new_n619), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n894), .A2(KEYINPUT117), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(KEYINPUT117), .B1(new_n894), .B2(new_n909), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n909), .A2(new_n889), .ZN(new_n912));
  OAI22_X1  g711(.A1(new_n910), .A2(new_n911), .B1(new_n891), .B2(new_n912), .ZN(G1344gat));
  NAND2_X1  g712(.A1(new_n867), .A2(new_n886), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(new_n211), .A3(new_n662), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT59), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT118), .B1(new_n904), .B2(new_n905), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT118), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n901), .B(new_n900), .C1(new_n856), .C2(new_n619), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n851), .B1(new_n920), .B2(new_n704), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n919), .B(new_n829), .C1(new_n921), .C2(new_n560), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n427), .A2(KEYINPUT57), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n918), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n859), .A2(new_n261), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT57), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n924), .A2(new_n662), .A3(new_n926), .A4(new_n897), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT119), .ZN(new_n928));
  OR2_X1    g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n211), .B1(new_n927), .B2(new_n928), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n917), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n908), .ZN(new_n932));
  AOI211_X1 g731(.A(KEYINPUT59), .B(new_n211), .C1(new_n932), .C2(new_n662), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n916), .B1(new_n931), .B2(new_n933), .ZN(G1345gat));
  OAI21_X1  g733(.A(G155gat), .B1(new_n908), .B2(new_n561), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n915), .A2(new_n215), .A3(new_n560), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1346gat));
  AOI21_X1  g736(.A(G162gat), .B1(new_n915), .B2(new_n681), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n704), .A2(new_n216), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n938), .B1(new_n932), .B2(new_n939), .ZN(G1347gat));
  NOR2_X1   g739(.A1(new_n430), .A2(new_n425), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n859), .A2(new_n717), .A3(new_n427), .A4(new_n941), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n942), .A2(new_n272), .A3(new_n619), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n859), .A2(new_n424), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n497), .A2(new_n347), .ZN(new_n945));
  XOR2_X1   g744(.A(new_n945), .B(KEYINPUT120), .Z(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT121), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT121), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n944), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(new_n783), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n943), .B1(new_n952), .B2(new_n272), .ZN(G1348gat));
  NAND3_X1  g752(.A1(new_n948), .A2(new_n662), .A3(new_n950), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n954), .A2(KEYINPUT122), .A3(new_n273), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n942), .A2(new_n273), .A3(new_n760), .ZN(new_n956));
  XOR2_X1   g755(.A(new_n956), .B(KEYINPUT123), .Z(new_n957));
  AOI21_X1  g756(.A(KEYINPUT122), .B1(new_n954), .B2(new_n273), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n955), .A2(new_n957), .A3(new_n958), .ZN(G1349gat));
  OAI21_X1  g758(.A(G183gat), .B1(new_n942), .B2(new_n561), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n560), .A2(new_n283), .A3(new_n287), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n960), .B1(new_n947), .B2(new_n961), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g762(.A1(new_n951), .A2(new_n284), .A3(new_n681), .ZN(new_n964));
  OAI21_X1  g763(.A(G190gat), .B1(new_n942), .B2(new_n704), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT61), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n966), .ZN(G1351gat));
  NOR3_X1   g766(.A1(new_n495), .A2(new_n430), .A3(new_n427), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n944), .A2(new_n968), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n969), .A2(G197gat), .A3(new_n619), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n970), .B(KEYINPUT124), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n697), .A2(new_n941), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n924), .A2(new_n926), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(new_n783), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(G197gat), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n971), .A2(new_n975), .ZN(G1352gat));
  NAND4_X1  g775(.A1(new_n924), .A2(new_n662), .A3(new_n926), .A4(new_n972), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(G204gat), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n760), .A2(G204gat), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n944), .A2(new_n968), .A3(new_n979), .ZN(new_n980));
  OR2_X1    g779(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n978), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n983), .B(KEYINPUT125), .ZN(G1353gat));
  NAND4_X1  g783(.A1(new_n944), .A2(new_n225), .A3(new_n560), .A4(new_n968), .ZN(new_n985));
  NAND4_X1  g784(.A1(new_n924), .A2(new_n560), .A3(new_n926), .A4(new_n972), .ZN(new_n986));
  AND3_X1   g785(.A1(new_n986), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n987));
  AOI21_X1  g786(.A(KEYINPUT63), .B1(new_n986), .B2(G211gat), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT126), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI211_X1 g790(.A(KEYINPUT126), .B(new_n985), .C1(new_n987), .C2(new_n988), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(G1354gat));
  NAND2_X1  g792(.A1(new_n681), .A2(G218gat), .ZN(new_n994));
  XNOR2_X1  g793(.A(new_n994), .B(KEYINPUT127), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n944), .A2(new_n681), .A3(new_n968), .ZN(new_n996));
  AOI22_X1  g795(.A1(new_n973), .A2(new_n995), .B1(new_n226), .B2(new_n996), .ZN(G1355gat));
endmodule


