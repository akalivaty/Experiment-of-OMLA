//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  NAND2_X1  g000(.A1(G234), .A2(G237), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND3_X1   g002(.A1(new_n187), .A2(G952), .A3(new_n188), .ZN(new_n189));
  AND3_X1   g003(.A1(new_n187), .A2(G902), .A3(G953), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT21), .B(G898), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n189), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G478), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(KEYINPUT15), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G902), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT93), .ZN(new_n198));
  INV_X1    g012(.A(G128), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(G143), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT93), .A3(G128), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(G143), .ZN(new_n204));
  AND3_X1   g018(.A1(new_n203), .A2(KEYINPUT95), .A3(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT95), .B1(new_n203), .B2(new_n204), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n197), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  AND3_X1   g021(.A1(new_n201), .A2(KEYINPUT93), .A3(G128), .ZN(new_n208));
  AOI21_X1  g022(.A(KEYINPUT93), .B1(new_n201), .B2(G128), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n204), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT95), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n203), .A2(KEYINPUT95), .A3(new_n204), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(G134), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n207), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G107), .ZN(new_n216));
  INV_X1    g030(.A(G122), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G116), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n216), .B1(new_n218), .B2(KEYINPUT14), .ZN(new_n219));
  XNOR2_X1  g033(.A(G116), .B(G122), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n219), .A2(new_n220), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(KEYINPUT97), .B1(new_n215), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT97), .ZN(new_n226));
  AOI211_X1 g040(.A(new_n226), .B(new_n223), .C1(new_n207), .C2(new_n214), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n220), .B(G107), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n212), .A2(new_n213), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(new_n197), .ZN(new_n230));
  XOR2_X1   g044(.A(KEYINPUT94), .B(KEYINPUT13), .Z(new_n231));
  OAI21_X1  g045(.A(new_n204), .B1(new_n231), .B2(new_n203), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n231), .A2(new_n203), .ZN(new_n233));
  OAI21_X1  g047(.A(G134), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(KEYINPUT96), .B1(new_n230), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n228), .ZN(new_n236));
  AND4_X1   g050(.A1(KEYINPUT96), .A2(new_n234), .A3(new_n207), .A4(new_n236), .ZN(new_n237));
  OAI22_X1  g051(.A1(new_n225), .A2(new_n227), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT9), .B(G234), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT74), .B(G217), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(new_n188), .A3(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n238), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n242), .ZN(new_n244));
  NOR3_X1   g058(.A1(new_n205), .A2(new_n206), .A3(new_n197), .ZN(new_n245));
  AOI21_X1  g059(.A(G134), .B1(new_n212), .B2(new_n213), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n224), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n226), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n215), .A2(KEYINPUT97), .A3(new_n224), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n234), .A2(new_n207), .A3(new_n236), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT96), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n230), .A2(KEYINPUT96), .A3(new_n234), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n244), .B1(new_n250), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n196), .B1(new_n243), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT98), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n238), .A2(new_n242), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n250), .A2(new_n255), .A3(new_n244), .ZN(new_n260));
  AOI21_X1  g074(.A(G902), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT98), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n195), .B1(new_n258), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n261), .A2(new_n262), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(new_n194), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT99), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  AOI211_X1 g081(.A(KEYINPUT98), .B(G902), .C1(new_n259), .C2(new_n260), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n194), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT99), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n258), .A2(new_n195), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n192), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G469), .ZN(new_n274));
  XNOR2_X1  g088(.A(G110), .B(G140), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n275), .B(KEYINPUT81), .ZN(new_n276));
  INV_X1    g090(.A(G227), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(G953), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n276), .B(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT10), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT82), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n199), .A2(KEYINPUT1), .ZN(new_n282));
  INV_X1    g096(.A(G146), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G143), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n201), .A2(G146), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n282), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT67), .ZN(new_n287));
  XNOR2_X1  g101(.A(G143), .B(G146), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT67), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n289), .A3(new_n282), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n288), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT1), .B1(new_n201), .B2(G146), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G128), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G104), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT3), .B1(new_n297), .B2(G107), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT3), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(new_n216), .A3(G104), .ZN(new_n300));
  INV_X1    g114(.A(G101), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n297), .A2(G107), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n298), .A2(new_n300), .A3(new_n301), .A4(new_n302), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n216), .A2(G104), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n297), .A2(G107), .ZN(new_n305));
  OAI21_X1  g119(.A(G101), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n281), .B1(new_n296), .B2(new_n307), .ZN(new_n308));
  AOI22_X1  g122(.A1(new_n287), .A2(new_n290), .B1(new_n292), .B2(new_n294), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n303), .A2(new_n306), .ZN(new_n310));
  NOR3_X1   g124(.A1(new_n309), .A2(KEYINPUT82), .A3(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n280), .B1(new_n308), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT68), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n293), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT1), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n315), .B1(G143), .B2(new_n283), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n199), .B1(new_n316), .B2(KEYINPUT68), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n201), .A2(KEYINPUT65), .A3(G146), .ZN(new_n318));
  AOI21_X1  g132(.A(KEYINPUT65), .B1(new_n201), .B2(G146), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT64), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(new_n201), .B2(G146), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n283), .A2(KEYINPUT64), .A3(G143), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n314), .A2(new_n317), .B1(new_n320), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n289), .B1(new_n288), .B2(new_n282), .ZN(new_n326));
  AND4_X1   g140(.A1(new_n289), .A2(new_n282), .A3(new_n284), .A4(new_n285), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(KEYINPUT70), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n284), .A2(KEYINPUT68), .A3(KEYINPUT1), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n314), .A2(G128), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n319), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n201), .A2(KEYINPUT65), .A3(G146), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n324), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT70), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n336), .A3(new_n291), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n329), .A2(KEYINPUT10), .A3(new_n337), .A4(new_n307), .ZN(new_n338));
  AND2_X1   g152(.A1(KEYINPUT0), .A2(G128), .ZN(new_n339));
  NOR2_X1   g153(.A1(KEYINPUT0), .A2(G128), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI22_X1  g155(.A1(new_n334), .A2(new_n341), .B1(new_n288), .B2(new_n339), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n298), .A2(new_n300), .A3(new_n302), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT4), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(G101), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(G101), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(KEYINPUT4), .A3(new_n303), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n342), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n312), .A2(new_n338), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT85), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n197), .A2(G137), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n197), .A2(G137), .ZN(new_n352));
  NAND2_X1  g166(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n351), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G137), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G134), .ZN(new_n357));
  OR2_X1    g171(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n357), .B1(new_n358), .B2(new_n353), .ZN(new_n359));
  OAI21_X1  g173(.A(G131), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n356), .A2(G134), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n361), .B1(new_n357), .B2(new_n353), .ZN(new_n362));
  INV_X1    g176(.A(G131), .ZN(new_n363));
  NOR2_X1   g177(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n352), .B1(new_n354), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n362), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT85), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n312), .A2(new_n368), .A3(new_n338), .A4(new_n348), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n350), .A2(new_n367), .A3(new_n369), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n360), .A2(new_n366), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n312), .A2(new_n371), .A3(new_n338), .A4(new_n348), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n279), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n296), .A2(new_n281), .A3(new_n307), .ZN(new_n374));
  OAI21_X1  g188(.A(KEYINPUT82), .B1(new_n309), .B2(new_n310), .ZN(new_n375));
  AOI22_X1  g189(.A1(new_n331), .A2(new_n334), .B1(new_n287), .B2(new_n290), .ZN(new_n376));
  AOI22_X1  g190(.A1(new_n374), .A2(new_n375), .B1(new_n376), .B2(new_n310), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(new_n371), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT12), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(KEYINPUT83), .A3(new_n379), .ZN(new_n380));
  OR2_X1    g194(.A1(new_n379), .A2(KEYINPUT83), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(KEYINPUT83), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n381), .B(new_n382), .C1(new_n377), .C2(new_n371), .ZN(new_n383));
  AND4_X1   g197(.A1(new_n372), .A2(new_n380), .A3(new_n279), .A4(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n274), .B(new_n196), .C1(new_n373), .C2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n274), .A2(new_n196), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n372), .ZN(new_n388));
  INV_X1    g202(.A(new_n279), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT84), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT84), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n372), .A2(new_n391), .A3(new_n279), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n370), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n380), .A2(new_n372), .A3(new_n383), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n389), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(G469), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n385), .A2(new_n387), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G221), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n398), .B1(new_n240), .B2(new_n196), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G140), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G125), .ZN(new_n403));
  INV_X1    g217(.A(G125), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G140), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(KEYINPUT79), .A3(new_n283), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT79), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n403), .A2(new_n405), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n408), .B1(new_n409), .B2(G146), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(G146), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(KEYINPUT71), .A2(G237), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(KEYINPUT71), .A2(G237), .ZN(new_n416));
  OAI211_X1 g230(.A(G214), .B(new_n188), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n201), .ZN(new_n418));
  XNOR2_X1  g232(.A(KEYINPUT71), .B(G237), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n419), .A2(G143), .A3(G214), .A4(new_n188), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(KEYINPUT18), .A2(G131), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n418), .A2(new_n420), .A3(new_n422), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n413), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT16), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n402), .A3(G125), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(KEYINPUT77), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n406), .A2(KEYINPUT76), .A3(KEYINPUT16), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT76), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n409), .B2(new_n427), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n283), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n421), .A2(KEYINPUT17), .A3(G131), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n429), .A2(new_n430), .A3(G146), .A4(new_n432), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  AND3_X1   g251(.A1(new_n418), .A2(new_n420), .A3(new_n363), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n363), .B1(new_n418), .B2(new_n420), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT17), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n426), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(G113), .B(G122), .ZN(new_n442));
  XNOR2_X1  g256(.A(KEYINPUT88), .B(G104), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n442), .B(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  AND2_X1   g259(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n444), .B(KEYINPUT89), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n426), .B(new_n447), .C1(new_n437), .C2(new_n440), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n196), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT91), .B(G475), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n406), .A2(KEYINPUT19), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n403), .A2(new_n405), .A3(KEYINPUT19), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n283), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n436), .B(new_n455), .C1(new_n438), .C2(new_n439), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n426), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n445), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(new_n448), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT20), .ZN(new_n460));
  NOR2_X1   g274(.A1(G475), .A2(G902), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n459), .A2(KEYINPUT90), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n461), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n463), .B1(new_n458), .B2(new_n448), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n462), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT90), .B1(new_n464), .B2(new_n460), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n452), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT92), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n464), .A2(new_n460), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT90), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n459), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT20), .B1(new_n473), .B2(new_n463), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n472), .A2(new_n462), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(KEYINPUT92), .A3(new_n452), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n273), .A2(new_n401), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(G214), .B1(G237), .B2(G902), .ZN(new_n480));
  XNOR2_X1  g294(.A(G110), .B(G122), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT8), .ZN(new_n482));
  OR2_X1    g296(.A1(KEYINPUT69), .A2(G119), .ZN(new_n483));
  NAND2_X1  g297(.A1(KEYINPUT69), .A2(G119), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(G116), .A3(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT86), .B(KEYINPUT5), .ZN(new_n486));
  OAI21_X1  g300(.A(G113), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G116), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(G119), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n487), .B1(new_n491), .B2(KEYINPUT5), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT2), .B(G113), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(new_n485), .A3(new_n489), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n307), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n485), .A2(new_n489), .A3(new_n486), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n498), .B(G113), .C1(new_n485), .C2(new_n486), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n307), .B1(new_n499), .B2(new_n495), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n482), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n335), .A2(new_n404), .A3(new_n291), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n502), .B1(new_n404), .B2(new_n342), .ZN(new_n503));
  INV_X1    g317(.A(G224), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT7), .B1(new_n504), .B2(G953), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n490), .A2(new_n493), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n495), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n345), .A3(new_n347), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n499), .A2(new_n307), .A3(new_n495), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n510), .A3(new_n481), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n501), .A2(new_n506), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n505), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n502), .B(new_n513), .C1(new_n404), .C2(new_n342), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT87), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(G902), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(G210), .B1(G237), .B2(G902), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n504), .A2(G953), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n503), .B(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n509), .A2(new_n510), .ZN(new_n521));
  INV_X1    g335(.A(new_n481), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(KEYINPUT6), .A3(new_n511), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT6), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n521), .A2(new_n525), .A3(new_n522), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n520), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n517), .A2(new_n518), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n518), .B1(new_n517), .B2(new_n527), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n480), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(G472), .A2(G902), .ZN(new_n531));
  OAI21_X1  g345(.A(G131), .B1(new_n352), .B2(new_n361), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n366), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n329), .A2(new_n337), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT30), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n536), .B1(new_n367), .B2(new_n342), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n334), .A2(new_n341), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n288), .A2(new_n339), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI22_X1  g355(.A1(new_n371), .A2(new_n541), .B1(new_n376), .B2(new_n533), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n536), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n538), .A2(new_n508), .A3(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n508), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n367), .A2(new_n342), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n535), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n419), .A2(G210), .A3(new_n188), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(KEYINPUT27), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT26), .B(G101), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT31), .B1(new_n544), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n538), .A2(new_n543), .A3(new_n508), .ZN(new_n554));
  XOR2_X1   g368(.A(KEYINPUT72), .B(KEYINPUT31), .Z(new_n555));
  NAND4_X1  g369(.A1(new_n554), .A2(new_n547), .A3(new_n551), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n542), .A2(new_n508), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n547), .A2(KEYINPUT28), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT28), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n535), .A2(new_n560), .A3(new_n545), .A4(new_n546), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n558), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(new_n551), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n531), .B1(new_n557), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT73), .B(KEYINPUT32), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n545), .B1(new_n535), .B2(new_n546), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(new_n559), .B2(new_n561), .ZN(new_n569));
  INV_X1    g383(.A(new_n551), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT29), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(G902), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n535), .A2(new_n545), .A3(new_n546), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n535), .A2(new_n537), .B1(new_n542), .B2(new_n536), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n574), .B1(new_n508), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n571), .B1(new_n576), .B2(new_n551), .ZN(new_n577));
  AOI211_X1 g391(.A(new_n570), .B(new_n558), .C1(new_n559), .C2(new_n561), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n573), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G472), .ZN(new_n580));
  OAI211_X1 g394(.A(KEYINPUT32), .B(new_n531), .C1(new_n557), .C2(new_n563), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n567), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(G234), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n241), .B1(new_n583), .B2(G902), .ZN(new_n584));
  XNOR2_X1  g398(.A(KEYINPUT22), .B(G137), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n398), .A2(new_n583), .A3(G953), .ZN(new_n586));
  XOR2_X1   g400(.A(new_n585), .B(new_n586), .Z(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n436), .A2(new_n411), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT23), .ZN(new_n590));
  XOR2_X1   g404(.A(KEYINPUT69), .B(G119), .Z(new_n591));
  OAI21_X1  g405(.A(new_n590), .B1(new_n591), .B2(G128), .ZN(new_n592));
  INV_X1    g406(.A(G110), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n483), .A2(G128), .A3(new_n484), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n199), .A2(KEYINPUT23), .A3(G119), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n592), .A2(new_n593), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT75), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n591), .A2(new_n598), .A3(G128), .ZN(new_n599));
  XNOR2_X1  g413(.A(KEYINPUT24), .B(G110), .ZN(new_n600));
  INV_X1    g414(.A(G119), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT75), .B1(new_n601), .B2(G128), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n599), .B(new_n600), .C1(new_n594), .C2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT78), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n597), .A2(new_n603), .A3(KEYINPUT78), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n589), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n434), .A2(new_n436), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n592), .A2(new_n595), .A3(new_n596), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n599), .B1(new_n594), .B2(new_n602), .ZN(new_n611));
  INV_X1    g425(.A(new_n600), .ZN(new_n612));
  AOI22_X1  g426(.A1(new_n610), .A2(G110), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n588), .B1(new_n608), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n589), .ZN(new_n616));
  INV_X1    g430(.A(new_n607), .ZN(new_n617));
  AOI21_X1  g431(.A(KEYINPUT78), .B1(new_n597), .B2(new_n603), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n609), .A2(new_n613), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(new_n620), .A3(new_n587), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n615), .A2(new_n621), .A3(new_n196), .ZN(new_n622));
  AND2_X1   g436(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n584), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n615), .A2(new_n621), .A3(new_n196), .A4(new_n626), .ZN(new_n627));
  AND2_X1   g441(.A1(new_n615), .A2(new_n621), .ZN(new_n628));
  AOI21_X1  g442(.A(G902), .B1(new_n241), .B2(new_n583), .ZN(new_n629));
  AOI22_X1  g443(.A1(new_n624), .A2(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n582), .A2(new_n630), .ZN(new_n631));
  OR3_X1    g445(.A1(new_n479), .A2(new_n530), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G101), .ZN(G3));
  OAI21_X1  g447(.A(new_n196), .B1(new_n557), .B2(new_n563), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(G472), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n635), .A2(new_n564), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n401), .A2(new_n630), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n530), .A2(new_n192), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT33), .B1(new_n243), .B2(new_n256), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT33), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n259), .A2(new_n640), .A3(new_n260), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n639), .A2(G478), .A3(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n193), .A2(new_n196), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n643), .B1(new_n261), .B2(new_n193), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n477), .A2(new_n638), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n637), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT34), .B(G104), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G6));
  AOI22_X1  g464(.A1(new_n474), .A2(new_n470), .B1(new_n450), .B2(new_n451), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n267), .A2(new_n272), .A3(new_n638), .A4(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n637), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT35), .B(G107), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  NAND2_X1  g470(.A1(new_n619), .A2(new_n620), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n588), .A2(KEYINPUT36), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(new_n659));
  AOI22_X1  g473(.A1(new_n624), .A2(new_n627), .B1(new_n629), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n530), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n636), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n479), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT100), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT37), .B(G110), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G12));
  INV_X1    g480(.A(G900), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n189), .B1(new_n190), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n267), .A2(new_n272), .A3(new_n651), .A4(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n582), .A2(new_n400), .A3(new_n397), .A4(new_n661), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G128), .ZN(G30));
  XOR2_X1   g489(.A(new_n668), .B(KEYINPUT39), .Z(new_n676));
  NAND2_X1  g490(.A1(new_n401), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n677), .B(KEYINPUT40), .Z(new_n678));
  NOR2_X1   g492(.A1(new_n576), .A2(new_n570), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n570), .A2(new_n547), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n196), .B1(new_n680), .B2(new_n568), .ZN(new_n681));
  OAI21_X1  g495(.A(G472), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n581), .A2(new_n682), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n553), .B(new_n556), .C1(new_n562), .C2(new_n551), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n565), .B1(new_n684), .B2(new_n531), .ZN(new_n685));
  OAI21_X1  g499(.A(KEYINPUT102), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT102), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n567), .A2(new_n687), .A3(new_n581), .A4(new_n682), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n660), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n267), .A2(new_n272), .ZN(new_n693));
  INV_X1    g507(.A(new_n529), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n517), .A2(new_n518), .A3(new_n527), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n480), .ZN(new_n699));
  NOR4_X1   g513(.A1(new_n693), .A2(new_n698), .A3(new_n478), .A4(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n678), .A2(new_n692), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G143), .ZN(G45));
  NOR2_X1   g516(.A1(new_n467), .A2(new_n468), .ZN(new_n703));
  AOI21_X1  g517(.A(KEYINPUT92), .B1(new_n475), .B2(new_n452), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n645), .B(new_n669), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n673), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  AND2_X1   g522(.A1(new_n582), .A2(new_n630), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n196), .B1(new_n373), .B2(new_n384), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(G469), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n711), .A2(new_n400), .A3(new_n385), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n647), .A2(new_n709), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NAND3_X1  g529(.A1(new_n653), .A2(new_n709), .A3(new_n712), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  AND2_X1   g531(.A1(new_n582), .A2(new_n691), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n699), .B1(new_n694), .B2(new_n695), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n711), .A2(new_n719), .A3(new_n400), .A4(new_n385), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n718), .A2(new_n273), .A3(new_n478), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G119), .ZN(G21));
  INV_X1    g537(.A(KEYINPUT103), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n635), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n634), .A2(KEYINPUT103), .A3(G472), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n553), .B(new_n556), .C1(new_n551), .C2(new_n569), .ZN(new_n727));
  AOI22_X1  g541(.A1(new_n725), .A2(new_n726), .B1(new_n531), .B2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n192), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(new_n729), .A3(new_n630), .A4(new_n712), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n267), .A2(new_n477), .A3(new_n272), .A4(new_n719), .ZN(new_n731));
  OR2_X1    g545(.A1(new_n731), .A2(KEYINPUT104), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(KEYINPUT104), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n730), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n217), .ZN(G24));
  NAND2_X1  g549(.A1(new_n727), .A2(new_n531), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n634), .A2(KEYINPUT103), .A3(G472), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT103), .B1(new_n634), .B2(G472), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n691), .B(new_n736), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n739), .A2(new_n705), .A3(new_n720), .ZN(new_n740));
  XOR2_X1   g554(.A(KEYINPUT105), .B(G125), .Z(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G27));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n696), .A2(new_n699), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n397), .A2(new_n744), .A3(new_n400), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n709), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n743), .B1(new_n747), .B2(new_n705), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n580), .A2(new_n581), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT32), .B1(new_n684), .B2(new_n531), .ZN(new_n750));
  OAI211_X1 g564(.A(KEYINPUT42), .B(new_n630), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n705), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT106), .B1(new_n752), .B2(new_n746), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT106), .ZN(new_n754));
  NOR4_X1   g568(.A1(new_n751), .A2(new_n745), .A3(new_n705), .A4(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n748), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT107), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n748), .B(KEYINPUT107), .C1(new_n753), .C2(new_n755), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G131), .ZN(G33));
  INV_X1    g575(.A(new_n747), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n671), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G134), .ZN(G36));
  AND2_X1   g578(.A1(new_n393), .A2(new_n395), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n765), .A2(KEYINPUT45), .ZN(new_n766));
  OAI21_X1  g580(.A(G469), .B1(new_n765), .B2(KEYINPUT45), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n768), .A2(new_n386), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n769), .A2(KEYINPUT46), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n385), .B1(new_n769), .B2(KEYINPUT46), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n400), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n676), .ZN(new_n774));
  INV_X1    g588(.A(new_n744), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n478), .A2(new_n645), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT43), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n636), .A2(new_n660), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n778), .A2(KEYINPUT44), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT44), .B1(new_n778), .B2(new_n779), .ZN(new_n781));
  NOR4_X1   g595(.A1(new_n774), .A2(new_n775), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n356), .ZN(G39));
  XNOR2_X1  g597(.A(new_n772), .B(KEYINPUT47), .ZN(new_n784));
  OR3_X1    g598(.A1(new_n775), .A2(new_n582), .A3(new_n630), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n784), .A2(new_n705), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(new_n402), .ZN(G42));
  NAND2_X1  g601(.A1(new_n712), .A2(new_n744), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n788), .B(new_n789), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n790), .A2(new_n189), .A3(new_n778), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n749), .A2(new_n750), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n630), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT48), .ZN(new_n794));
  INV_X1    g608(.A(G952), .ZN(new_n795));
  AND4_X1   g609(.A1(new_n189), .A2(new_n778), .A3(new_n630), .A4(new_n728), .ZN(new_n796));
  AOI211_X1 g610(.A(new_n795), .B(G953), .C1(new_n796), .C2(new_n721), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n477), .A2(new_n645), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n790), .A2(new_n189), .A3(new_n630), .A4(new_n690), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n794), .B(new_n797), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n784), .A2(KEYINPUT115), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n784), .A2(KEYINPUT115), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n711), .A2(new_n385), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n399), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT116), .Z(new_n806));
  NAND3_X1  g620(.A1(new_n802), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n796), .A2(new_n744), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(KEYINPUT51), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n778), .A2(new_n189), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n728), .A2(new_n630), .A3(new_n712), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n698), .A2(new_n699), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT50), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n800), .A2(new_n477), .A3(new_n645), .ZN(new_n816));
  INV_X1    g630(.A(new_n739), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n816), .B1(new_n817), .B2(new_n791), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT51), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n810), .B(new_n819), .C1(KEYINPUT118), .C2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n819), .A2(KEYINPUT118), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n808), .B1(new_n784), .B2(new_n805), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT51), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n801), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n798), .A2(KEYINPUT109), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n264), .A2(new_n266), .ZN(new_n828));
  OAI22_X1  g642(.A1(new_n798), .A2(KEYINPUT109), .B1(new_n477), .B2(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n638), .B(new_n637), .C1(new_n827), .C2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n632), .A3(new_n663), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n716), .A2(new_n713), .A3(new_n722), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n734), .A2(new_n833), .A3(KEYINPUT108), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT108), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n712), .A2(new_n582), .A3(new_n630), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n646), .B2(new_n652), .ZN(new_n837));
  AND4_X1   g651(.A1(new_n478), .A2(new_n718), .A3(new_n273), .A4(new_n721), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n730), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n731), .A2(KEYINPUT104), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n731), .A2(KEYINPUT104), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n835), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n832), .B1(new_n834), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n817), .A2(new_n706), .A3(new_n746), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n828), .A2(new_n651), .A3(new_n669), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n746), .A2(new_n847), .A3(new_n718), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n763), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n758), .A2(new_n850), .A3(new_n759), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n845), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n397), .A2(new_n400), .A3(new_n669), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n689), .A2(new_n855), .A3(new_n660), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n856), .B1(new_n841), .B2(new_n842), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n672), .B1(new_n670), .B2(new_n705), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n740), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n857), .A2(new_n859), .A3(KEYINPUT52), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT110), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n857), .A2(new_n859), .A3(KEYINPUT110), .A4(KEYINPUT52), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT52), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n689), .A2(new_n855), .A3(new_n660), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n866), .B1(new_n732), .B2(new_n733), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n706), .A2(new_n728), .A3(new_n721), .A4(new_n691), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n674), .A2(new_n707), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n865), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT111), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n857), .A2(new_n859), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT111), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(new_n873), .A3(new_n865), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT112), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n864), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n873), .B1(new_n872), .B2(new_n865), .ZN(new_n878));
  AOI211_X1 g692(.A(KEYINPUT111), .B(KEYINPUT52), .C1(new_n857), .C2(new_n859), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n862), .A2(new_n863), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT112), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n854), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n870), .A2(KEYINPUT113), .A3(new_n860), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT113), .B1(new_n870), .B2(new_n860), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n853), .B1(new_n852), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n883), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n831), .A2(new_n849), .A3(new_n853), .ZN(new_n890));
  OR3_X1    g704(.A1(new_n734), .A2(new_n833), .A3(KEYINPUT114), .ZN(new_n891));
  OAI21_X1  g705(.A(KEYINPUT114), .B1(new_n734), .B2(new_n833), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n890), .A2(new_n756), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n893), .B1(new_n882), .B2(new_n877), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT53), .B1(new_n852), .B2(new_n886), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n894), .A2(new_n895), .A3(KEYINPUT54), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n889), .A2(new_n896), .ZN(new_n897));
  AOI22_X1  g711(.A1(new_n825), .A2(new_n897), .B1(new_n795), .B2(new_n188), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n804), .B(KEYINPUT49), .Z(new_n899));
  NAND4_X1  g713(.A1(new_n698), .A2(new_n400), .A3(new_n480), .A4(new_n630), .ZN(new_n900));
  NOR4_X1   g714(.A1(new_n899), .A2(new_n689), .A3(new_n776), .A4(new_n900), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n898), .A2(new_n901), .ZN(G75));
  NOR2_X1   g716(.A1(new_n894), .A2(new_n895), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n903), .A2(new_n196), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(G210), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT56), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n524), .A2(new_n526), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(new_n520), .Z(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT55), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n905), .A2(new_n906), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n188), .A2(G952), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT56), .B1(new_n904), .B2(G210), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n915), .B1(new_n916), .B2(new_n910), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n905), .A2(new_n906), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n918), .A2(KEYINPUT119), .A3(new_n909), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n914), .B1(new_n917), .B2(new_n919), .ZN(G51));
  NAND2_X1  g734(.A1(new_n903), .A2(new_n888), .ZN(new_n921));
  OAI21_X1  g735(.A(KEYINPUT54), .B1(new_n894), .B2(new_n895), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g737(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n387), .B(new_n924), .ZN(new_n925));
  OAI22_X1  g739(.A1(new_n923), .A2(new_n925), .B1(new_n373), .B2(new_n384), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n904), .A2(new_n768), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n912), .B1(new_n926), .B2(new_n927), .ZN(G54));
  INV_X1    g742(.A(KEYINPUT121), .ZN(new_n929));
  AND2_X1   g743(.A1(KEYINPUT58), .A2(G475), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n904), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n929), .B1(new_n931), .B2(new_n473), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n912), .B1(new_n931), .B2(new_n473), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n904), .A2(KEYINPUT121), .A3(new_n459), .A4(new_n930), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(G60));
  NAND2_X1  g749(.A1(new_n639), .A2(new_n641), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n643), .B(KEYINPUT59), .Z(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g752(.A(KEYINPUT122), .B(new_n913), .C1(new_n923), .C2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n937), .B1(new_n889), .B2(new_n896), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n940), .A2(new_n639), .A3(new_n641), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n938), .B1(new_n921), .B2(new_n922), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(new_n912), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n939), .A2(new_n941), .A3(new_n944), .ZN(G63));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n946));
  NAND2_X1  g760(.A1(G217), .A2(G902), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT60), .ZN(new_n948));
  INV_X1    g762(.A(new_n893), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n880), .A2(KEYINPUT112), .A3(new_n881), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n876), .B1(new_n864), .B2(new_n875), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n852), .A2(new_n886), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n853), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n948), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n955), .A2(new_n628), .ZN(new_n956));
  INV_X1    g770(.A(new_n948), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n659), .B(new_n957), .C1(new_n894), .C2(new_n895), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n913), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n946), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n957), .B1(new_n894), .B2(new_n895), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT123), .ZN(new_n962));
  INV_X1    g776(.A(new_n628), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n962), .B1(new_n961), .B2(new_n963), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n958), .A2(KEYINPUT61), .A3(new_n913), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT124), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(KEYINPUT123), .B1(new_n955), .B2(new_n628), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n970));
  AND4_X1   g784(.A1(KEYINPUT124), .A2(new_n967), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n960), .B1(new_n968), .B2(new_n971), .ZN(G66));
  OAI21_X1  g786(.A(G953), .B1(new_n191), .B2(new_n504), .ZN(new_n973));
  OAI21_X1  g787(.A(KEYINPUT108), .B1(new_n734), .B2(new_n833), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n839), .A2(new_n835), .A3(new_n843), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n831), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n973), .B1(new_n976), .B2(G953), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n907), .B1(G898), .B2(new_n188), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n977), .B(new_n978), .ZN(G69));
  NOR2_X1   g793(.A1(new_n453), .A2(new_n454), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n575), .B(new_n980), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n786), .A2(new_n782), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n762), .B(new_n676), .C1(new_n827), .C2(new_n829), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n701), .A2(new_n859), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT62), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n984), .B(new_n985), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n982), .A2(new_n983), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n981), .B1(new_n987), .B2(G953), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT125), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n981), .B1(G900), .B2(G953), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n763), .A2(new_n859), .ZN(new_n991));
  INV_X1    g805(.A(new_n774), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n792), .A2(new_n630), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n993), .B1(new_n732), .B2(new_n733), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n991), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n982), .A2(new_n760), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n990), .B1(new_n996), .B2(G953), .ZN(new_n997));
  OAI21_X1  g811(.A(G953), .B1(new_n277), .B2(new_n667), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT126), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n988), .A2(new_n997), .ZN(new_n1001));
  OAI22_X1  g815(.A1(new_n989), .A2(new_n1000), .B1(new_n998), .B2(new_n1001), .ZN(G72));
  NAND2_X1  g816(.A1(G472), .A2(G902), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT63), .Z(new_n1004));
  OAI21_X1  g818(.A(new_n1004), .B1(new_n996), .B2(new_n845), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n1005), .A2(new_n547), .A3(new_n570), .A4(new_n554), .ZN(new_n1006));
  INV_X1    g820(.A(new_n679), .ZN(new_n1007));
  INV_X1    g821(.A(new_n1004), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1008), .B1(new_n987), .B2(new_n976), .ZN(new_n1009));
  OAI211_X1 g823(.A(new_n1006), .B(new_n913), .C1(new_n1007), .C2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n883), .A2(new_n887), .ZN(new_n1011));
  INV_X1    g825(.A(new_n576), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n570), .ZN(new_n1013));
  OR2_X1    g827(.A1(new_n1013), .A2(KEYINPUT127), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n544), .A2(new_n552), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1015), .B1(new_n1013), .B2(KEYINPUT127), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1008), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1010), .B1(new_n1011), .B2(new_n1017), .ZN(G57));
endmodule


