//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n805, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n977, new_n978, new_n979, new_n980, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016, new_n1017;
  AOI21_X1  g000(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n202));
  OAI21_X1  g001(.A(new_n202), .B1(G169gat), .B2(G176gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204));
  AOI22_X1  g003(.A1(new_n204), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT27), .B(G183gat), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  AOI21_X1  g006(.A(KEYINPUT28), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G183gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT27), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT27), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G183gat), .ZN(new_n212));
  AND4_X1   g011(.A1(KEYINPUT28), .A2(new_n210), .A3(new_n212), .A4(new_n207), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n203), .B(new_n205), .C1(new_n208), .C2(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(G183gat), .A2(G190gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT24), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT24), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n218), .A2(G183gat), .A3(G190gat), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n215), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n204), .A2(KEYINPUT23), .ZN(new_n222));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G169gat), .B2(G176gat), .ZN(new_n225));
  AND3_X1   g024(.A1(new_n222), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT25), .B1(new_n221), .B2(new_n226), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n222), .A2(KEYINPUT25), .A3(new_n225), .A4(new_n223), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n217), .A2(new_n219), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT65), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n215), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n228), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n214), .B1(new_n227), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G113gat), .ZN(new_n236));
  INV_X1    g035(.A(G120gat), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT1), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G134gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G127gat), .ZN(new_n240));
  INV_X1    g039(.A(G127gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G134gat), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n238), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n236), .A2(KEYINPUT66), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n236), .A2(KEYINPUT66), .ZN(new_n245));
  OAI21_X1  g044(.A(G120gat), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n238), .B1(new_n236), .B2(new_n237), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n240), .A2(new_n242), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n243), .A2(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n235), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G227gat), .A2(G233gat), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n251), .B(KEYINPUT64), .Z(new_n252));
  NAND3_X1  g051(.A1(new_n229), .A2(new_n232), .A3(new_n231), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(new_n226), .A3(KEYINPUT25), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT25), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n222), .A2(new_n223), .A3(new_n225), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n255), .B1(new_n256), .B2(new_n220), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n247), .A2(new_n248), .ZN(new_n259));
  XNOR2_X1  g058(.A(G127gat), .B(G134gat), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT66), .B(G113gat), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n238), .B(new_n260), .C1(new_n261), .C2(new_n237), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n258), .A2(new_n263), .A3(new_n214), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n250), .A2(new_n252), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT32), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT33), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(G15gat), .B(G43gat), .Z(new_n269));
  XNOR2_X1  g068(.A(G71gat), .B(G99gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n266), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n271), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n265), .B(KEYINPUT32), .C1(new_n267), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n252), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n235), .A2(new_n249), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n263), .B1(new_n258), .B2(new_n214), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT67), .B(KEYINPUT34), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT34), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n283), .A2(KEYINPUT67), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n276), .B(new_n285), .C1(new_n277), .C2(new_n278), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n275), .A2(new_n287), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n272), .A2(new_n274), .A3(new_n282), .A4(new_n286), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n252), .B1(new_n250), .B2(new_n264), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n286), .B(KEYINPUT68), .C1(new_n291), .C2(new_n280), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT68), .B1(new_n282), .B2(new_n286), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n275), .B(KEYINPUT69), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(new_n289), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT68), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n287), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n292), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT69), .B1(new_n299), .B2(new_n275), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  MUX2_X1   g100(.A(new_n290), .B(new_n301), .S(KEYINPUT36), .Z(new_n302));
  INV_X1    g101(.A(KEYINPUT82), .ZN(new_n303));
  INV_X1    g102(.A(G22gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(G228gat), .A2(G233gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT3), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT29), .ZN(new_n307));
  INV_X1    g106(.A(G197gat), .ZN(new_n308));
  INV_X1    g107(.A(G204gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G197gat), .A2(G204gat), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT22), .ZN(new_n312));
  NAND2_X1  g111(.A1(G211gat), .A2(G218gat), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n310), .A2(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G211gat), .ZN(new_n315));
  INV_X1    g114(.A(G218gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n317), .A2(new_n313), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n307), .B1(new_n314), .B2(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n314), .A2(new_n318), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n306), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G155gat), .A2(G162gat), .ZN(new_n322));
  OR2_X1    g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323));
  INV_X1    g122(.A(G141gat), .ZN(new_n324));
  INV_X1    g123(.A(G148gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G141gat), .A2(G148gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n322), .B(new_n323), .C1(new_n328), .C2(KEYINPUT2), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT75), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n323), .A2(new_n330), .A3(new_n322), .ZN(new_n331));
  AND2_X1   g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333));
  OAI21_X1  g132(.A(KEYINPUT75), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n326), .A2(new_n335), .A3(new_n327), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n331), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  AND2_X1   g136(.A1(G141gat), .A2(G148gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(G141gat), .A2(G148gat), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT74), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n322), .A2(KEYINPUT2), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n329), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n321), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G197gat), .B(G204gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n313), .A2(new_n312), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT70), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n348), .A3(new_n318), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n317), .A2(new_n348), .A3(new_n313), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n314), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n306), .B(new_n329), .C1(new_n337), .C2(new_n342), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n352), .B1(new_n353), .B2(new_n307), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n344), .B1(new_n354), .B2(KEYINPUT79), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT79), .ZN(new_n356));
  AOI211_X1 g155(.A(new_n356), .B(new_n352), .C1(new_n307), .C2(new_n353), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n305), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT80), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n360), .B(new_n305), .C1(new_n355), .C2(new_n357), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT29), .B1(new_n349), .B2(new_n351), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n343), .B1(new_n363), .B2(KEYINPUT3), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT81), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n353), .A2(new_n307), .ZN(new_n367));
  INV_X1    g166(.A(new_n352), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g168(.A(KEYINPUT81), .B(new_n343), .C1(new_n363), .C2(KEYINPUT3), .ZN(new_n370));
  INV_X1    g169(.A(new_n305), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n366), .A2(new_n369), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n304), .B1(new_n362), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n372), .ZN(new_n374));
  AOI211_X1 g173(.A(G22gat), .B(new_n374), .C1(new_n359), .C2(new_n361), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n303), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n369), .A2(new_n356), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n354), .A2(KEYINPUT79), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n377), .A2(new_n378), .A3(new_n344), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n360), .B1(new_n379), .B2(new_n305), .ZN(new_n380));
  INV_X1    g179(.A(new_n361), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n372), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G22gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n362), .A2(new_n304), .A3(new_n372), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(KEYINPUT82), .A3(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(G78gat), .B(G106gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT31), .B(G50gat), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n386), .B(new_n387), .Z(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n376), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n383), .A2(KEYINPUT82), .A3(new_n384), .A4(new_n388), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(G8gat), .B(G36gat), .Z(new_n393));
  XNOR2_X1  g192(.A(new_n393), .B(KEYINPUT72), .ZN(new_n394));
  XNOR2_X1  g193(.A(G64gat), .B(G92gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(G226gat), .ZN(new_n397));
  INV_X1    g196(.A(G233gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n399), .A2(KEYINPUT29), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT71), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n235), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n258), .A2(KEYINPUT71), .A3(new_n214), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n401), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n399), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n235), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n352), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n235), .A2(new_n400), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n403), .A2(new_n404), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n368), .B(new_n409), .C1(new_n410), .C2(new_n406), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n396), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n408), .A2(new_n411), .A3(new_n396), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n408), .A2(new_n411), .A3(KEYINPUT30), .A4(new_n396), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n416), .A2(KEYINPUT73), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(KEYINPUT73), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n415), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n421), .B1(new_n343), .B2(new_n263), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n328), .A2(KEYINPUT74), .B1(KEYINPUT2), .B2(new_n322), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n423), .A2(new_n331), .A3(new_n336), .A4(new_n334), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n424), .A2(new_n249), .A3(KEYINPUT4), .A4(new_n329), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n249), .B1(new_n343), .B2(KEYINPUT3), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n427), .A2(KEYINPUT76), .A3(new_n353), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT76), .B1(new_n427), .B2(new_n353), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n420), .B(new_n426), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT77), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT78), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n424), .A2(new_n249), .A3(new_n329), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n343), .A2(new_n263), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n420), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n432), .B1(new_n437), .B2(KEYINPUT5), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT5), .ZN(new_n439));
  AOI211_X1 g238(.A(KEYINPUT78), .B(new_n439), .C1(new_n435), .C2(new_n436), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n343), .A2(KEYINPUT3), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(new_n353), .A3(new_n263), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT76), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n427), .A2(KEYINPUT76), .A3(new_n353), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT77), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n420), .A4(new_n426), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n431), .A2(new_n441), .A3(new_n449), .ZN(new_n450));
  OR2_X1    g249(.A1(new_n430), .A2(KEYINPUT5), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(G1gat), .B(G29gat), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n453), .B(KEYINPUT0), .ZN(new_n454));
  XNOR2_X1  g253(.A(G57gat), .B(G85gat), .ZN(new_n455));
  XOR2_X1   g254(.A(new_n454), .B(new_n455), .Z(new_n456));
  AOI21_X1  g255(.A(KEYINPUT6), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n456), .B1(new_n450), .B2(new_n451), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n458), .A2(KEYINPUT6), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n419), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n302), .B1(new_n392), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n413), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT37), .ZN(new_n465));
  INV_X1    g264(.A(new_n410), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n466), .A2(new_n399), .B1(new_n400), .B2(new_n235), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n465), .B1(new_n467), .B2(new_n352), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n368), .B1(new_n405), .B2(new_n407), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT38), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n408), .A2(new_n465), .A3(new_n411), .ZN(new_n471));
  INV_X1    g270(.A(new_n396), .ZN(new_n472));
  AND2_X1   g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n464), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT84), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n450), .A2(new_n475), .A3(new_n451), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n475), .B1(new_n450), .B2(new_n451), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n476), .A2(new_n477), .A3(new_n456), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n450), .A2(new_n451), .ZN(new_n480));
  INV_X1    g279(.A(new_n456), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n461), .B(new_n474), .C1(new_n478), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT85), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n480), .A2(KEYINPUT84), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n450), .A2(new_n475), .A3(new_n451), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(new_n481), .A3(new_n486), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n487), .A2(new_n457), .B1(KEYINPUT6), .B2(new_n458), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT85), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(new_n489), .A3(new_n474), .ZN(new_n490));
  INV_X1    g289(.A(new_n473), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n465), .B1(new_n408), .B2(new_n411), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT38), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n484), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n447), .A2(new_n426), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n436), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n433), .A2(new_n434), .A3(new_n420), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(KEYINPUT39), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n456), .B1(new_n496), .B2(KEYINPUT39), .ZN(new_n500));
  OAI22_X1  g299(.A1(new_n499), .A2(new_n500), .B1(KEYINPUT83), .B2(KEYINPUT40), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n496), .A2(KEYINPUT39), .ZN(new_n502));
  NOR2_X1   g301(.A1(KEYINPUT83), .A2(KEYINPUT40), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n502), .A2(new_n456), .A3(new_n503), .A4(new_n498), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(KEYINPUT83), .A2(KEYINPUT40), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n419), .A3(new_n506), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n391), .B(new_n390), .C1(new_n507), .C2(new_n478), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n463), .B1(new_n494), .B2(new_n509), .ZN(new_n510));
  NOR3_X1   g309(.A1(new_n419), .A2(KEYINPUT35), .A3(new_n290), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n511), .A2(new_n391), .A3(new_n390), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n512), .A2(new_n488), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n390), .A2(new_n391), .A3(new_n301), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT86), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT86), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n390), .A2(new_n301), .A3(new_n516), .A4(new_n391), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n515), .A2(new_n462), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n513), .B1(new_n518), .B2(KEYINPUT35), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n510), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(G113gat), .B(G141gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(G197gat), .ZN(new_n522));
  XOR2_X1   g321(.A(KEYINPUT11), .B(G169gat), .Z(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  XOR2_X1   g323(.A(new_n524), .B(KEYINPUT12), .Z(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n526), .A2(G1gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT16), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n526), .B1(new_n528), .B2(G1gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT88), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n531), .B1(new_n526), .B2(G1gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n530), .A2(G8gat), .A3(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(G8gat), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n527), .B(new_n529), .C1(new_n531), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT89), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n533), .A2(KEYINPUT89), .A3(new_n535), .ZN(new_n539));
  NOR2_X1   g338(.A1(G29gat), .A2(G36gat), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT14), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G29gat), .A2(G36gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G43gat), .B(G50gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(KEYINPUT15), .A3(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n545), .A2(KEYINPUT15), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(KEYINPUT15), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n543), .B(KEYINPUT87), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n547), .A2(new_n542), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n538), .A2(new_n539), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT91), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n538), .A2(KEYINPUT91), .A3(new_n539), .A4(new_n552), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n533), .A2(KEYINPUT89), .A3(new_n535), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT89), .B1(new_n533), .B2(new_n535), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n551), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n555), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT90), .B(KEYINPUT13), .ZN(new_n561));
  NAND2_X1  g360(.A1(G229gat), .A2(G233gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n536), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n551), .A2(KEYINPUT17), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT17), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n566), .B1(new_n546), .B2(new_n550), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n564), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  AND3_X1   g367(.A1(new_n559), .A2(new_n568), .A3(new_n562), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n560), .A2(new_n563), .B1(new_n569), .B2(KEYINPUT18), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT92), .ZN(new_n571));
  OAI22_X1  g370(.A1(new_n570), .A2(new_n571), .B1(KEYINPUT18), .B2(new_n569), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n560), .A2(new_n563), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n569), .A2(KEYINPUT18), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n573), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n525), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n559), .A2(new_n568), .A3(new_n562), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT18), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n525), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n570), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT93), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n570), .A2(KEYINPUT93), .A3(new_n579), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n576), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n520), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT94), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT94), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n520), .A2(new_n588), .A3(new_n585), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT21), .ZN(new_n591));
  XNOR2_X1  g390(.A(G57gat), .B(G64gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(G71gat), .ZN(new_n594));
  INV_X1    g393(.A(G78gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G71gat), .A2(G78gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT9), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n593), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n597), .B(new_n596), .C1(new_n592), .C2(new_n599), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT95), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n601), .A2(new_n602), .A3(KEYINPUT95), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n538), .B(new_n539), .C1(new_n591), .C2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT97), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n591), .ZN(new_n610));
  XNOR2_X1  g409(.A(G127gat), .B(G155gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n610), .B(new_n611), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n609), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT96), .ZN(new_n615));
  XOR2_X1   g414(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G183gat), .B(G211gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n613), .B(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G134gat), .B(G162gat), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(KEYINPUT98), .B(KEYINPUT7), .Z(new_n626));
  INV_X1    g425(.A(G85gat), .ZN(new_n627));
  INV_X1    g426(.A(G92gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT98), .B(KEYINPUT7), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n631), .B1(new_n627), .B2(new_n628), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G99gat), .B(G106gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n627), .A2(KEYINPUT99), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT99), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(G85gat), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n635), .A2(new_n637), .A3(new_n628), .ZN(new_n638));
  NAND2_X1  g437(.A1(G99gat), .A2(G106gat), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT8), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  AND4_X1   g441(.A1(KEYINPUT100), .A2(new_n633), .A3(new_n634), .A4(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n641), .B1(new_n630), .B2(new_n632), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT100), .B1(new_n644), .B2(new_n634), .ZN(new_n645));
  OAI21_X1  g444(.A(KEYINPUT101), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT100), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n633), .A2(new_n642), .ZN(new_n648));
  INV_X1    g447(.A(new_n634), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT101), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n644), .A2(KEYINPUT100), .A3(new_n634), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n648), .A2(new_n649), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n646), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n655), .B1(new_n567), .B2(new_n565), .ZN(new_n656));
  NAND3_X1  g455(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(G190gat), .B(G218gat), .Z(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n655), .A2(new_n552), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n660), .B1(new_n658), .B2(new_n661), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n625), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n664), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n666), .A2(new_n624), .A3(new_n662), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n621), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n607), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT10), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n603), .B1(new_n648), .B2(new_n649), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n673), .B1(new_n643), .B2(new_n645), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT102), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n673), .B(KEYINPUT102), .C1(new_n643), .C2(new_n645), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n671), .A2(new_n672), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n605), .A2(KEYINPUT10), .A3(new_n606), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n655), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(G230gat), .A2(G233gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT103), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n655), .A2(new_n607), .B1(new_n676), .B2(new_n677), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n688), .A2(new_n686), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(G120gat), .B(G148gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(G176gat), .B(G204gat), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n692), .B(new_n693), .Z(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n685), .B1(new_n679), .B2(new_n682), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(new_n689), .ZN(new_n698));
  AOI21_X1  g497(.A(KEYINPUT104), .B1(new_n698), .B2(new_n694), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n700));
  NOR4_X1   g499(.A1(new_n697), .A2(new_n689), .A3(new_n700), .A4(new_n695), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n696), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n670), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n460), .A2(new_n461), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n460), .A2(KEYINPUT105), .A3(new_n461), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n590), .A2(new_n705), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g512(.A(new_n704), .B1(new_n587), .B2(new_n589), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT106), .B(KEYINPUT16), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(G8gat), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n714), .A2(new_n419), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT42), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n714), .A2(KEYINPUT42), .A3(new_n419), .A4(new_n716), .ZN(new_n720));
  INV_X1    g519(.A(new_n589), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n588), .B1(new_n520), .B2(new_n585), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n419), .B(new_n705), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n723), .A2(new_n724), .A3(G8gat), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n723), .B2(G8gat), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n719), .B(new_n720), .C1(new_n725), .C2(new_n726), .ZN(G1325gat));
  INV_X1    g526(.A(new_n290), .ZN(new_n728));
  AOI21_X1  g527(.A(G15gat), .B1(new_n714), .B2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n302), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G15gat), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT108), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n729), .B1(new_n714), .B2(new_n732), .ZN(G1326gat));
  INV_X1    g532(.A(new_n392), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n714), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(KEYINPUT43), .B(G22gat), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1327gat));
  NOR3_X1   g536(.A1(new_n702), .A2(new_n620), .A3(new_n668), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n590), .A2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT45), .ZN(new_n740));
  INV_X1    g539(.A(G29gat), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n711), .A2(new_n741), .ZN(new_n742));
  OR3_X1    g541(.A1(new_n739), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n669), .B1(new_n510), .B2(new_n519), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI211_X1 g545(.A(KEYINPUT44), .B(new_n669), .C1(new_n510), .C2(new_n519), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n620), .B(KEYINPUT109), .Z(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n585), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n749), .A2(new_n750), .A3(new_n702), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n746), .A2(new_n747), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G29gat), .B1(new_n752), .B2(new_n710), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n740), .B1(new_n739), .B2(new_n742), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n743), .A2(new_n753), .A3(new_n754), .ZN(G1328gat));
  INV_X1    g554(.A(new_n419), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n756), .A2(G36gat), .ZN(new_n757));
  OR3_X1    g556(.A1(new_n739), .A2(KEYINPUT46), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(G36gat), .B1(new_n752), .B2(new_n756), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT46), .B1(new_n739), .B2(new_n757), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(G1329gat));
  NOR2_X1   g560(.A1(new_n290), .A2(G43gat), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n590), .A2(new_n738), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n764));
  OAI21_X1  g563(.A(G43gat), .B1(new_n752), .B2(new_n302), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n764), .B1(new_n763), .B2(new_n765), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n766), .A2(new_n767), .ZN(G1330gat));
  NOR2_X1   g567(.A1(new_n392), .A2(G50gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n590), .A2(new_n738), .A3(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT48), .ZN(new_n771));
  OAI21_X1  g570(.A(G50gat), .B1(new_n752), .B2(new_n392), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n771), .B1(new_n770), .B2(new_n772), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(G1331gat));
  NOR4_X1   g574(.A1(new_n703), .A2(new_n621), .A3(new_n669), .A4(new_n585), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT111), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(new_n520), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT112), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n777), .A2(new_n520), .A3(KEYINPUT112), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(new_n710), .ZN(new_n783));
  XOR2_X1   g582(.A(new_n783), .B(G57gat), .Z(G1332gat));
  XNOR2_X1  g583(.A(new_n419), .B(KEYINPUT113), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT114), .B1(new_n782), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n780), .A2(new_n789), .A3(new_n781), .A4(new_n786), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT49), .ZN(new_n792));
  INV_X1    g591(.A(G64gat), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n788), .A2(new_n792), .A3(new_n793), .A4(new_n790), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(G1333gat));
  OAI21_X1  g596(.A(G71gat), .B1(new_n782), .B2(new_n302), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n780), .A2(new_n594), .A3(new_n728), .A4(new_n781), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n798), .A2(KEYINPUT50), .A3(new_n799), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(G1334gat));
  NOR2_X1   g603(.A1(new_n782), .A2(new_n392), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(new_n595), .ZN(G1335gat));
  NOR2_X1   g605(.A1(new_n620), .A2(new_n585), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n520), .A2(KEYINPUT51), .A3(new_n669), .A4(new_n807), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n669), .B(new_n807), .C1(new_n510), .C2(new_n519), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n703), .B1(new_n808), .B2(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n635), .A2(new_n637), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n813), .A3(new_n711), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n703), .A2(new_n585), .A3(new_n620), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n746), .A2(new_n747), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n746), .A2(KEYINPUT115), .A3(new_n747), .A4(new_n815), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n818), .A2(new_n711), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n814), .B1(new_n820), .B2(new_n813), .ZN(G1336gat));
  XNOR2_X1  g620(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n785), .A2(G92gat), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n812), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(G92gat), .B1(new_n816), .B2(new_n785), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT117), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n809), .A2(new_n810), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n809), .A2(new_n810), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n702), .B(new_n823), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n822), .ZN(new_n830));
  AND4_X1   g629(.A1(KEYINPUT117), .A2(new_n825), .A3(new_n829), .A4(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(new_n823), .ZN(new_n832));
  AOI211_X1 g631(.A(new_n703), .B(new_n832), .C1(new_n808), .C2(new_n811), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n419), .A3(new_n819), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n833), .B1(new_n834), .B2(G92gat), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT52), .ZN(new_n836));
  OAI22_X1  g635(.A1(new_n826), .A2(new_n831), .B1(new_n835), .B2(new_n836), .ZN(G1337gat));
  INV_X1    g636(.A(G99gat), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n812), .A2(new_n838), .A3(new_n728), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n818), .A2(new_n730), .A3(new_n819), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(new_n838), .ZN(G1338gat));
  NOR2_X1   g640(.A1(new_n392), .A2(G106gat), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n812), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n844));
  OAI21_X1  g643(.A(G106gat), .B1(new_n816), .B2(new_n392), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n818), .A2(new_n734), .A3(new_n819), .ZN(new_n847));
  AOI22_X1  g646(.A1(new_n847), .A2(G106gat), .B1(new_n812), .B2(new_n842), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n846), .B1(new_n848), .B2(new_n844), .ZN(G1339gat));
  NAND3_X1  g648(.A1(new_n670), .A2(new_n750), .A3(new_n703), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n559), .A2(new_n568), .ZN(new_n851));
  OAI22_X1  g650(.A1(new_n560), .A2(new_n563), .B1(new_n562), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n524), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n702), .A2(new_n584), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n700), .B1(new_n691), .B2(new_n695), .ZN(new_n855));
  INV_X1    g654(.A(new_n701), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT118), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n681), .B1(new_n688), .B2(new_n672), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT54), .B1(new_n859), .B2(new_n685), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n683), .A2(new_n686), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n859), .A2(new_n685), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n687), .A2(new_n863), .A3(KEYINPUT118), .A4(KEYINPUT54), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n694), .B1(new_n697), .B2(new_n865), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n862), .A2(KEYINPUT55), .A3(new_n864), .A4(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n857), .A2(new_n867), .A3(new_n585), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n683), .A2(new_n865), .A3(new_n686), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n695), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n687), .A2(new_n863), .A3(KEYINPUT54), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n858), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(KEYINPUT55), .B1(new_n872), .B2(new_n864), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n854), .B1(new_n868), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n857), .A2(new_n867), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n665), .A2(new_n584), .A3(new_n667), .A4(new_n853), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  AOI22_X1  g677(.A1(new_n874), .A2(new_n668), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n850), .B1(new_n879), .B2(new_n749), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n734), .A2(new_n290), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n880), .A2(new_n711), .A3(new_n785), .A4(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(G113gat), .B1(new_n882), .B2(new_n750), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n880), .A2(new_n711), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n515), .A2(new_n517), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n785), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n585), .A2(new_n261), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n883), .B1(new_n887), .B2(new_n888), .ZN(G1340gat));
  NOR3_X1   g688(.A1(new_n882), .A2(new_n237), .A3(new_n703), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n886), .A2(new_n702), .A3(new_n785), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n890), .B1(new_n891), .B2(new_n237), .ZN(G1341gat));
  OAI21_X1  g691(.A(G127gat), .B1(new_n882), .B2(new_n748), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n620), .A2(new_n241), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n887), .B2(new_n894), .ZN(G1342gat));
  NAND4_X1  g694(.A1(new_n886), .A2(new_n239), .A3(new_n756), .A4(new_n669), .ZN(new_n896));
  OR2_X1    g695(.A1(new_n896), .A2(KEYINPUT56), .ZN(new_n897));
  OAI21_X1  g696(.A(G134gat), .B1(new_n882), .B2(new_n668), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(KEYINPUT56), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(G1343gat));
  INV_X1    g699(.A(KEYINPUT57), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n880), .A2(new_n901), .A3(new_n734), .ZN(new_n902));
  INV_X1    g701(.A(new_n785), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n710), .A2(new_n730), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n862), .A2(new_n864), .A3(new_n866), .ZN(new_n905));
  XOR2_X1   g704(.A(KEYINPUT119), .B(KEYINPUT55), .Z(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n907), .A2(new_n585), .A3(new_n857), .A4(new_n867), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n669), .B1(new_n908), .B2(new_n854), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n875), .A2(new_n873), .A3(new_n877), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n621), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n392), .B1(new_n911), .B2(new_n850), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n902), .B(new_n904), .C1(new_n901), .C2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT121), .B1(new_n913), .B2(new_n750), .ZN(new_n914));
  INV_X1    g713(.A(new_n904), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n911), .A2(new_n850), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n734), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n915), .B1(new_n917), .B2(KEYINPUT57), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT121), .ZN(new_n919));
  NAND4_X1  g718(.A1(new_n918), .A2(new_n919), .A3(new_n585), .A4(new_n902), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n914), .A2(G141gat), .A3(new_n920), .ZN(new_n921));
  XOR2_X1   g720(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n922));
  NOR2_X1   g721(.A1(new_n730), .A2(new_n392), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n884), .A2(new_n785), .A3(new_n923), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n750), .A2(G141gat), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n921), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(G141gat), .B1(new_n913), .B2(new_n750), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n924), .A2(new_n925), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT58), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n927), .A2(new_n931), .ZN(G1344gat));
  NAND3_X1  g731(.A1(new_n924), .A2(new_n325), .A3(new_n702), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT59), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n392), .A2(KEYINPUT57), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(KEYINPUT122), .B1(new_n909), .B2(new_n910), .ZN(new_n937));
  INV_X1    g736(.A(new_n906), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n938), .B1(new_n872), .B2(new_n864), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n854), .B1(new_n868), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(new_n668), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n878), .A2(new_n876), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n937), .A2(new_n944), .A3(new_n621), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n936), .B1(new_n945), .B2(new_n850), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n901), .B1(new_n880), .B2(new_n734), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n948), .A2(new_n702), .A3(new_n904), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n934), .B1(new_n949), .B2(G148gat), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n913), .A2(new_n703), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n951), .A2(KEYINPUT59), .A3(new_n325), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n933), .B1(new_n950), .B2(new_n952), .ZN(G1345gat));
  INV_X1    g752(.A(G155gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n924), .A2(new_n954), .A3(new_n620), .ZN(new_n955));
  OAI21_X1  g754(.A(G155gat), .B1(new_n913), .B2(new_n748), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(G1346gat));
  OAI21_X1  g756(.A(G162gat), .B1(new_n913), .B2(new_n668), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n668), .A2(G162gat), .A3(new_n419), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n884), .A2(new_n923), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(KEYINPUT123), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT123), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n958), .A2(new_n960), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n964), .ZN(G1347gat));
  NOR2_X1   g764(.A1(new_n711), .A2(new_n756), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n880), .A2(new_n881), .A3(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(G169gat), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n967), .A2(new_n968), .A3(new_n750), .ZN(new_n969));
  AND4_X1   g768(.A1(new_n885), .A2(new_n880), .A3(new_n710), .A4(new_n903), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(new_n585), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n969), .B1(new_n968), .B2(new_n971), .ZN(G1348gat));
  INV_X1    g771(.A(G176gat), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n970), .A2(new_n973), .A3(new_n702), .ZN(new_n974));
  OAI21_X1  g773(.A(G176gat), .B1(new_n967), .B2(new_n703), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(G1349gat));
  NAND3_X1  g775(.A1(new_n970), .A2(new_n206), .A3(new_n620), .ZN(new_n977));
  OAI21_X1  g776(.A(G183gat), .B1(new_n967), .B2(new_n748), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n980));
  XOR2_X1   g779(.A(new_n979), .B(new_n980), .Z(G1350gat));
  NAND3_X1  g780(.A1(new_n970), .A2(new_n207), .A3(new_n669), .ZN(new_n982));
  OAI21_X1  g781(.A(G190gat), .B1(new_n967), .B2(new_n668), .ZN(new_n983));
  AND2_X1   g782(.A1(new_n983), .A2(KEYINPUT61), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n983), .A2(KEYINPUT61), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(G1351gat));
  NAND2_X1  g785(.A1(new_n923), .A2(new_n903), .ZN(new_n987));
  INV_X1    g786(.A(new_n987), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n880), .A2(new_n710), .A3(new_n988), .ZN(new_n989));
  INV_X1    g788(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g789(.A(G197gat), .B1(new_n990), .B2(new_n585), .ZN(new_n991));
  INV_X1    g790(.A(KEYINPUT125), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n992), .B1(new_n966), .B2(new_n302), .ZN(new_n993));
  NOR4_X1   g792(.A1(new_n711), .A2(KEYINPUT125), .A3(new_n756), .A4(new_n730), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n995), .A2(new_n308), .A3(new_n750), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n991), .B1(new_n948), .B2(new_n996), .ZN(G1352gat));
  NOR2_X1   g796(.A1(new_n703), .A2(G204gat), .ZN(new_n998));
  NAND4_X1  g797(.A1(new_n880), .A2(new_n710), .A3(new_n988), .A4(new_n998), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT62), .ZN(new_n1000));
  XNOR2_X1  g799(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  NOR4_X1   g800(.A1(new_n946), .A2(new_n947), .A3(new_n703), .A4(new_n995), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n1001), .B1(new_n1002), .B2(new_n309), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT126), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g804(.A(KEYINPUT126), .B(new_n1001), .C1(new_n1002), .C2(new_n309), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1005), .A2(new_n1006), .ZN(G1353gat));
  NAND3_X1  g806(.A1(new_n990), .A2(new_n315), .A3(new_n620), .ZN(new_n1008));
  NOR4_X1   g807(.A1(new_n711), .A2(new_n756), .A3(new_n730), .A4(new_n621), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n948), .A2(new_n1009), .ZN(new_n1010));
  AND3_X1   g809(.A1(new_n1010), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1011));
  AOI21_X1  g810(.A(KEYINPUT63), .B1(new_n1010), .B2(G211gat), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1008), .B1(new_n1011), .B2(new_n1012), .ZN(G1354gat));
  AOI21_X1  g812(.A(G218gat), .B1(new_n990), .B2(new_n669), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n669), .A2(G218gat), .ZN(new_n1015));
  XNOR2_X1  g814(.A(new_n1015), .B(KEYINPUT127), .ZN(new_n1016));
  NOR2_X1   g815(.A1(new_n995), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g816(.A(new_n1014), .B1(new_n948), .B2(new_n1017), .ZN(G1355gat));
endmodule


