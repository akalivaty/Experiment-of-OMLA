//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n557,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  OR2_X1    g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n465), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n469), .B1(new_n463), .B2(new_n464), .ZN(new_n470));
  AND2_X1   g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n463), .A2(new_n464), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  INV_X1    g051(.A(G124), .ZN(new_n477));
  NOR2_X1   g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI21_X1  g053(.A(G2104), .B1(new_n466), .B2(G112), .ZN(new_n479));
  OAI22_X1  g054(.A1(new_n476), .A2(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n480), .B1(G136), .B2(new_n465), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT68), .Z(G162));
  INV_X1    g057(.A(new_n467), .ZN(new_n483));
  INV_X1    g058(.A(G102), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(G114), .A2(G2104), .ZN(new_n486));
  XOR2_X1   g061(.A(KEYINPUT3), .B(G2104), .Z(new_n487));
  INV_X1    g062(.A(G126), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n485), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n475), .A2(G138), .A3(new_n466), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n465), .A2(new_n493), .A3(G138), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT69), .B1(new_n498), .B2(KEYINPUT6), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(new_n501), .A3(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n498), .A2(KEYINPUT6), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT5), .B(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G88), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n500), .B1(new_n501), .B2(G651), .ZN(new_n509));
  NOR3_X1   g084(.A1(new_n498), .A2(KEYINPUT69), .A3(KEYINPUT6), .ZN(new_n510));
  OAI211_X1 g085(.A(G543), .B(new_n504), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n514), .A2(new_n498), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n508), .A2(new_n513), .A3(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT5), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G543), .ZN(new_n521));
  AND3_X1   g096(.A1(new_n519), .A2(new_n521), .A3(KEYINPUT70), .ZN(new_n522));
  AOI21_X1  g097(.A(KEYINPUT70), .B1(new_n519), .B2(new_n521), .ZN(new_n523));
  OAI211_X1 g098(.A(G63), .B(G651), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n503), .A2(G89), .A3(new_n504), .A4(new_n505), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n511), .A2(KEYINPUT71), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n503), .A2(new_n530), .A3(G543), .A4(new_n504), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n529), .A2(G51), .A3(new_n531), .ZN(new_n532));
  AND3_X1   g107(.A1(new_n526), .A2(new_n528), .A3(new_n532), .ZN(G168));
  INV_X1    g108(.A(G64), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n519), .A2(new_n521), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT70), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n519), .A2(new_n521), .A3(KEYINPUT70), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n534), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AND2_X1   g114(.A1(G77), .A2(G543), .ZN(new_n540));
  OAI21_X1  g115(.A(G651), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n529), .A2(G52), .A3(new_n531), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n507), .A2(G90), .ZN(new_n543));
  AND3_X1   g118(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(G171));
  NAND2_X1  g119(.A1(new_n537), .A2(new_n538), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n545), .A2(G56), .ZN(new_n546));
  AND2_X1   g121(.A1(G68), .A2(G543), .ZN(new_n547));
  OAI21_X1  g122(.A(G651), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n529), .A2(G43), .A3(new_n531), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n507), .A2(G81), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n549), .A2(KEYINPUT72), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g126(.A(KEYINPUT72), .B1(new_n549), .B2(new_n550), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n548), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(new_n557));
  XOR2_X1   g132(.A(new_n557), .B(KEYINPUT73), .Z(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(G188));
  NAND3_X1  g136(.A1(new_n512), .A2(KEYINPUT9), .A3(G53), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n507), .A2(G91), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n505), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(new_n498), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n511), .B2(new_n567), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n562), .A2(new_n563), .A3(new_n565), .A4(new_n568), .ZN(G299));
  NAND3_X1  g144(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(G301));
  NAND3_X1  g145(.A1(new_n526), .A2(new_n528), .A3(new_n532), .ZN(G286));
  OAI21_X1  g146(.A(G651), .B1(new_n545), .B2(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n507), .A2(G87), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n512), .A2(G49), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  NAND2_X1  g150(.A1(new_n507), .A2(G86), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n512), .A2(G48), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n505), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n578));
  OR2_X1    g153(.A1(new_n578), .A2(new_n498), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(G305));
  AOI22_X1  g155(.A1(new_n545), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n581), .A2(new_n498), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n529), .A2(new_n531), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G47), .ZN(new_n584));
  XNOR2_X1  g159(.A(KEYINPUT74), .B(G85), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n507), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n582), .A2(new_n584), .A3(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n507), .A2(KEYINPUT10), .A3(G92), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT10), .ZN(new_n590));
  INV_X1    g165(.A(G92), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n506), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n535), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n589), .A2(new_n592), .B1(G651), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n583), .A2(G54), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n588), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n588), .B1(new_n599), .B2(G868), .ZN(G321));
  NAND2_X1  g176(.A1(G286), .A2(G868), .ZN(new_n602));
  XOR2_X1   g177(.A(G299), .B(KEYINPUT75), .Z(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G868), .ZN(G297));
  OAI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(G868), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND3_X1  g182(.A1(new_n596), .A2(new_n597), .A3(new_n606), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT76), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  AND2_X1   g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n554), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(KEYINPUT77), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(KEYINPUT77), .B2(new_n611), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n475), .A2(new_n467), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT12), .Z(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT13), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2100), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n465), .A2(G135), .ZN(new_n620));
  NOR2_X1   g195(.A1(G99), .A2(G2105), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(new_n466), .B2(G111), .ZN(new_n622));
  INV_X1    g197(.A(G123), .ZN(new_n623));
  OAI221_X1 g198(.A(new_n620), .B1(new_n621), .B2(new_n622), .C1(new_n623), .C2(new_n476), .ZN(new_n624));
  INV_X1    g199(.A(G2096), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n619), .A2(new_n626), .ZN(G156));
  XNOR2_X1  g202(.A(G1341), .B(G1348), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2435), .ZN(new_n632));
  XOR2_X1   g207(.A(G2427), .B(G2438), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(KEYINPUT14), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(KEYINPUT80), .ZN(new_n636));
  INV_X1    g211(.A(G2451), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT80), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n634), .A2(new_n638), .A3(KEYINPUT14), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n637), .B1(new_n636), .B2(new_n639), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n630), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n636), .A2(new_n639), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(G2451), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n645), .A2(G2454), .A3(new_n640), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT79), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n643), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n649), .B1(new_n643), .B2(new_n646), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  NOR3_X1   g229(.A1(new_n651), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n643), .A2(new_n646), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(new_n648), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n653), .B1(new_n657), .B2(new_n650), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n629), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n654), .B1(new_n651), .B2(new_n652), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n657), .A2(new_n653), .A3(new_n650), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n660), .A2(new_n661), .A3(new_n628), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n659), .A2(G14), .A3(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(G401));
  XNOR2_X1  g239(.A(G2072), .B(G2078), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT81), .ZN(new_n666));
  XOR2_X1   g241(.A(G2084), .B(G2090), .Z(new_n667));
  XOR2_X1   g242(.A(G2067), .B(G2678), .Z(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n666), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT18), .Z(new_n671));
  INV_X1    g246(.A(KEYINPUT82), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n666), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT17), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n674), .A2(new_n667), .A3(new_n668), .ZN(new_n675));
  INV_X1    g250(.A(new_n667), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(new_n674), .B2(new_n668), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n666), .A2(new_n669), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n671), .B(new_n675), .C1(new_n677), .C2(new_n678), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n679), .A2(G2100), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT83), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(G2100), .ZN(new_n682));
  AND3_X1   g257(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n681), .B1(new_n680), .B2(new_n682), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n625), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n680), .A2(new_n682), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(KEYINPUT83), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n687), .A2(G2096), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G227));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  XOR2_X1   g268(.A(G1956), .B(G2474), .Z(new_n694));
  XOR2_X1   g269(.A(G1961), .B(G1966), .Z(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n693), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n694), .A2(new_n695), .ZN(new_n699));
  AOI22_X1  g274(.A1(new_n697), .A2(KEYINPUT20), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n699), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n701), .A2(new_n693), .A3(new_n696), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n700), .B(new_n702), .C1(KEYINPUT20), .C2(new_n697), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT84), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n703), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1991), .B(G1996), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(G1981), .B(G1986), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(G229));
  OR2_X1    g285(.A1(G29), .A2(G32), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n467), .A2(G105), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT92), .Z(new_n713));
  INV_X1    g288(.A(new_n476), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n714), .A2(G129), .B1(G141), .B2(new_n465), .ZN(new_n715));
  NAND3_X1  g290(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT26), .Z(new_n717));
  NAND3_X1  g292(.A1(new_n713), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n711), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT27), .B(G1996), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n719), .A2(G26), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n714), .A2(G128), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n465), .A2(G140), .ZN(new_n725));
  OR2_X1    g300(.A1(G104), .A2(G2105), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n726), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n723), .B1(new_n729), .B2(new_n719), .ZN(new_n730));
  MUX2_X1   g305(.A(new_n723), .B(new_n730), .S(KEYINPUT28), .Z(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT88), .B(G2067), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G2084), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G34), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(new_n719), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n473), .B2(new_n719), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n733), .B1(new_n734), .B2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(G16), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G20), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(KEYINPUT96), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT23), .ZN(new_n743));
  INV_X1    g318(.A(G299), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(new_n740), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1956), .ZN(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT31), .B(G11), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT93), .Z(new_n748));
  NAND2_X1  g323(.A1(G164), .A2(G29), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G27), .B2(G29), .ZN(new_n750));
  INV_X1    g325(.A(G2078), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n751), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT30), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(G28), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(G28), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n755), .A2(new_n756), .A3(new_n719), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n624), .B2(new_n719), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n734), .B2(new_n738), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n752), .A2(new_n753), .A3(new_n759), .ZN(new_n760));
  NOR4_X1   g335(.A1(new_n739), .A2(new_n746), .A3(new_n748), .A4(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G29), .A2(G33), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n467), .A2(G103), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n465), .A2(G139), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n475), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n765), .B(new_n766), .C1(new_n466), .C2(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT90), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n762), .B1(new_n769), .B2(G29), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(G2072), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n740), .A2(G21), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G168), .B2(new_n740), .ZN(new_n773));
  INV_X1    g348(.A(G1966), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n761), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n740), .A2(G19), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n554), .B2(new_n740), .ZN(new_n780));
  MUX2_X1   g355(.A(new_n779), .B(new_n780), .S(KEYINPUT87), .Z(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(G1341), .Z(new_n782));
  NOR2_X1   g357(.A1(G29), .A2(G35), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G162), .B2(G29), .ZN(new_n784));
  INV_X1    g359(.A(G2090), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT94), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G5), .B2(G16), .ZN(new_n790));
  OR3_X1    g365(.A1(new_n789), .A2(G5), .A3(G16), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n790), .B(new_n791), .C1(G301), .C2(new_n740), .ZN(new_n792));
  INV_X1    g367(.A(G1961), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n788), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n740), .A2(G4), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n599), .B2(new_n740), .ZN(new_n797));
  INV_X1    g372(.A(G1348), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n778), .A2(new_n782), .A3(new_n795), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n740), .A2(G24), .ZN(new_n801));
  INV_X1    g376(.A(G290), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n802), .B2(new_n740), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1986), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n740), .A2(G22), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G166), .B2(new_n740), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1971), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n740), .A2(G23), .ZN(new_n808));
  INV_X1    g383(.A(G288), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(new_n740), .ZN(new_n810));
  XOR2_X1   g385(.A(new_n810), .B(KEYINPUT33), .Z(new_n811));
  AOI21_X1  g386(.A(new_n807), .B1(new_n811), .B2(G1976), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n740), .A2(G6), .ZN(new_n813));
  INV_X1    g388(.A(G305), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(new_n740), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT32), .B(G1981), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  OAI211_X1 g392(.A(new_n812), .B(new_n817), .C1(G1976), .C2(new_n811), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n804), .B1(new_n818), .B2(KEYINPUT34), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n465), .A2(G131), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT85), .ZN(new_n821));
  OR2_X1    g396(.A1(G95), .A2(G2105), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n822), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n714), .A2(G119), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n821), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  MUX2_X1   g400(.A(G25), .B(new_n825), .S(G29), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT86), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT35), .B(G1991), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n819), .B(new_n829), .C1(KEYINPUT34), .C2(new_n818), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(KEYINPUT36), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(KEYINPUT36), .ZN(new_n832));
  AOI211_X1 g407(.A(new_n722), .B(new_n800), .C1(new_n831), .C2(new_n832), .ZN(G311));
  AOI21_X1  g408(.A(new_n800), .B1(new_n831), .B2(new_n832), .ZN(new_n834));
  INV_X1    g409(.A(new_n722), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(G150));
  INV_X1    g411(.A(G67), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(new_n537), .B2(new_n538), .ZN(new_n838));
  AND2_X1   g413(.A1(G80), .A2(G543), .ZN(new_n839));
  OAI21_X1  g414(.A(G651), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n529), .A2(G55), .A3(new_n531), .ZN(new_n841));
  XOR2_X1   g416(.A(KEYINPUT97), .B(G93), .Z(new_n842));
  NAND2_X1  g417(.A1(new_n507), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n840), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n840), .A2(new_n841), .A3(KEYINPUT98), .A4(new_n843), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(new_n553), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n548), .B(new_n844), .C1(new_n551), .C2(new_n552), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT38), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n598), .A2(new_n606), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT39), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(G860), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n853), .A2(new_n855), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT99), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n848), .A2(new_n857), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT37), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(KEYINPUT100), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n861), .A2(new_n866), .A3(new_n863), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(G145));
  INV_X1    g443(.A(KEYINPUT40), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n624), .B(new_n473), .ZN(new_n870));
  XNOR2_X1  g445(.A(G162), .B(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n718), .B(new_n729), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n872), .A2(new_n496), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n718), .B(new_n728), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(G164), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n873), .A2(new_n875), .A3(new_n768), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n873), .A2(new_n875), .ZN(new_n877));
  INV_X1    g452(.A(new_n769), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n825), .A2(new_n617), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n714), .A2(G130), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n465), .A2(G142), .ZN(new_n882));
  OR2_X1    g457(.A1(G106), .A2(G2105), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n883), .B(G2104), .C1(G118), .C2(new_n466), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n881), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n825), .A2(new_n617), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n880), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n825), .A2(new_n617), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n885), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n879), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT102), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT101), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n889), .A2(new_n890), .A3(new_n885), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n886), .B1(new_n880), .B2(new_n887), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n891), .A2(KEYINPUT101), .A3(new_n888), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n878), .B1(new_n873), .B2(new_n875), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n901), .B1(new_n768), .B2(new_n877), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n893), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NOR3_X1   g478(.A1(new_n879), .A2(new_n899), .A3(KEYINPUT102), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n871), .B(new_n892), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n900), .A2(new_n902), .A3(new_n893), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT102), .B1(new_n879), .B2(new_n899), .ZN(new_n908));
  AOI22_X1  g483(.A1(new_n907), .A2(new_n908), .B1(new_n899), .B2(new_n879), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n905), .B(new_n906), .C1(new_n871), .C2(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n910), .A2(KEYINPUT103), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT103), .ZN(new_n912));
  OAI22_X1  g487(.A1(new_n903), .A2(new_n904), .B1(new_n900), .B2(new_n902), .ZN(new_n913));
  INV_X1    g488(.A(new_n871), .ZN(new_n914));
  AOI21_X1  g489(.A(G37), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n912), .B1(new_n915), .B2(new_n905), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n869), .B1(new_n911), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n910), .A2(KEYINPUT103), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(new_n912), .A3(new_n905), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n919), .A3(KEYINPUT40), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(G395));
  INV_X1    g496(.A(new_n851), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n610), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n851), .A2(new_n609), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n598), .A2(new_n744), .ZN(new_n926));
  AOI21_X1  g501(.A(G299), .B1(new_n596), .B2(new_n597), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT104), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n599), .A2(G299), .ZN(new_n932));
  INV_X1    g507(.A(new_n927), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n932), .A2(KEYINPUT41), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT41), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n935), .B1(new_n926), .B2(new_n927), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n923), .A2(new_n924), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n925), .A2(new_n939), .A3(new_n929), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n931), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT42), .ZN(new_n942));
  NAND2_X1  g517(.A1(G166), .A2(G288), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n809), .A2(G303), .ZN(new_n944));
  AOI21_X1  g519(.A(G290), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(G290), .A2(new_n944), .A3(new_n943), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(new_n814), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n947), .ZN(new_n949));
  OAI21_X1  g524(.A(G305), .B1(new_n949), .B2(new_n945), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT42), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n931), .A2(new_n952), .A3(new_n938), .A4(new_n940), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n942), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n951), .B1(new_n942), .B2(new_n953), .ZN(new_n955));
  OAI21_X1  g530(.A(G868), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n956), .B1(G868), .B2(new_n848), .ZN(G295));
  OAI21_X1  g532(.A(new_n956), .B1(G868), .B2(new_n848), .ZN(G331));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n959), .B1(G168), .B2(G301), .ZN(new_n960));
  NAND3_X1  g535(.A1(G171), .A2(KEYINPUT106), .A3(G286), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n963), .B1(G171), .B2(G286), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n526), .A2(new_n532), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n965), .A2(KEYINPUT105), .A3(new_n528), .A4(G301), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n962), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n851), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n962), .A2(new_n967), .A3(new_n849), .A4(new_n850), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n969), .A2(KEYINPUT107), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n968), .A2(new_n851), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(new_n937), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n969), .A2(new_n929), .A3(new_n970), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(new_n951), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(new_n906), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n951), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n948), .A2(new_n950), .A3(KEYINPUT108), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n974), .A2(new_n975), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT43), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT109), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n979), .A2(new_n980), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n936), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n937), .A2(KEYINPUT110), .ZN(new_n987));
  AOI211_X1 g562(.A(new_n986), .B(new_n987), .C1(new_n969), .C2(new_n970), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n928), .B1(new_n971), .B2(new_n973), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n984), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n990), .A2(new_n991), .A3(new_n906), .A4(new_n976), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n993), .B(KEYINPUT43), .C1(new_n977), .C2(new_n981), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n983), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT44), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n991), .B1(new_n977), .B2(new_n981), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n990), .A2(new_n906), .A3(new_n976), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n998), .B1(new_n999), .B2(new_n991), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(KEYINPUT44), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n997), .A2(new_n1001), .ZN(G397));
  NAND3_X1  g577(.A1(new_n468), .A2(new_n472), .A3(G40), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n1003), .B(KEYINPUT111), .ZN(new_n1004));
  INV_X1    g579(.A(G1384), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT45), .B1(new_n496), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  OR2_X1    g582(.A1(new_n1007), .A2(G1996), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(new_n718), .ZN(new_n1009));
  XOR2_X1   g584(.A(new_n1009), .B(KEYINPUT112), .Z(new_n1010));
  XOR2_X1   g585(.A(new_n1007), .B(KEYINPUT113), .Z(new_n1011));
  NAND3_X1  g586(.A1(new_n1011), .A2(G1996), .A3(new_n718), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n728), .B(G2067), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1010), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  XOR2_X1   g590(.A(new_n825), .B(new_n828), .Z(new_n1016));
  INV_X1    g591(.A(KEYINPUT114), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1016), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1011), .B1(KEYINPUT114), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1015), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1007), .ZN(new_n1022));
  XNOR2_X1  g597(.A(G290), .B(G1986), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1025));
  OR2_X1    g600(.A1(new_n1025), .A2(KEYINPUT116), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n1027));
  INV_X1    g602(.A(G8), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1027), .B1(G166), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1025), .A2(KEYINPUT116), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1026), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(G1384), .B1(new_n490), .B2(new_n495), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1032), .A2(KEYINPUT50), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n1034));
  AOI211_X1 g609(.A(new_n1034), .B(G1384), .C1(new_n490), .C2(new_n495), .ZN(new_n1035));
  OR2_X1    g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1036), .A2(new_n785), .A3(new_n1004), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT115), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n496), .A2(new_n1005), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT45), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1032), .A2(KEYINPUT45), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(new_n1004), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1971), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1037), .B1(new_n1038), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT115), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1047));
  OAI211_X1 g622(.A(G8), .B(new_n1031), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1028), .B1(new_n1037), .B2(new_n1045), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT119), .B1(new_n1049), .B2(new_n1031), .ZN(new_n1050));
  XNOR2_X1  g625(.A(G305), .B(KEYINPUT49), .ZN(new_n1051));
  INV_X1    g626(.A(G1981), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1052), .B1(new_n579), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1028), .B1(new_n1004), .B2(new_n1032), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1976), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1057), .B1(new_n1060), .B2(G288), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT52), .ZN(new_n1062));
  AOI21_X1  g637(.A(KEYINPUT52), .B1(G288), .B2(new_n1060), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1057), .B(new_n1063), .C1(new_n1060), .C2(G288), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1059), .A2(new_n1062), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1048), .A2(new_n1050), .A3(new_n1065), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1049), .A2(KEYINPUT119), .A3(new_n1031), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  XNOR2_X1  g643(.A(KEYINPUT121), .B(G2084), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1036), .A2(new_n1004), .A3(new_n1069), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1043), .A2(KEYINPUT120), .A3(new_n774), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT120), .B1(new_n1043), .B2(new_n774), .ZN(new_n1072));
  OAI211_X1 g647(.A(G168), .B(new_n1070), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT124), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(G8), .A3(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1078), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1073), .A2(G8), .A3(new_n1076), .A4(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(G8), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1079), .B(new_n1081), .C1(G168), .C2(new_n1083), .ZN(new_n1084));
  AOI211_X1 g659(.A(new_n1040), .B(G1384), .C1(new_n490), .C2(new_n495), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1006), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1086), .A2(new_n751), .A3(new_n1004), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT125), .B(KEYINPUT53), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1004), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n793), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1089), .B(new_n1091), .C1(new_n1092), .C2(new_n1087), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(G171), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT62), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1068), .B1(new_n1084), .B2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT56), .B(G2072), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1041), .A2(new_n1004), .A3(new_n1042), .A4(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT123), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT123), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1086), .A2(new_n1101), .A3(new_n1004), .A4(new_n1098), .ZN(new_n1102));
  INV_X1    g677(.A(G1956), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1090), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1100), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT57), .ZN(new_n1107));
  OAI21_X1  g682(.A(G299), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1108), .B(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1105), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1110), .A2(new_n1100), .A3(new_n1102), .A4(new_n1104), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT61), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1090), .A2(new_n798), .ZN(new_n1117));
  INV_X1    g692(.A(G2067), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1004), .A2(new_n1118), .A3(new_n1032), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1117), .A2(new_n598), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n598), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1121));
  OAI21_X1  g696(.A(KEYINPUT60), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n598), .A2(KEYINPUT60), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1117), .A2(new_n1119), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1004), .A2(new_n1032), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT58), .B(G1341), .Z(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1127), .B1(new_n1043), .B2(G1996), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n554), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT59), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1128), .A2(new_n1131), .A3(new_n554), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1124), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1112), .A2(KEYINPUT61), .A3(new_n1113), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1116), .A2(new_n1122), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1113), .A2(new_n1121), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1135), .A2(new_n1136), .A3(new_n1112), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1003), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1092), .A2(G2078), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1041), .A2(new_n1042), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(KEYINPUT126), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1141), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1142));
  OAI21_X1  g717(.A(KEYINPUT127), .B1(new_n1142), .B2(G171), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT54), .ZN(new_n1144));
  AND2_X1   g719(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT127), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1145), .A2(new_n1146), .A3(G301), .A4(new_n1141), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1143), .A2(new_n1094), .A3(new_n1144), .A4(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1144), .B1(new_n1093), .B2(G301), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(G301), .B2(new_n1142), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1137), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1093), .A2(new_n1095), .A3(G171), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n1084), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1097), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1048), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n1065), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1059), .A2(new_n1060), .A3(new_n809), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1158), .B1(G1981), .B2(G305), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1057), .B(KEYINPUT118), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1083), .A2(G286), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT63), .B1(new_n1068), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT63), .ZN(new_n1164));
  OAI21_X1  g739(.A(G8), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1031), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AND4_X1   g742(.A1(new_n1048), .A2(new_n1167), .A3(new_n1065), .A4(new_n1162), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1157), .B(new_n1161), .C1(new_n1163), .C2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1024), .B1(new_n1155), .B2(new_n1169), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1007), .A2(G290), .A3(G1986), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT48), .ZN(new_n1172));
  NOR2_X1   g747(.A1(new_n1021), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1011), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n825), .A2(new_n828), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1015), .A2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n729), .A2(new_n1118), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1174), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1011), .B1(new_n718), .B2(new_n1013), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1008), .B(KEYINPUT46), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1181), .B(KEYINPUT47), .Z(new_n1182));
  NOR3_X1   g757(.A1(new_n1173), .A2(new_n1178), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1170), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g759(.A1(new_n910), .A2(new_n663), .A3(new_n690), .ZN(new_n1186));
  NOR2_X1   g760(.A1(G229), .A2(new_n461), .ZN(new_n1187));
  AND3_X1   g761(.A1(new_n1186), .A2(new_n995), .A3(new_n1187), .ZN(G308));
  NAND3_X1  g762(.A1(new_n1186), .A2(new_n995), .A3(new_n1187), .ZN(G225));
endmodule


