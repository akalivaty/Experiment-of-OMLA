//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:57 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1283, new_n1284, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1351, new_n1352, new_n1353;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n213), .B(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n216));
  INV_X1    g0016(.A(G77), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  INV_X1    g0018(.A(G264), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n205), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n211), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n209), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n202), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n215), .B(new_n225), .C1(new_n227), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT65), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G68), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n226), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n209), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(G150), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  OAI22_X1  g0054(.A1(new_n250), .A2(new_n251), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G50), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n209), .B1(new_n201), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n249), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(new_n226), .A3(new_n248), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n256), .B1(new_n208), .B2(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n259), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n261), .A2(new_n262), .B1(new_n256), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n258), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(new_n265), .B(KEYINPUT9), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G223), .A3(G1698), .ZN(new_n272));
  INV_X1    g0072(.A(G1698), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n271), .A2(G222), .A3(new_n273), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n272), .B(new_n274), .C1(new_n217), .C2(new_n271), .ZN(new_n275));
  AND2_X1   g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(new_n226), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(KEYINPUT66), .B1(new_n276), .B2(new_n226), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT66), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n280), .A2(new_n281), .A3(G1), .A4(G13), .ZN(new_n282));
  INV_X1    g0082(.A(G41), .ZN(new_n283));
  INV_X1    g0083(.A(G45), .ZN(new_n284));
  AOI21_X1  g0084(.A(G1), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n279), .A2(G274), .A3(new_n282), .A4(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n279), .A2(new_n282), .ZN(new_n287));
  INV_X1    g0087(.A(new_n285), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(G226), .A3(new_n288), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n278), .A2(G190), .A3(new_n286), .A4(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n278), .A2(new_n286), .A3(new_n289), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G200), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n266), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT10), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT10), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n266), .A2(new_n295), .A3(new_n290), .A4(new_n292), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  XOR2_X1   g0097(.A(KEYINPUT67), .B(G179), .Z(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n291), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n291), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n300), .A2(new_n265), .A3(new_n302), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n288), .A2(new_n279), .A3(G244), .A4(new_n282), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(new_n286), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT68), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT68), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n304), .A2(new_n286), .A3(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(G232), .A2(G1698), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n273), .A2(G238), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n271), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n311), .B(new_n277), .C1(G107), .C2(new_n271), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n306), .A2(new_n308), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G200), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT69), .ZN(new_n315));
  OAI21_X1  g0115(.A(G77), .B1(new_n209), .B2(G1), .ZN(new_n316));
  OR3_X1    g0116(.A1(new_n260), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n315), .B1(new_n260), .B2(new_n316), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n263), .A2(new_n217), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n250), .A2(new_n254), .B1(new_n209), .B2(new_n217), .ZN(new_n321));
  XNOR2_X1  g0121(.A(KEYINPUT15), .B(G87), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(new_n251), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n249), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n319), .A2(new_n320), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n313), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(G190), .ZN(new_n327));
  INV_X1    g0127(.A(new_n325), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n328), .B1(new_n301), .B2(new_n313), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n326), .A2(new_n298), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n314), .A2(new_n327), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n297), .A2(new_n303), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G58), .ZN(new_n333));
  INV_X1    g0133(.A(G68), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(G20), .B1(new_n335), .B2(new_n201), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n253), .A2(G159), .ZN(new_n337));
  AND2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n268), .A2(KEYINPUT74), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT74), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G33), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(new_n341), .A3(new_n267), .ZN(new_n342));
  AND2_X1   g0142(.A1(KEYINPUT3), .A2(G33), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT7), .ZN(new_n344));
  NOR3_X1   g0144(.A1(new_n343), .A2(new_n344), .A3(G20), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n269), .A2(new_n209), .A3(new_n270), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n342), .A2(new_n345), .B1(new_n346), .B2(new_n344), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n338), .B1(new_n347), .B2(new_n334), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT16), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT74), .B(G33), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n209), .B(new_n269), .C1(new_n351), .C2(new_n267), .ZN(new_n352));
  OAI21_X1  g0152(.A(G68), .B1(new_n352), .B2(KEYINPUT7), .ZN(new_n353));
  NOR2_X1   g0153(.A1(KEYINPUT3), .A2(G33), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n339), .A2(new_n341), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n354), .B1(new_n355), .B2(KEYINPUT3), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n344), .B1(new_n356), .B2(new_n209), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n338), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n350), .B(new_n249), .C1(new_n358), .C2(new_n349), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n250), .B1(new_n208), .B2(G20), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(new_n261), .B1(new_n263), .B2(new_n250), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n269), .B1(new_n351), .B2(new_n267), .ZN(new_n363));
  NOR2_X1   g0163(.A1(G223), .A2(G1698), .ZN(new_n364));
  INV_X1    g0164(.A(G226), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(G1698), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n363), .A2(new_n366), .B1(G33), .B2(G87), .ZN(new_n367));
  INV_X1    g0167(.A(new_n277), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n287), .A2(G232), .A3(new_n288), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n286), .ZN(new_n371));
  OAI21_X1  g0171(.A(G169), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n369), .A2(new_n371), .A3(new_n298), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT75), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n369), .A2(new_n371), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(new_n299), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT75), .B1(new_n378), .B2(new_n372), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n362), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT18), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n377), .A2(G190), .ZN(new_n382));
  OAI21_X1  g0182(.A(G200), .B1(new_n369), .B2(new_n371), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n382), .A2(new_n359), .A3(new_n361), .A4(new_n383), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n384), .B(KEYINPUT17), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n375), .B1(new_n373), .B2(new_n374), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n378), .A2(KEYINPUT75), .A3(new_n372), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT18), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n388), .A2(new_n389), .A3(new_n362), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n332), .A2(new_n381), .A3(new_n385), .A4(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n365), .A2(new_n273), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n232), .A2(G1698), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n392), .B(new_n393), .C1(new_n343), .C2(new_n354), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT70), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G97), .ZN(new_n396));
  AND3_X1   g0196(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n395), .B1(new_n394), .B2(new_n396), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n397), .A2(new_n398), .A3(new_n368), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n288), .A2(new_n279), .A3(G238), .A4(new_n282), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n286), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT13), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT13), .ZN(new_n403));
  INV_X1    g0203(.A(new_n401), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n394), .A2(new_n396), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n277), .B1(new_n405), .B2(new_n395), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n403), .B(new_n404), .C1(new_n406), .C2(new_n397), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT71), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n402), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  OAI211_X1 g0209(.A(KEYINPUT71), .B(KEYINPUT13), .C1(new_n399), .C2(new_n401), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(G169), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT14), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT14), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n409), .A2(new_n413), .A3(G169), .A4(new_n410), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n402), .A2(new_n407), .A3(G179), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n412), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n251), .A2(new_n217), .B1(new_n209), .B2(G68), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT72), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n417), .A2(new_n418), .B1(new_n256), .B2(new_n254), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n417), .A2(new_n418), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n249), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT11), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI211_X1 g0223(.A(KEYINPUT11), .B(new_n249), .C1(new_n419), .C2(new_n420), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT73), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n423), .A2(KEYINPUT73), .A3(new_n424), .ZN(new_n428));
  OAI21_X1  g0228(.A(KEYINPUT12), .B1(new_n259), .B2(G68), .ZN(new_n429));
  OR3_X1    g0229(.A1(new_n259), .A2(KEYINPUT12), .A3(G68), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n334), .B1(new_n208), .B2(G20), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n429), .A2(new_n430), .B1(new_n261), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n427), .A2(new_n428), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n416), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n433), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n409), .A2(G200), .A3(new_n410), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n402), .A2(new_n407), .A3(G190), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n391), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n218), .A2(G1698), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n271), .A2(KEYINPUT4), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n271), .A2(G250), .A3(G1698), .ZN(new_n444));
  NAND2_X1  g0244(.A1(G33), .A2(G283), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT77), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n267), .B1(new_n339), .B2(new_n341), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n447), .B(new_n442), .C1(new_n448), .C2(new_n354), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT4), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n447), .B1(new_n363), .B2(new_n442), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n446), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n277), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n279), .A2(G274), .A3(new_n282), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT79), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT5), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n456), .B1(new_n457), .B2(G41), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n283), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n284), .A2(G1), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n457), .A2(G41), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n458), .A2(new_n459), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  OR2_X1    g0262(.A1(new_n455), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(G257), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n287), .A2(new_n462), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(G169), .B1(new_n454), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n263), .A2(new_n204), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n260), .B1(new_n208), .B2(G33), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n469), .B1(new_n471), .B2(new_n204), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n253), .A2(G77), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G97), .A2(G107), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT6), .B1(new_n206), .B2(new_n474), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n205), .A2(KEYINPUT6), .A3(G97), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n473), .B1(new_n477), .B2(new_n209), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n345), .A2(new_n342), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n346), .A2(new_n344), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n205), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n249), .B1(new_n478), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(KEYINPUT76), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT76), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n484), .B(new_n249), .C1(new_n478), .C2(new_n481), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n472), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n468), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT78), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n453), .A2(new_n488), .A3(new_n277), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n488), .B1(new_n453), .B2(new_n277), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n298), .B(new_n467), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(new_n322), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(new_n259), .ZN(new_n495));
  XNOR2_X1  g0295(.A(KEYINPUT82), .B(KEYINPUT19), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n396), .A2(new_n209), .ZN(new_n497));
  INV_X1    g0297(.A(G87), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(new_n204), .A3(new_n205), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n496), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n251), .A2(new_n204), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(new_n496), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n363), .A2(new_n209), .A3(G68), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n495), .B1(new_n505), .B2(new_n249), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(new_n322), .B2(new_n471), .ZN(new_n507));
  AND4_X1   g0307(.A1(G274), .A2(new_n279), .A3(new_n282), .A4(new_n460), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n355), .A2(G116), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n218), .A2(G1698), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(G238), .B2(G1698), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n509), .B1(new_n356), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n508), .B1(new_n512), .B2(new_n277), .ZN(new_n513));
  INV_X1    g0313(.A(G250), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n460), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(new_n279), .A3(new_n282), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT81), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n515), .A2(new_n279), .A3(KEYINPUT81), .A4(new_n282), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n513), .A2(new_n299), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n301), .B1(new_n513), .B2(new_n520), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n507), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n340), .A2(G33), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n268), .A2(KEYINPUT74), .ZN(new_n525));
  OAI21_X1  g0325(.A(KEYINPUT3), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n511), .B1(new_n526), .B2(new_n269), .ZN(new_n527));
  INV_X1    g0327(.A(new_n509), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n277), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(new_n508), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n529), .A2(new_n520), .A3(G190), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT83), .ZN(new_n532));
  INV_X1    g0332(.A(new_n249), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n533), .B1(new_n503), .B2(new_n504), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n471), .A2(new_n498), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n534), .A2(new_n535), .A3(new_n495), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n529), .A2(new_n520), .A3(new_n530), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G200), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT83), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n513), .A2(new_n539), .A3(G190), .A4(new_n520), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n532), .A2(new_n536), .A3(new_n538), .A4(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n523), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n454), .A2(new_n467), .ZN(new_n543));
  INV_X1    g0343(.A(G190), .ZN(new_n544));
  OAI21_X1  g0344(.A(KEYINPUT80), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n466), .B1(new_n453), .B2(new_n277), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT80), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n546), .A2(new_n547), .A3(G190), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n545), .A2(new_n486), .A3(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(G200), .ZN(new_n550));
  INV_X1    g0350(.A(new_n491), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n489), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n550), .B1(new_n552), .B2(new_n467), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n493), .B(new_n542), .C1(new_n549), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n205), .A2(G20), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(G13), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n557), .A2(G1), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n556), .B(new_n558), .C1(KEYINPUT86), .C2(KEYINPUT25), .ZN(new_n559));
  NAND2_X1  g0359(.A1(KEYINPUT86), .A2(KEYINPUT25), .ZN(new_n560));
  OR2_X1    g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n560), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n561), .A2(new_n562), .B1(new_n470), .B2(G107), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT22), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n564), .A2(new_n498), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n209), .B(new_n565), .C1(new_n448), .C2(new_n354), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT23), .ZN(new_n568));
  AOI22_X1  g0368(.A1(KEYINPUT84), .A2(new_n568), .B1(new_n205), .B2(G20), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(KEYINPUT84), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT84), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT23), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n569), .B1(new_n556), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n343), .A2(new_n354), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n209), .A2(G87), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n564), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n355), .A2(new_n209), .A3(G116), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n574), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(KEYINPUT24), .B1(new_n567), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(G116), .ZN(new_n581));
  NOR3_X1   g0381(.A1(new_n351), .A2(G20), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n570), .A2(new_n555), .ZN(new_n583));
  XNOR2_X1  g0383(.A(KEYINPUT84), .B(KEYINPUT23), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n583), .B1(new_n584), .B2(new_n555), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT24), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n586), .A2(new_n587), .A3(new_n566), .A4(new_n577), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n580), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT85), .B1(new_n589), .B2(new_n249), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT85), .ZN(new_n591));
  AOI211_X1 g0391(.A(new_n591), .B(new_n533), .C1(new_n580), .C2(new_n588), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n563), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(G250), .A2(G1698), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n464), .B2(G1698), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n363), .A2(new_n595), .B1(G294), .B2(new_n355), .ZN(new_n596));
  OAI221_X1 g0396(.A(new_n463), .B1(new_n465), .B2(new_n219), .C1(new_n368), .C2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n301), .ZN(new_n598));
  INV_X1    g0398(.A(new_n465), .ZN(new_n599));
  INV_X1    g0399(.A(new_n595), .ZN(new_n600));
  INV_X1    g0400(.A(G294), .ZN(new_n601));
  OAI22_X1  g0401(.A1(new_n356), .A2(new_n600), .B1(new_n601), .B2(new_n351), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n599), .A2(G264), .B1(new_n602), .B2(new_n277), .ZN(new_n603));
  INV_X1    g0403(.A(G179), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n604), .A3(new_n463), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n598), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n593), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n597), .A2(new_n550), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(G190), .B2(new_n597), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n610), .B(new_n563), .C1(new_n590), .C2(new_n592), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n462), .A2(G270), .A3(new_n279), .A4(new_n282), .ZN(new_n613));
  NOR2_X1   g0413(.A1(G257), .A2(G1698), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n614), .B1(new_n219), .B2(G1698), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n448), .B2(new_n354), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n575), .A2(G303), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n463), .B(new_n613), .C1(new_n618), .C2(new_n368), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n445), .B(new_n209), .C1(G33), .C2(new_n204), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n581), .A2(G20), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(new_n249), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT20), .ZN(new_n623));
  XNOR2_X1  g0423(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n259), .A2(G116), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(new_n470), .B2(G116), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n301), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n619), .A2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT21), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n619), .A2(new_n627), .A3(KEYINPUT21), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n613), .B1(new_n455), .B2(new_n462), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n368), .B1(new_n616), .B2(new_n617), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n632), .A2(new_n633), .A3(new_n604), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n624), .A2(new_n626), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n630), .A2(new_n631), .A3(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n632), .A2(new_n633), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(G190), .ZN(new_n639));
  INV_X1    g0439(.A(new_n635), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n639), .B(new_n640), .C1(new_n550), .C2(new_n638), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NOR4_X1   g0442(.A1(new_n441), .A2(new_n554), .A3(new_n612), .A4(new_n642), .ZN(G372));
  INV_X1    g0443(.A(new_n303), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n378), .A2(new_n372), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n362), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n646), .B(new_n389), .ZN(new_n647));
  INV_X1    g0447(.A(new_n415), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n648), .B1(new_n411), .B2(KEYINPUT14), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n435), .B1(new_n649), .B2(new_n414), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n329), .A2(new_n330), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n650), .B1(new_n438), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n385), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n647), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n644), .B1(new_n655), .B2(new_n297), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT87), .B1(new_n521), .B2(new_n522), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n537), .A2(G169), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT87), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n513), .A2(new_n299), .A3(new_n520), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n662), .A2(KEYINPUT89), .A3(new_n507), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT89), .B1(new_n662), .B2(new_n507), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n563), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n589), .A2(new_n249), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n591), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n589), .A2(KEYINPUT85), .A3(new_n249), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n666), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n637), .B1(new_n670), .B2(new_n606), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT88), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n537), .A2(new_n672), .A3(G200), .ZN(new_n673));
  INV_X1    g0473(.A(new_n535), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n506), .A2(new_n531), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n672), .B1(new_n537), .B2(G200), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI22_X1  g0477(.A1(new_n662), .A2(new_n507), .B1(new_n673), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n671), .A2(new_n611), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n493), .B1(new_n549), .B2(new_n553), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n665), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT26), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n523), .A2(new_n541), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n493), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n487), .A2(new_n492), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n678), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n684), .B1(new_n682), .B2(new_n686), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n656), .B1(new_n689), .B2(new_n441), .ZN(G369));
  NAND3_X1  g0490(.A1(new_n630), .A2(new_n631), .A3(new_n636), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n558), .A2(new_n209), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(KEYINPUT27), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n693), .A2(G213), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(G343), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n640), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n691), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n642), .B2(new_n699), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n701), .A2(G330), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n670), .A2(new_n698), .ZN(new_n703));
  OAI22_X1  g0503(.A1(new_n612), .A2(new_n703), .B1(new_n608), .B2(new_n698), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n691), .A2(new_n698), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n708), .A2(new_n608), .A3(new_n611), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n608), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n710), .B1(new_n711), .B2(new_n698), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n706), .A2(new_n712), .ZN(G399));
  INV_X1    g0513(.A(new_n212), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G41), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n499), .A2(G116), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(G1), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n228), .B2(new_n716), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  INV_X1    g0520(.A(G330), .ZN(new_n721));
  OAI22_X1  g0521(.A1(new_n596), .A2(new_n368), .B1(new_n465), .B2(new_n219), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n537), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n546), .A2(new_n723), .A3(new_n634), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT90), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n725), .B1(new_n724), .B2(new_n726), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n467), .B1(new_n490), .B2(new_n491), .ZN(new_n730));
  AND4_X1   g0530(.A1(new_n298), .A2(new_n597), .A3(new_n619), .A4(new_n537), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n634), .A2(new_n520), .A3(new_n603), .A4(new_n513), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n543), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n730), .A2(new_n731), .B1(new_n733), .B2(KEYINPUT30), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n698), .B1(new_n729), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(KEYINPUT91), .B1(new_n735), .B2(KEYINPUT31), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n726), .B1(new_n732), .B2(new_n543), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(KEYINPUT90), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n730), .A2(new_n731), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n733), .A2(KEYINPUT30), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n738), .A2(new_n739), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n697), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT91), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n736), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n697), .A2(KEYINPUT31), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n748), .B1(new_n734), .B2(new_n737), .ZN(new_n749));
  INV_X1    g0549(.A(new_n554), .ZN(new_n750));
  AND4_X1   g0550(.A1(new_n630), .A2(new_n641), .A3(new_n631), .A4(new_n636), .ZN(new_n751));
  AND4_X1   g0551(.A1(new_n608), .A2(new_n751), .A3(new_n611), .A4(new_n698), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n749), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n721), .B1(new_n747), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT29), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n755), .B(new_n698), .C1(new_n681), .C2(new_n687), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n608), .A2(new_n637), .B1(new_n670), .B2(new_n610), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n730), .A2(G200), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n759), .A2(new_n486), .A3(new_n548), .A4(new_n545), .ZN(new_n760));
  NAND4_X1  g0560(.A1(new_n758), .A2(new_n493), .A3(new_n760), .A4(new_n678), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n686), .A2(KEYINPUT26), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n685), .A2(new_n682), .A3(new_n542), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n761), .A2(new_n665), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n755), .B1(new_n764), .B2(new_n698), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n754), .A2(new_n757), .A3(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n720), .B1(new_n766), .B2(G1), .ZN(G364));
  NOR2_X1   g0567(.A1(new_n557), .A2(G20), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n208), .B1(new_n768), .B2(G45), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n715), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n702), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(G330), .B2(new_n701), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n212), .A2(new_n271), .ZN(new_n774));
  INV_X1    g0574(.A(G355), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n774), .A2(new_n775), .B1(G116), .B2(new_n212), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n714), .A2(new_n363), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(new_n284), .B2(new_n229), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n246), .A2(G45), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI211_X1 g0581(.A(G1), .B(G13), .C1(new_n209), .C2(G169), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT93), .Z(new_n783));
  NOR2_X1   g0583(.A1(G13), .A2(G33), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n209), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT92), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT94), .Z(new_n788));
  OAI21_X1  g0588(.A(new_n771), .B1(new_n781), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n209), .A2(G179), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G190), .A2(G200), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n271), .B1(new_n793), .B2(G329), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n544), .A2(G179), .A3(G200), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n209), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n794), .B1(new_n601), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n298), .A2(new_n209), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n791), .ZN(new_n799));
  INV_X1    g0599(.A(G311), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n544), .A2(G200), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n798), .A2(new_n802), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n797), .B(new_n801), .C1(G322), .C2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(G326), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n798), .A2(G190), .A3(G200), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n798), .A2(new_n544), .A3(G200), .ZN(new_n807));
  XOR2_X1   g0607(.A(KEYINPUT33), .B(G317), .Z(new_n808));
  OAI22_X1  g0608(.A1(new_n805), .A2(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n790), .A2(G190), .A3(G200), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n810), .A2(KEYINPUT96), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(KEYINPUT96), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n809), .B1(G303), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n790), .A2(new_n544), .A3(G200), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT97), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT98), .Z(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(G283), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n804), .B(new_n815), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n818), .A2(G107), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n814), .A2(G87), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n822), .A2(new_n271), .A3(new_n823), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT99), .Z(new_n825));
  INV_X1    g0625(.A(new_n796), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(G97), .ZN(new_n827));
  INV_X1    g0627(.A(new_n803), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n827), .B1(new_n828), .B2(new_n333), .ZN(new_n829));
  INV_X1    g0629(.A(G159), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n792), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(KEYINPUT95), .B(KEYINPUT32), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n831), .B(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n217), .B2(new_n799), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n256), .A2(new_n806), .B1(new_n807), .B2(new_n334), .ZN(new_n835));
  OR3_X1    g0635(.A1(new_n829), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n821), .B1(new_n825), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n783), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n789), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n701), .B2(new_n786), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n773), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G396));
  NAND2_X1  g0642(.A1(new_n652), .A2(new_n698), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n327), .A2(new_n314), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n325), .A2(new_n697), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n651), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n689), .A2(new_n697), .B1(new_n844), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n844), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n698), .B(new_n851), .C1(new_n681), .C2(new_n687), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n754), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n853), .A2(new_n771), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n850), .A2(new_n754), .A3(new_n852), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n271), .B1(new_n793), .B2(G311), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n827), .B(new_n857), .C1(new_n828), .C2(new_n601), .ZN(new_n858));
  INV_X1    g0658(.A(new_n799), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n858), .B1(G116), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n818), .A2(G87), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n814), .A2(G107), .ZN(new_n862));
  INV_X1    g0662(.A(new_n807), .ZN(new_n863));
  INV_X1    g0663(.A(new_n806), .ZN(new_n864));
  AOI22_X1  g0664(.A1(G283), .A2(new_n863), .B1(new_n864), .B2(G303), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n860), .A2(new_n861), .A3(new_n862), .A4(new_n865), .ZN(new_n866));
  AOI22_X1  g0666(.A1(G159), .A2(new_n859), .B1(new_n803), .B2(G143), .ZN(new_n867));
  INV_X1    g0667(.A(G137), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n867), .B1(new_n868), .B2(new_n806), .C1(new_n252), .C2(new_n807), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT34), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n818), .A2(G68), .ZN(new_n872));
  INV_X1    g0672(.A(G132), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n363), .B1(new_n873), .B2(new_n792), .C1(new_n333), .C2(new_n796), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n814), .B2(G50), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n871), .A2(new_n872), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n869), .A2(new_n870), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n866), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n838), .ZN(new_n879));
  INV_X1    g0679(.A(new_n771), .ZN(new_n880));
  INV_X1    g0680(.A(new_n784), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n783), .A2(new_n881), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n882), .B(KEYINPUT100), .Z(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n880), .B1(new_n884), .B2(new_n217), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n879), .B(new_n885), .C1(new_n851), .C2(new_n881), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n856), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(G384));
  NOR2_X1   g0688(.A1(new_n768), .A2(new_n208), .ZN(new_n889));
  INV_X1    g0689(.A(new_n695), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n647), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n362), .A2(new_n890), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n647), .B2(new_n385), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n893), .A2(new_n384), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n646), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT37), .B1(new_n388), .B2(new_n362), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n896), .A2(KEYINPUT37), .B1(new_n897), .B2(new_n895), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n892), .B1(new_n894), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n381), .A2(new_n385), .A3(new_n390), .ZN(new_n900));
  AND2_X1   g0700(.A1(new_n358), .A2(new_n349), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n249), .B1(new_n358), .B2(new_n349), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n361), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n890), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n897), .A2(new_n895), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n903), .A2(new_n645), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(new_n904), .A3(new_n384), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT37), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n906), .A2(KEYINPUT38), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT39), .B1(new_n899), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n906), .A2(new_n911), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n892), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n915), .A2(new_n912), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n913), .B1(new_n916), .B2(KEYINPUT39), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n434), .A2(new_n697), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n891), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n852), .A2(new_n843), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(KEYINPUT103), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT103), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n852), .A2(new_n922), .A3(new_n843), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n915), .A2(new_n912), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT104), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n433), .A2(new_n926), .A3(new_n697), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n926), .B1(new_n433), .B2(new_n697), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n434), .A2(new_n930), .A3(new_n438), .ZN(new_n931));
  INV_X1    g0731(.A(new_n929), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n927), .ZN(new_n933));
  INV_X1    g0733(.A(new_n438), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n933), .B1(new_n650), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n924), .A2(new_n925), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n919), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n440), .B1(new_n757), .B2(new_n765), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n656), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n939), .B(new_n941), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n931), .A2(new_n935), .A3(new_n851), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n750), .A2(new_n752), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n743), .A2(new_n745), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n742), .A2(KEYINPUT31), .A3(new_n697), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n943), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n925), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT40), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n899), .B2(new_n912), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n949), .A2(new_n950), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n947), .A2(new_n440), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n953), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n954), .A2(G330), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n889), .B1(new_n942), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n942), .B2(new_n956), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n477), .B(KEYINPUT101), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT35), .ZN(new_n961));
  OAI211_X1 g0761(.A(G116), .B(new_n227), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(new_n961), .B2(new_n960), .ZN(new_n963));
  XNOR2_X1  g0763(.A(KEYINPUT102), .B(KEYINPUT36), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n963), .B(new_n964), .ZN(new_n965));
  NOR3_X1   g0765(.A1(new_n228), .A2(new_n217), .A3(new_n335), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n334), .A2(G50), .ZN(new_n967));
  OAI211_X1 g0767(.A(G1), .B(new_n557), .C1(new_n966), .C2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n958), .A2(new_n965), .A3(new_n968), .ZN(G367));
  NAND2_X1  g0769(.A1(new_n777), .A2(new_n238), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n212), .B2(new_n322), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n864), .A2(G143), .B1(G77), .B2(new_n817), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n333), .B2(new_n813), .C1(new_n830), .C2(new_n807), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n271), .B1(new_n792), .B2(new_n868), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(G68), .B2(new_n826), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n975), .B1(new_n256), .B2(new_n799), .C1(new_n828), .C2(new_n252), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n863), .A2(G294), .B1(G97), .B2(new_n817), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n800), .B2(new_n806), .ZN(new_n978));
  AOI22_X1  g0778(.A1(G283), .A2(new_n859), .B1(new_n803), .B2(G303), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n814), .A2(KEYINPUT46), .A3(G116), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n796), .A2(new_n205), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n363), .B(new_n981), .C1(G317), .C2(new_n793), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT46), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n813), .B2(new_n581), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n979), .A2(new_n980), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n973), .A2(new_n976), .B1(new_n978), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT47), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n838), .B1(new_n986), .B2(new_n987), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n771), .B1(new_n788), .B2(new_n971), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n665), .A2(new_n536), .A3(new_n698), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n536), .A2(new_n698), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n991), .B1(new_n678), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n786), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n990), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n766), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n486), .A2(new_n698), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n680), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n685), .A2(new_n697), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n712), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT44), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT108), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n705), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n712), .A2(new_n1001), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT45), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1003), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n705), .A2(new_n1004), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n709), .B1(new_n704), .B2(new_n708), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(new_n702), .Z(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n997), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n715), .B(new_n1018), .Z(new_n1019));
  OAI21_X1  g0819(.A(new_n769), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n999), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n685), .B1(new_n1021), .B2(new_n711), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n709), .B1(new_n999), .B2(new_n1000), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT42), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n1022), .A2(new_n697), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT43), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n1025), .A2(new_n1026), .B1(new_n1027), .B2(new_n994), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n994), .A2(new_n1027), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n705), .A2(new_n1001), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(KEYINPUT105), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1030), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1031), .A2(KEYINPUT105), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT106), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1034), .B(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n996), .B1(new_n1020), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(G387));
  OR2_X1    g0839(.A1(new_n704), .A2(new_n786), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n774), .A2(new_n717), .B1(G107), .B2(new_n212), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n235), .A2(G45), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n717), .ZN(new_n1043));
  AOI211_X1 g0843(.A(G45), .B(new_n1043), .C1(G68), .C2(G77), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n250), .A2(G50), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT50), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n778), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1041), .B1(new_n1042), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n771), .B1(new_n1048), .B2(new_n788), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT109), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n814), .A2(G77), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n807), .B2(new_n250), .C1(new_n830), .C2(new_n806), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n826), .A2(new_n494), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1053), .B(new_n363), .C1(new_n252), .C2(new_n792), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n828), .A2(new_n256), .B1(new_n334), .B2(new_n799), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n1052), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n204), .B2(new_n819), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G303), .A2(new_n859), .B1(new_n803), .B2(G317), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(KEYINPUT110), .B(G322), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1058), .B1(new_n800), .B2(new_n807), .C1(new_n806), .C2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT48), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n814), .A2(G294), .B1(G283), .B2(new_n826), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT111), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1067), .A2(KEYINPUT49), .A3(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n356), .B1(new_n805), .B2(new_n792), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n817), .B2(G116), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(KEYINPUT49), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1057), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1050), .B1(new_n1074), .B2(new_n838), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1075), .A2(KEYINPUT112), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT112), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1077), .B(new_n1050), .C1(new_n1074), .C2(new_n838), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1040), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(KEYINPUT113), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT113), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1081), .B(new_n1040), .C1(new_n1076), .C2(new_n1078), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1080), .A2(new_n1082), .B1(new_n770), .B2(new_n1016), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n997), .A2(new_n1015), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n766), .A2(new_n1016), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1084), .A2(new_n715), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1083), .A2(new_n1086), .ZN(G393));
  INV_X1    g0887(.A(new_n1010), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1009), .B(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1089), .A2(new_n1085), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1090), .A2(new_n716), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1085), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n769), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n999), .A2(new_n995), .A3(new_n1000), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n828), .A2(new_n830), .B1(new_n252), .B2(new_n806), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT51), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n813), .A2(new_n334), .B1(new_n807), .B2(new_n256), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n799), .A2(new_n250), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n826), .A2(G77), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n793), .A2(G143), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1100), .A2(new_n363), .A3(new_n1101), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n1098), .A2(new_n1099), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1097), .A2(new_n861), .A3(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n813), .A2(new_n820), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1059), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n271), .B1(new_n793), .B2(new_n1106), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1107), .B1(new_n581), .B2(new_n796), .C1(new_n799), .C2(new_n601), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1105), .B(new_n1108), .C1(G303), .C2(new_n863), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n864), .A2(G317), .B1(new_n803), .B2(G311), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1110), .B(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1109), .A2(new_n1112), .A3(new_n822), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n783), .B1(new_n1104), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n243), .A2(new_n778), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n1115), .B(new_n788), .C1(G97), .C2(new_n714), .ZN(new_n1116));
  NOR3_X1   g0916(.A1(new_n1114), .A2(new_n1116), .A3(new_n880), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1095), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(KEYINPUT115), .B1(new_n1094), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT115), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1121), .B(new_n1118), .C1(new_n1089), .C2(new_n769), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1093), .A2(new_n1123), .ZN(G390));
  NAND3_X1  g0924(.A1(new_n943), .A2(new_n947), .A3(G330), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT116), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n943), .A2(new_n947), .A3(KEYINPUT116), .A4(G330), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AND3_X1   g0929(.A1(new_n852), .A2(new_n922), .A3(new_n843), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n922), .B1(new_n852), .B2(new_n843), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n937), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n918), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n917), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n899), .A2(new_n912), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n1133), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n764), .A2(new_n698), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n843), .B1(new_n1137), .B2(new_n849), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1136), .B1(new_n1138), .B2(new_n937), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1129), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1139), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n744), .B1(new_n743), .B2(new_n745), .ZN(new_n1142));
  AOI211_X1 g0942(.A(KEYINPUT91), .B(KEYINPUT31), .C1(new_n742), .C2(new_n697), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n753), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1144), .A2(G330), .A3(new_n943), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(KEYINPUT117), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT117), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1144), .A2(new_n1147), .A3(G330), .A4(new_n943), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n918), .B1(new_n924), .B2(new_n937), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1141), .B(new_n1149), .C1(new_n1150), .C2(new_n917), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1140), .A2(new_n1151), .A3(new_n770), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(KEYINPUT121), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT121), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1140), .A2(new_n1151), .A3(new_n1154), .A4(new_n770), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n880), .B1(new_n884), .B2(new_n250), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n271), .B1(new_n793), .B2(G294), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1100), .B(new_n1158), .C1(new_n828), .C2(new_n581), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n823), .B1(new_n807), .B2(new_n205), .C1(new_n820), .C2(new_n806), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1159), .B(new_n1160), .C1(G97), .C2(new_n859), .ZN(new_n1161));
  XOR2_X1   g0961(.A(KEYINPUT54), .B(G143), .Z(new_n1162));
  NAND2_X1  g0962(.A1(new_n859), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n575), .B1(new_n793), .B2(G125), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1163), .B(new_n1164), .C1(new_n830), .C2(new_n796), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n864), .A2(G128), .B1(G50), .B2(new_n817), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n868), .B2(new_n807), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1165), .B(new_n1167), .C1(G132), .C2(new_n803), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n813), .A2(new_n252), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT53), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1161), .A2(new_n872), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1157), .B1(new_n783), .B2(new_n1171), .C1(new_n917), .C2(new_n881), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1138), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT119), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n947), .A2(new_n1174), .A3(G330), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n851), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1174), .B1(new_n947), .B2(G330), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n936), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1144), .A2(G330), .A3(new_n851), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n936), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1180), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1173), .A2(new_n1178), .B1(new_n1181), .B2(new_n924), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n947), .A2(new_n440), .A3(G330), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(KEYINPUT118), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT118), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n947), .A2(new_n440), .A3(new_n1185), .A4(G330), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1187), .A2(new_n940), .A3(new_n656), .ZN(new_n1188));
  OAI21_X1  g0988(.A(KEYINPUT120), .B1(new_n1182), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1138), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1149), .A2(new_n1178), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n937), .B1(new_n754), .B2(new_n851), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n924), .B1(new_n1129), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1191), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT120), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1188), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1189), .A2(new_n1197), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1140), .A2(new_n1151), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n715), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1140), .A2(new_n1151), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n1197), .B2(new_n1189), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1156), .B(new_n1172), .C1(new_n1200), .C2(new_n1202), .ZN(G378));
  NAND2_X1  g1003(.A1(new_n949), .A2(new_n950), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n948), .A2(new_n951), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(G330), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n297), .A2(new_n303), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n265), .A2(new_n890), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1207), .B(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1209), .B(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1206), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n952), .A2(G330), .A3(new_n1211), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n939), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1213), .A2(new_n938), .A3(new_n919), .A4(new_n1214), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1212), .A2(new_n784), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n771), .B1(new_n883), .B2(G50), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n799), .A2(new_n868), .B1(new_n252), .B2(new_n796), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n814), .A2(new_n1162), .B1(new_n864), .B2(G125), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n873), .B2(new_n807), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1221), .B(new_n1223), .C1(G128), .C2(new_n803), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n817), .A2(G159), .ZN(new_n1228));
  AOI211_X1 g1028(.A(G33), .B(G41), .C1(new_n793), .C2(G124), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n864), .A2(G116), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n863), .A2(G97), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n817), .A2(G58), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1051), .A2(new_n1231), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n826), .A2(G68), .B1(G283), .B2(new_n793), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n828), .B2(new_n205), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n283), .B(new_n356), .C1(new_n799), .C2(new_n322), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1234), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(KEYINPUT58), .ZN(new_n1239));
  OR2_X1    g1039(.A1(new_n1238), .A2(KEYINPUT58), .ZN(new_n1240));
  AOI21_X1  g1040(.A(G50), .B1(new_n268), .B2(new_n283), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n363), .B2(G41), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1230), .A2(new_n1239), .A3(new_n1240), .A4(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1220), .B1(new_n1243), .B2(new_n838), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(new_n1218), .A2(new_n770), .B1(new_n1219), .B2(new_n1244), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1188), .B(KEYINPUT122), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1195), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1247));
  AOI211_X1 g1047(.A(KEYINPUT120), .B(new_n1188), .C1(new_n1191), .C2(new_n1193), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1246), .B1(new_n1249), .B2(new_n1201), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT57), .B1(new_n1250), .B2(new_n1218), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1246), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1218), .A2(KEYINPUT57), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n715), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1245), .B1(new_n1251), .B2(new_n1255), .ZN(G375));
  NOR2_X1   g1056(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1198), .A2(new_n1019), .A3(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n880), .B1(new_n884), .B2(new_n334), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n271), .B1(new_n793), .B2(G303), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1053), .B(new_n1260), .C1(new_n828), .C2(new_n820), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(G116), .A2(new_n863), .B1(new_n864), .B2(G294), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n204), .B2(new_n813), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n1261), .B(new_n1263), .C1(G107), .C2(new_n859), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n818), .A2(G77), .ZN(new_n1265));
  INV_X1    g1065(.A(G128), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n363), .B1(new_n1266), .B2(new_n792), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n828), .A2(new_n868), .B1(new_n252), .B2(new_n799), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n1267), .B(new_n1268), .C1(G50), .C2(new_n826), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(G132), .A2(new_n864), .B1(new_n863), .B2(new_n1162), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n814), .A2(G159), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1270), .A2(new_n1233), .A3(new_n1271), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1264), .A2(new_n1265), .B1(new_n1269), .B2(new_n1272), .ZN(new_n1273));
  OAI221_X1 g1073(.A(new_n1259), .B1(new_n783), .B2(new_n1273), .C1(new_n937), .C2(new_n881), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(new_n1182), .B2(new_n769), .ZN(new_n1275));
  OR2_X1    g1075(.A1(new_n1258), .A2(new_n1275), .ZN(G381));
  NAND3_X1  g1076(.A1(new_n1083), .A2(new_n841), .A3(new_n1086), .ZN(new_n1277));
  OR3_X1    g1077(.A1(G381), .A2(G384), .A3(new_n1277), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n1091), .A2(new_n1092), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1038), .A2(new_n1279), .ZN(new_n1280));
  NOR4_X1   g1080(.A1(new_n1278), .A2(G375), .A3(G378), .A4(new_n1280), .ZN(new_n1281));
  XOR2_X1   g1081(.A(new_n1281), .B(KEYINPUT123), .Z(G407));
  INV_X1    g1082(.A(G378), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n696), .ZN(new_n1284));
  OAI211_X1 g1084(.A(G407), .B(G213), .C1(G375), .C2(new_n1284), .ZN(G409));
  NAND2_X1  g1085(.A1(G393), .A2(G396), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1277), .ZN(new_n1287));
  AOI22_X1  g1087(.A1(new_n1038), .A2(new_n1279), .B1(new_n1287), .B2(KEYINPUT126), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1020), .A2(new_n1037), .ZN(new_n1289));
  OAI21_X1  g1089(.A(G390), .B1(new_n1289), .B2(new_n996), .ZN(new_n1290));
  OR2_X1    g1090(.A1(new_n1287), .A2(KEYINPUT126), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1288), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1291), .B1(new_n1288), .B2(new_n1290), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  OAI211_X1 g1095(.A(G378), .B(new_n1245), .C1(new_n1251), .C2(new_n1255), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1172), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n716), .B1(new_n1249), .B2(new_n1201), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1297), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1301));
  NOR3_X1   g1101(.A1(new_n1253), .A2(new_n1019), .A3(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1245), .ZN(new_n1303));
  OAI211_X1 g1103(.A(new_n1300), .B(new_n1156), .C1(new_n1302), .C2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1296), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(G213), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1306), .A2(G343), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1275), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT60), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1182), .A2(new_n1188), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1310), .B1(new_n1249), .B2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n715), .B1(new_n1257), .B2(KEYINPUT60), .ZN(new_n1313));
  OAI211_X1 g1113(.A(G384), .B(new_n1309), .C1(new_n1312), .C2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1189), .A2(new_n1197), .A3(new_n1311), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1313), .B1(KEYINPUT60), .B2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n887), .B1(new_n1316), .B2(new_n1275), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1314), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1305), .A2(new_n1308), .A3(new_n1319), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(new_n1320), .B(KEYINPUT62), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1305), .A2(new_n1308), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1314), .A2(new_n1317), .A3(KEYINPUT125), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1307), .A2(G2897), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT125), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1318), .A2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1318), .A2(new_n1326), .A3(new_n1324), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1322), .A2(new_n1328), .A3(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT61), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1295), .B1(new_n1321), .B2(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1307), .B1(new_n1296), .B2(new_n1304), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1334), .A2(KEYINPUT63), .A3(new_n1319), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1330), .A2(new_n1331), .A3(new_n1294), .A4(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT63), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1320), .A2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(KEYINPUT124), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT124), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1320), .A2(new_n1341), .A3(new_n1338), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1340), .A2(new_n1342), .ZN(new_n1343));
  AOI21_X1  g1143(.A(KEYINPUT127), .B1(new_n1337), .B2(new_n1343), .ZN(new_n1344));
  AOI211_X1 g1144(.A(KEYINPUT124), .B(KEYINPUT63), .C1(new_n1334), .C2(new_n1319), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1341), .B1(new_n1320), .B2(new_n1338), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT127), .ZN(new_n1348));
  NOR3_X1   g1148(.A1(new_n1347), .A2(new_n1336), .A3(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1333), .B1(new_n1344), .B2(new_n1349), .ZN(G405));
  NAND2_X1  g1150(.A1(G375), .A2(new_n1283), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(new_n1296), .ZN(new_n1352));
  XNOR2_X1  g1152(.A(new_n1352), .B(new_n1319), .ZN(new_n1353));
  XNOR2_X1  g1153(.A(new_n1353), .B(new_n1295), .ZN(G402));
endmodule


