

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U324 ( .A(n461), .B(n460), .ZN(n572) );
  XNOR2_X1 U325 ( .A(n381), .B(n380), .ZN(n386) );
  NAND2_X1 U326 ( .A1(G227GAT), .A2(G233GAT), .ZN(n292) );
  XOR2_X1 U327 ( .A(KEYINPUT45), .B(n396), .Z(n293) );
  INV_X1 U328 ( .A(KEYINPUT114), .ZN(n399) );
  INV_X1 U329 ( .A(KEYINPUT9), .ZN(n378) );
  XNOR2_X1 U330 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U331 ( .A(n435), .B(n292), .ZN(n436) );
  INV_X1 U332 ( .A(KEYINPUT94), .ZN(n458) );
  XNOR2_X1 U333 ( .A(n437), .B(n436), .ZN(n439) );
  XNOR2_X1 U334 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U335 ( .A(KEYINPUT104), .B(KEYINPUT37), .ZN(n475) );
  XNOR2_X1 U336 ( .A(n557), .B(n395), .ZN(n585) );
  XNOR2_X1 U337 ( .A(n476), .B(n475), .ZN(n515) );
  INV_X1 U338 ( .A(G190GAT), .ZN(n451) );
  XNOR2_X1 U339 ( .A(n447), .B(n446), .ZN(n531) );
  XNOR2_X1 U340 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U341 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n480) );
  XNOR2_X1 U342 ( .A(n454), .B(n453), .ZN(G1351GAT) );
  XNOR2_X1 U343 ( .A(n481), .B(n480), .ZN(G1330GAT) );
  XOR2_X1 U344 ( .A(KEYINPUT89), .B(KEYINPUT82), .Z(n295) );
  XNOR2_X1 U345 ( .A(KEYINPUT24), .B(KEYINPUT88), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U347 ( .A(KEYINPUT23), .B(n296), .Z(n298) );
  NAND2_X1 U348 ( .A1(G228GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U349 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U350 ( .A(n299), .B(KEYINPUT22), .Z(n304) );
  XOR2_X1 U351 ( .A(KEYINPUT2), .B(G162GAT), .Z(n301) );
  XNOR2_X1 U352 ( .A(KEYINPUT86), .B(G155GAT), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U354 ( .A(KEYINPUT3), .B(n302), .Z(n430) );
  XNOR2_X1 U355 ( .A(n430), .B(KEYINPUT87), .ZN(n303) );
  XNOR2_X1 U356 ( .A(n304), .B(n303), .ZN(n307) );
  XOR2_X1 U357 ( .A(G78GAT), .B(G148GAT), .Z(n306) );
  XNOR2_X1 U358 ( .A(G106GAT), .B(G204GAT), .ZN(n305) );
  XNOR2_X1 U359 ( .A(n306), .B(n305), .ZN(n348) );
  XNOR2_X1 U360 ( .A(n307), .B(n348), .ZN(n315) );
  XNOR2_X1 U361 ( .A(G50GAT), .B(G22GAT), .ZN(n308) );
  XNOR2_X1 U362 ( .A(n308), .B(G141GAT), .ZN(n336) );
  XOR2_X1 U363 ( .A(KEYINPUT84), .B(KEYINPUT21), .Z(n310) );
  XNOR2_X1 U364 ( .A(G218GAT), .B(KEYINPUT83), .ZN(n309) );
  XNOR2_X1 U365 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U366 ( .A(n311), .B(KEYINPUT85), .Z(n313) );
  XNOR2_X1 U367 ( .A(G197GAT), .B(G211GAT), .ZN(n312) );
  XNOR2_X1 U368 ( .A(n313), .B(n312), .ZN(n327) );
  XOR2_X1 U369 ( .A(n336), .B(n327), .Z(n314) );
  XNOR2_X1 U370 ( .A(n315), .B(n314), .ZN(n467) );
  XOR2_X1 U371 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n317) );
  XNOR2_X1 U372 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n317), .B(n316), .ZN(n433) );
  XOR2_X1 U374 ( .A(G92GAT), .B(G64GAT), .Z(n347) );
  XOR2_X1 U375 ( .A(n433), .B(n347), .Z(n319) );
  NAND2_X1 U376 ( .A1(G226GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U377 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U378 ( .A(KEYINPUT74), .B(KEYINPUT93), .Z(n321) );
  XNOR2_X1 U379 ( .A(G8GAT), .B(G204GAT), .ZN(n320) );
  XNOR2_X1 U380 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U381 ( .A(n323), .B(n322), .Z(n329) );
  XOR2_X1 U382 ( .A(G190GAT), .B(G183GAT), .Z(n325) );
  XNOR2_X1 U383 ( .A(G36GAT), .B(G176GAT), .ZN(n324) );
  XNOR2_X1 U384 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U385 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n457) );
  XNOR2_X1 U387 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n409) );
  XOR2_X1 U388 ( .A(KEYINPUT30), .B(G197GAT), .Z(n331) );
  XNOR2_X1 U389 ( .A(G169GAT), .B(G113GAT), .ZN(n330) );
  XNOR2_X1 U390 ( .A(n331), .B(n330), .ZN(n340) );
  XOR2_X1 U391 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n333) );
  NAND2_X1 U392 ( .A1(G229GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U393 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U394 ( .A(n334), .B(KEYINPUT29), .Z(n338) );
  XNOR2_X1 U395 ( .A(G15GAT), .B(G8GAT), .ZN(n335) );
  XNOR2_X1 U396 ( .A(n335), .B(G1GAT), .ZN(n368) );
  XNOR2_X1 U397 ( .A(n336), .B(n368), .ZN(n337) );
  XNOR2_X1 U398 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U399 ( .A(n340), .B(n339), .ZN(n345) );
  XOR2_X1 U400 ( .A(G29GAT), .B(KEYINPUT8), .Z(n342) );
  XNOR2_X1 U401 ( .A(G43GAT), .B(G36GAT), .ZN(n341) );
  XNOR2_X1 U402 ( .A(n342), .B(n341), .ZN(n344) );
  XOR2_X1 U403 ( .A(KEYINPUT68), .B(KEYINPUT7), .Z(n343) );
  XNOR2_X1 U404 ( .A(n344), .B(n343), .ZN(n391) );
  XOR2_X1 U405 ( .A(n345), .B(n391), .Z(n547) );
  INV_X1 U406 ( .A(n547), .ZN(n574) );
  XOR2_X1 U407 ( .A(KEYINPUT69), .B(n574), .Z(n560) );
  INV_X1 U408 ( .A(n560), .ZN(n534) );
  XNOR2_X1 U409 ( .A(G71GAT), .B(G57GAT), .ZN(n346) );
  XNOR2_X1 U410 ( .A(n346), .B(KEYINPUT13), .ZN(n360) );
  XOR2_X1 U411 ( .A(n360), .B(n347), .Z(n350) );
  XOR2_X1 U412 ( .A(G176GAT), .B(G120GAT), .Z(n445) );
  XNOR2_X1 U413 ( .A(n445), .B(n348), .ZN(n349) );
  XNOR2_X1 U414 ( .A(n350), .B(n349), .ZN(n357) );
  XOR2_X1 U415 ( .A(G99GAT), .B(G85GAT), .Z(n377) );
  XOR2_X1 U416 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n352) );
  XNOR2_X1 U417 ( .A(KEYINPUT70), .B(KEYINPUT31), .ZN(n351) );
  XNOR2_X1 U418 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U419 ( .A(n377), .B(n353), .Z(n355) );
  NAND2_X1 U420 ( .A1(G230GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U421 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U422 ( .A(n357), .B(n356), .Z(n477) );
  XOR2_X1 U423 ( .A(KEYINPUT15), .B(KEYINPUT77), .Z(n363) );
  XOR2_X1 U424 ( .A(KEYINPUT14), .B(KEYINPUT75), .Z(n359) );
  XNOR2_X1 U425 ( .A(KEYINPUT12), .B(KEYINPUT76), .ZN(n358) );
  XNOR2_X1 U426 ( .A(n359), .B(n358), .ZN(n361) );
  XNOR2_X1 U427 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U429 ( .A(G78GAT), .B(G155GAT), .Z(n365) );
  XNOR2_X1 U430 ( .A(G22GAT), .B(G211GAT), .ZN(n364) );
  XNOR2_X1 U431 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U432 ( .A(n367), .B(n366), .Z(n376) );
  XOR2_X1 U433 ( .A(G183GAT), .B(G127GAT), .Z(n444) );
  XOR2_X1 U434 ( .A(n444), .B(n368), .Z(n370) );
  NAND2_X1 U435 ( .A1(G231GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U436 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U437 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n372) );
  XNOR2_X1 U438 ( .A(KEYINPUT74), .B(G64GAT), .ZN(n371) );
  XNOR2_X1 U439 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U440 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U441 ( .A(n376), .B(n375), .ZN(n582) );
  XOR2_X1 U442 ( .A(G190GAT), .B(G134GAT), .Z(n434) );
  XNOR2_X1 U443 ( .A(n434), .B(n377), .ZN(n381) );
  XOR2_X1 U444 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n379) );
  XOR2_X1 U445 ( .A(G92GAT), .B(G106GAT), .Z(n383) );
  XNOR2_X1 U446 ( .A(G50GAT), .B(G162GAT), .ZN(n382) );
  XNOR2_X1 U447 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U448 ( .A(G218GAT), .B(n384), .ZN(n385) );
  XNOR2_X1 U449 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U450 ( .A(KEYINPUT71), .B(KEYINPUT73), .Z(n388) );
  NAND2_X1 U451 ( .A1(G232GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U452 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U453 ( .A(n390), .B(n389), .ZN(n394) );
  INV_X1 U454 ( .A(n391), .ZN(n392) );
  XOR2_X1 U455 ( .A(n392), .B(KEYINPUT72), .Z(n393) );
  XNOR2_X2 U456 ( .A(n394), .B(n393), .ZN(n557) );
  XNOR2_X1 U457 ( .A(KEYINPUT36), .B(KEYINPUT103), .ZN(n395) );
  NOR2_X1 U458 ( .A1(n582), .A2(n585), .ZN(n396) );
  NOR2_X1 U459 ( .A1(n477), .A2(n293), .ZN(n397) );
  XNOR2_X1 U460 ( .A(n397), .B(KEYINPUT113), .ZN(n398) );
  NOR2_X1 U461 ( .A1(n534), .A2(n398), .ZN(n400) );
  XNOR2_X1 U462 ( .A(n400), .B(n399), .ZN(n407) );
  XNOR2_X1 U463 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n401) );
  INV_X1 U464 ( .A(n477), .ZN(n579) );
  XNOR2_X1 U465 ( .A(n401), .B(n579), .ZN(n549) );
  NAND2_X1 U466 ( .A1(n547), .A2(n549), .ZN(n402) );
  XNOR2_X1 U467 ( .A(n402), .B(KEYINPUT46), .ZN(n403) );
  XNOR2_X1 U468 ( .A(KEYINPUT112), .B(n582), .ZN(n568) );
  NAND2_X1 U469 ( .A1(n403), .A2(n568), .ZN(n404) );
  NOR2_X1 U470 ( .A1(n557), .A2(n404), .ZN(n405) );
  XNOR2_X1 U471 ( .A(KEYINPUT47), .B(n405), .ZN(n406) );
  NAND2_X1 U472 ( .A1(n407), .A2(n406), .ZN(n408) );
  XNOR2_X1 U473 ( .A(n409), .B(n408), .ZN(n528) );
  NOR2_X1 U474 ( .A1(n457), .A2(n528), .ZN(n411) );
  XNOR2_X1 U475 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n410) );
  XNOR2_X1 U476 ( .A(n411), .B(n410), .ZN(n431) );
  XOR2_X1 U477 ( .A(G57GAT), .B(G148GAT), .Z(n413) );
  XNOR2_X1 U478 ( .A(G141GAT), .B(G127GAT), .ZN(n412) );
  XNOR2_X1 U479 ( .A(n413), .B(n412), .ZN(n417) );
  XOR2_X1 U480 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n415) );
  XNOR2_X1 U481 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n414) );
  XNOR2_X1 U482 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U483 ( .A(n417), .B(n416), .Z(n428) );
  XOR2_X1 U484 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n419) );
  XNOR2_X1 U485 ( .A(KEYINPUT6), .B(KEYINPUT90), .ZN(n418) );
  XNOR2_X1 U486 ( .A(n419), .B(n418), .ZN(n426) );
  XOR2_X1 U487 ( .A(G113GAT), .B(KEYINPUT0), .Z(n435) );
  XOR2_X1 U488 ( .A(G85GAT), .B(G134GAT), .Z(n421) );
  XNOR2_X1 U489 ( .A(G29GAT), .B(G120GAT), .ZN(n420) );
  XNOR2_X1 U490 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U491 ( .A(n435), .B(n422), .Z(n424) );
  NAND2_X1 U492 ( .A1(G225GAT), .A2(G233GAT), .ZN(n423) );
  XNOR2_X1 U493 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U494 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U495 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U496 ( .A(n430), .B(n429), .ZN(n517) );
  NOR2_X1 U497 ( .A1(n431), .A2(n517), .ZN(n573) );
  NAND2_X1 U498 ( .A1(n467), .A2(n573), .ZN(n432) );
  XNOR2_X1 U499 ( .A(n432), .B(KEYINPUT55), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n434), .B(n433), .ZN(n437) );
  XNOR2_X1 U501 ( .A(G43GAT), .B(G99GAT), .ZN(n438) );
  XNOR2_X1 U502 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U503 ( .A(G71GAT), .B(KEYINPUT80), .Z(n441) );
  XNOR2_X1 U504 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n440) );
  XNOR2_X1 U505 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U506 ( .A(n443), .B(n442), .ZN(n447) );
  XOR2_X1 U507 ( .A(n445), .B(n444), .Z(n446) );
  NAND2_X1 U508 ( .A1(n448), .A2(n531), .ZN(n449) );
  XNOR2_X1 U509 ( .A(KEYINPUT122), .B(n449), .ZN(n569) );
  INV_X1 U510 ( .A(n557), .ZN(n450) );
  NOR2_X1 U511 ( .A1(n569), .A2(n450), .ZN(n454) );
  XNOR2_X1 U512 ( .A(KEYINPUT58), .B(KEYINPUT126), .ZN(n452) );
  INV_X1 U513 ( .A(n457), .ZN(n519) );
  NAND2_X1 U514 ( .A1(n531), .A2(n519), .ZN(n455) );
  NAND2_X1 U515 ( .A1(n467), .A2(n455), .ZN(n456) );
  XNOR2_X1 U516 ( .A(KEYINPUT25), .B(n456), .ZN(n464) );
  XOR2_X1 U517 ( .A(n457), .B(KEYINPUT27), .Z(n466) );
  NOR2_X1 U518 ( .A1(n531), .A2(n467), .ZN(n461) );
  XNOR2_X1 U519 ( .A(KEYINPUT95), .B(KEYINPUT26), .ZN(n459) );
  AND2_X1 U520 ( .A1(n466), .A2(n572), .ZN(n462) );
  XNOR2_X1 U521 ( .A(n462), .B(KEYINPUT96), .ZN(n463) );
  NOR2_X1 U522 ( .A1(n464), .A2(n463), .ZN(n465) );
  NOR2_X1 U523 ( .A1(n465), .A2(n517), .ZN(n472) );
  NAND2_X1 U524 ( .A1(n466), .A2(n517), .ZN(n527) );
  XNOR2_X1 U525 ( .A(KEYINPUT81), .B(n531), .ZN(n469) );
  XOR2_X1 U526 ( .A(n467), .B(KEYINPUT28), .Z(n468) );
  XNOR2_X1 U527 ( .A(KEYINPUT65), .B(n468), .ZN(n530) );
  NAND2_X1 U528 ( .A1(n469), .A2(n530), .ZN(n470) );
  NOR2_X1 U529 ( .A1(n527), .A2(n470), .ZN(n471) );
  NOR2_X1 U530 ( .A1(n472), .A2(n471), .ZN(n473) );
  XOR2_X1 U531 ( .A(KEYINPUT97), .B(n473), .Z(n484) );
  NOR2_X1 U532 ( .A1(n585), .A2(n484), .ZN(n474) );
  NAND2_X1 U533 ( .A1(n474), .A2(n582), .ZN(n476) );
  NOR2_X1 U534 ( .A1(n477), .A2(n560), .ZN(n485) );
  NAND2_X1 U535 ( .A1(n515), .A2(n485), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n478), .B(KEYINPUT38), .ZN(n479) );
  XNOR2_X1 U537 ( .A(KEYINPUT105), .B(n479), .ZN(n502) );
  NAND2_X1 U538 ( .A1(n502), .A2(n531), .ZN(n481) );
  NOR2_X1 U539 ( .A1(n557), .A2(n582), .ZN(n482) );
  XOR2_X1 U540 ( .A(KEYINPUT16), .B(n482), .Z(n483) );
  NOR2_X1 U541 ( .A1(n484), .A2(n483), .ZN(n504) );
  AND2_X1 U542 ( .A1(n485), .A2(n504), .ZN(n494) );
  NAND2_X1 U543 ( .A1(n494), .A2(n517), .ZN(n486) );
  XNOR2_X1 U544 ( .A(KEYINPUT34), .B(n486), .ZN(n487) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(n487), .ZN(G1324GAT) );
  NAND2_X1 U546 ( .A1(n519), .A2(n494), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n488), .B(KEYINPUT98), .ZN(n489) );
  XNOR2_X1 U548 ( .A(G8GAT), .B(n489), .ZN(G1325GAT) );
  XOR2_X1 U549 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n491) );
  NAND2_X1 U550 ( .A1(n494), .A2(n531), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(n493) );
  XOR2_X1 U552 ( .A(G15GAT), .B(KEYINPUT99), .Z(n492) );
  XNOR2_X1 U553 ( .A(n493), .B(n492), .ZN(G1326GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT101), .B(KEYINPUT102), .Z(n496) );
  INV_X1 U555 ( .A(n530), .ZN(n522) );
  NAND2_X1 U556 ( .A1(n494), .A2(n522), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U558 ( .A(G22GAT), .B(n497), .ZN(G1327GAT) );
  XOR2_X1 U559 ( .A(G29GAT), .B(KEYINPUT39), .Z(n499) );
  NAND2_X1 U560 ( .A1(n502), .A2(n517), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  NAND2_X1 U562 ( .A1(n502), .A2(n519), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n500), .B(KEYINPUT106), .ZN(n501) );
  XNOR2_X1 U564 ( .A(G36GAT), .B(n501), .ZN(G1329GAT) );
  NAND2_X1 U565 ( .A1(n522), .A2(n502), .ZN(n503) );
  XNOR2_X1 U566 ( .A(G50GAT), .B(n503), .ZN(G1331GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n507) );
  XNOR2_X1 U568 ( .A(KEYINPUT107), .B(n549), .ZN(n563) );
  NOR2_X1 U569 ( .A1(n547), .A2(n563), .ZN(n516) );
  NAND2_X1 U570 ( .A1(n504), .A2(n516), .ZN(n505) );
  XOR2_X1 U571 ( .A(KEYINPUT108), .B(n505), .Z(n512) );
  NAND2_X1 U572 ( .A1(n512), .A2(n517), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U574 ( .A(G57GAT), .B(n508), .ZN(G1332GAT) );
  NAND2_X1 U575 ( .A1(n512), .A2(n519), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n509), .B(KEYINPUT110), .ZN(n510) );
  XNOR2_X1 U577 ( .A(G64GAT), .B(n510), .ZN(G1333GAT) );
  NAND2_X1 U578 ( .A1(n512), .A2(n531), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n511), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U581 ( .A1(n522), .A2(n512), .ZN(n513) );
  XNOR2_X1 U582 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  AND2_X1 U583 ( .A1(n516), .A2(n515), .ZN(n523) );
  NAND2_X1 U584 ( .A1(n523), .A2(n517), .ZN(n518) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(n518), .ZN(G1336GAT) );
  NAND2_X1 U586 ( .A1(n519), .A2(n523), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n520), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n523), .A2(n531), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n521), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n525) );
  NAND2_X1 U591 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  NOR2_X1 U594 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U595 ( .A(KEYINPUT116), .B(n529), .Z(n546) );
  NAND2_X1 U596 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U597 ( .A1(n546), .A2(n532), .ZN(n533) );
  XOR2_X1 U598 ( .A(KEYINPUT117), .B(n533), .Z(n541) );
  NAND2_X1 U599 ( .A1(n534), .A2(n541), .ZN(n535) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(n535), .ZN(G1340GAT) );
  INV_X1 U601 ( .A(n541), .ZN(n538) );
  NOR2_X1 U602 ( .A1(n563), .A2(n538), .ZN(n537) );
  XNOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  NOR2_X1 U605 ( .A1(n568), .A2(n538), .ZN(n539) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(n539), .Z(n540) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U609 ( .A1(n541), .A2(n557), .ZN(n542) );
  XNOR2_X1 U610 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U611 ( .A(G134GAT), .B(n544), .ZN(G1343GAT) );
  INV_X1 U612 ( .A(n572), .ZN(n545) );
  NOR2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n558) );
  NAND2_X1 U614 ( .A1(n547), .A2(n558), .ZN(n548) );
  XNOR2_X1 U615 ( .A(G141GAT), .B(n548), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n551) );
  NAND2_X1 U617 ( .A1(n558), .A2(n549), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(n553) );
  XOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT53), .Z(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(KEYINPUT120), .ZN(n556) );
  INV_X1 U622 ( .A(n582), .ZN(n554) );
  NAND2_X1 U623 ( .A1(n558), .A2(n554), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(G1346GAT) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U627 ( .A1(n569), .A2(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(KEYINPUT123), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(G1348GAT) );
  XNOR2_X1 U630 ( .A(KEYINPUT57), .B(KEYINPUT124), .ZN(n567) );
  XNOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n565) );
  NOR2_X1 U632 ( .A1(n569), .A2(n563), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  NOR2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G183GAT), .B(KEYINPUT125), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(G1350GAT) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n584) );
  NOR2_X1 U639 ( .A1(n584), .A2(n574), .ZN(n578) );
  XOR2_X1 U640 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT127), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n584), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n584), .ZN(n583) );
  XOR2_X1 U648 ( .A(G211GAT), .B(n583), .Z(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(n586), .Z(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

