//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  INV_X1    g0013(.A(G97), .ZN(new_n214));
  INV_X1    g0014(.A(G257), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT65), .ZN(new_n217));
  AOI21_X1  g0017(.A(new_n210), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n218), .B1(new_n217), .B2(new_n216), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G20), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT66), .Z(new_n223));
  NOR2_X1   g0023(.A1(new_n220), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(G250), .B1(G257), .B2(G264), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n201), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI22_X1  g0033(.A1(new_n227), .A2(KEYINPUT0), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(new_n234), .B1(KEYINPUT0), .B2(new_n227), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT64), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n237));
  NOR3_X1   g0037(.A1(new_n223), .A2(new_n236), .A3(new_n237), .ZN(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G226), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G250), .B(G257), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G264), .B(G270), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n243), .B(new_n247), .ZN(G358));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT69), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G50), .B(G68), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G58), .B(G77), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  INV_X1    g0056(.A(G200), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  OAI211_X1 g0059(.A(G1), .B(G13), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G33), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n261), .A2(new_n263), .A3(G226), .A4(G1698), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT78), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT3), .B(G33), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT78), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n266), .A2(new_n267), .A3(G226), .A4(G1698), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G1698), .ZN(new_n270));
  AND3_X1   g0070(.A1(new_n261), .A2(new_n263), .A3(new_n270), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n271), .A2(G223), .B1(G33), .B2(G87), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n260), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G274), .ZN(new_n275));
  INV_X1    g0075(.A(G1), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n276), .B1(G41), .B2(G45), .ZN(new_n277));
  NOR3_X1   g0077(.A1(new_n274), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n277), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n274), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G232), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n257), .B1(new_n273), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G190), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n278), .B1(G232), .B2(new_n281), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n261), .A2(new_n263), .A3(G223), .A4(new_n270), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n287), .B1(new_n258), .B2(new_n212), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n288), .B1(new_n268), .B2(new_n265), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n285), .B(new_n286), .C1(new_n289), .C2(new_n260), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n261), .A2(new_n263), .ZN(new_n292));
  AOI21_X1  g0092(.A(KEYINPUT7), .B1(new_n292), .B2(new_n232), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT7), .ZN(new_n294));
  AOI211_X1 g0094(.A(new_n294), .B(G20), .C1(new_n261), .C2(new_n263), .ZN(new_n295));
  OAI21_X1  g0095(.A(G68), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G58), .ZN(new_n297));
  INV_X1    g0097(.A(G68), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(G20), .B1(new_n299), .B2(new_n201), .ZN(new_n300));
  NOR2_X1   g0100(.A1(G20), .A2(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G159), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n296), .A2(KEYINPUT16), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT16), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n294), .B1(new_n266), .B2(G20), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n292), .A2(KEYINPUT7), .A3(new_n232), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n298), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n306), .B1(new_n309), .B2(new_n303), .ZN(new_n310));
  NAND3_X1  g0110(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n231), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT70), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT70), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n311), .A2(new_n314), .A3(new_n231), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n305), .A2(new_n310), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G13), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n318), .A2(new_n232), .A3(G1), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT8), .B(G58), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n321), .B1(new_n276), .B2(G20), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n320), .A2(new_n322), .B1(new_n321), .B2(new_n319), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT79), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n291), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n320), .A2(new_n322), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n321), .A2(new_n319), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n313), .A2(new_n315), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n296), .A2(new_n304), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n330), .B1(new_n331), .B2(new_n306), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n329), .B1(new_n332), .B2(new_n305), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n284), .A2(new_n290), .ZN(new_n334));
  AOI21_X1  g0134(.A(KEYINPUT79), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(KEYINPUT17), .B1(new_n326), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(G169), .B1(new_n273), .B2(new_n283), .ZN(new_n337));
  INV_X1    g0137(.A(G179), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n286), .B1(new_n289), .B2(new_n260), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT18), .ZN(new_n341));
  AND3_X1   g0141(.A1(new_n340), .A2(new_n324), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n341), .B1(new_n340), .B2(new_n324), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n333), .A2(new_n334), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT17), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n336), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT80), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n348), .B(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n271), .A2(G222), .ZN(new_n351));
  INV_X1    g0151(.A(G77), .ZN(new_n352));
  INV_X1    g0152(.A(G223), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n266), .A2(G1698), .ZN(new_n354));
  OAI221_X1 g0154(.A(new_n351), .B1(new_n352), .B2(new_n266), .C1(new_n353), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n274), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n278), .B1(G226), .B2(new_n281), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(G169), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n319), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n276), .A2(G20), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n330), .A2(G50), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n203), .A2(G20), .ZN(new_n365));
  INV_X1    g0165(.A(G150), .ZN(new_n366));
  INV_X1    g0166(.A(new_n301), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n232), .A2(G33), .ZN(new_n368));
  OAI221_X1 g0168(.A(new_n365), .B1(new_n366), .B2(new_n367), .C1(new_n368), .C2(new_n321), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n369), .A2(new_n316), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n364), .B1(new_n370), .B2(KEYINPUT71), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n369), .A2(new_n316), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT71), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n372), .A2(new_n373), .B1(new_n202), .B2(new_n319), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n360), .B(new_n375), .C1(G179), .C2(new_n358), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(KEYINPUT9), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT9), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n371), .A2(new_n379), .A3(new_n374), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT76), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n358), .A2(new_n285), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n381), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n358), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(new_n257), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n382), .B1(new_n381), .B2(new_n384), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT10), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT10), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n358), .A2(KEYINPUT75), .A3(G200), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n384), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT75), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n394), .B1(new_n395), .B2(new_n388), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n381), .A2(KEYINPUT74), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n381), .A2(KEYINPUT74), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n377), .B1(new_n391), .B2(new_n399), .ZN(new_n400));
  AOI22_X1  g0200(.A1(new_n301), .A2(G50), .B1(G20), .B2(new_n298), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n352), .B2(new_n368), .ZN(new_n402));
  AND2_X1   g0202(.A1(new_n316), .A2(new_n402), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n403), .A2(KEYINPUT11), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n319), .A2(new_n298), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n405), .B(KEYINPUT12), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n403), .A2(KEYINPUT11), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n320), .A2(G68), .A3(new_n362), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n404), .A2(new_n406), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT14), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n271), .A2(G226), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n266), .A2(G232), .A3(G1698), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G97), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n274), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT13), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n278), .B1(G238), .B2(new_n281), .ZN(new_n417));
  AND3_X1   g0217(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n416), .B1(new_n415), .B2(new_n417), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n410), .B(G169), .C1(new_n418), .C2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n419), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n420), .B1(new_n423), .B2(new_n338), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n410), .B1(new_n423), .B2(G169), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n409), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n418), .A2(new_n419), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n409), .B1(new_n427), .B2(G190), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT77), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n423), .B2(G200), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n429), .B(G200), .C1(new_n418), .C2(new_n419), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n428), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n426), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(G238), .ZN(new_n435));
  INV_X1    g0235(.A(G107), .ZN(new_n436));
  OAI22_X1  g0236(.A1(new_n354), .A2(new_n435), .B1(new_n436), .B2(new_n266), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n266), .A2(G232), .A3(new_n270), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n274), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n278), .B1(G244), .B2(new_n281), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(G190), .ZN(new_n442));
  XOR2_X1   g0242(.A(new_n442), .B(KEYINPUT72), .Z(new_n443));
  AOI21_X1  g0243(.A(new_n321), .B1(KEYINPUT73), .B2(new_n367), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(KEYINPUT73), .B2(new_n367), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT15), .B(G87), .ZN(new_n446));
  OAI221_X1 g0246(.A(new_n445), .B1(new_n232), .B2(new_n352), .C1(new_n368), .C2(new_n446), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n447), .A2(new_n316), .B1(new_n352), .B2(new_n319), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n320), .A2(G77), .A3(new_n362), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n441), .A2(new_n257), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n443), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n441), .A2(new_n338), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n450), .B(new_n455), .C1(G169), .C2(new_n441), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n434), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n350), .A2(new_n400), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT81), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n350), .A2(new_n400), .A3(KEYINPUT81), .A4(new_n458), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G45), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(G1), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n466), .B(KEYINPUT84), .C1(KEYINPUT5), .C2(new_n259), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n276), .B(G45), .C1(new_n259), .C2(KEYINPUT5), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT84), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n259), .A2(KEYINPUT5), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n467), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(G264), .A3(new_n260), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n292), .A2(new_n215), .A3(new_n270), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n261), .A2(new_n263), .A3(G250), .A4(new_n270), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G294), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n274), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n468), .A2(new_n469), .B1(KEYINPUT5), .B2(new_n259), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n479), .A2(G274), .A3(new_n260), .A4(new_n467), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n473), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  OR2_X1    g0281(.A1(new_n481), .A2(G179), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n359), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n261), .A2(new_n263), .A3(new_n232), .A4(G87), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT22), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT22), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n266), .A2(new_n487), .A3(new_n232), .A4(G87), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G116), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n490), .A2(G20), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT23), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n232), .B2(G107), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n436), .A2(KEYINPUT23), .A3(G20), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT24), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT24), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n489), .A2(new_n498), .A3(new_n495), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n330), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n276), .A2(G33), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n330), .A2(new_n361), .A3(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(new_n436), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n319), .A2(new_n436), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n504), .B(KEYINPUT25), .ZN(new_n505));
  OR2_X1    g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n484), .A2(new_n507), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n489), .A2(new_n498), .A3(new_n495), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n498), .B1(new_n489), .B2(new_n495), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n316), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n481), .A2(G200), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n503), .A2(new_n505), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n473), .A2(new_n478), .A3(G190), .A4(new_n480), .ZN(new_n514));
  AND4_X1   g0314(.A1(new_n511), .A2(new_n512), .A3(new_n513), .A4(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n508), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n330), .A2(G116), .A3(new_n361), .A4(new_n501), .ZN(new_n517));
  INV_X1    g0317(.A(G116), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n319), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n311), .A2(new_n231), .B1(G20), .B2(new_n518), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G283), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n521), .B(new_n232), .C1(G33), .C2(new_n214), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT20), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n520), .A2(KEYINPUT20), .A3(new_n522), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n517), .B(new_n519), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n472), .A2(G270), .A3(new_n260), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n261), .A2(new_n263), .A3(G264), .A4(G1698), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n261), .A2(new_n263), .A3(G257), .A4(new_n270), .ZN(new_n528));
  INV_X1    g0328(.A(G303), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n527), .B(new_n528), .C1(new_n529), .C2(new_n266), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n274), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n526), .A2(new_n531), .A3(new_n480), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n525), .A2(new_n532), .A3(G169), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT21), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n532), .A2(G200), .ZN(new_n536));
  INV_X1    g0336(.A(new_n525), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n526), .A2(new_n531), .A3(G190), .A4(new_n480), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n526), .A2(new_n480), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n540), .A2(new_n525), .A3(G179), .A4(new_n531), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n525), .A2(new_n532), .A3(KEYINPUT21), .A4(G169), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n535), .A2(new_n539), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT88), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n541), .A2(new_n542), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n546), .A2(KEYINPUT88), .A3(new_n535), .A4(new_n539), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n361), .A2(G97), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(new_n502), .B2(new_n214), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n436), .B1(new_n307), .B2(new_n308), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n301), .A2(G77), .ZN(new_n553));
  NAND2_X1  g0353(.A1(KEYINPUT6), .A2(G97), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n554), .A2(G107), .ZN(new_n555));
  XNOR2_X1  g0355(.A(G97), .B(G107), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT6), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n553), .B1(new_n558), .B2(new_n232), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n316), .B1(new_n552), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT82), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(KEYINPUT82), .B(new_n316), .C1(new_n552), .C2(new_n559), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n551), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n271), .A2(KEYINPUT83), .A3(KEYINPUT4), .A4(G244), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n261), .A2(new_n263), .A3(G250), .A4(G1698), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n566), .A2(new_n521), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT83), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n261), .A2(new_n263), .A3(G244), .A4(new_n270), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT4), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n569), .A2(new_n570), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n565), .A2(new_n567), .A3(new_n571), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n274), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n274), .B1(new_n479), .B2(new_n467), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(G257), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n480), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G200), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n573), .A2(new_n274), .B1(G257), .B2(new_n575), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n579), .A2(G190), .A3(new_n480), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n564), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n551), .ZN(new_n582));
  OAI21_X1  g0382(.A(G107), .B1(new_n293), .B2(new_n295), .ZN(new_n583));
  AND2_X1   g0383(.A1(G97), .A2(G107), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n557), .B1(new_n584), .B2(new_n205), .ZN(new_n585));
  INV_X1    g0385(.A(new_n555), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n587), .A2(G20), .B1(G77), .B2(new_n301), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT82), .B1(new_n589), .B2(new_n316), .ZN(new_n590));
  AOI211_X1 g0390(.A(new_n561), .B(new_n330), .C1(new_n583), .C2(new_n588), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n582), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT85), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n564), .A2(KEYINPUT85), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n579), .A2(G179), .A3(new_n480), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n574), .A2(new_n480), .A3(new_n576), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n597), .B1(new_n598), .B2(new_n359), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n581), .B1(new_n596), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n502), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(G87), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n266), .A2(new_n232), .A3(G68), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT19), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n232), .B1(new_n413), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(G87), .B2(new_n206), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n604), .B1(new_n368), .B2(new_n214), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n603), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n608), .A2(new_n316), .B1(new_n319), .B2(new_n446), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n466), .A2(new_n275), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n213), .B1(new_n465), .B2(G1), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n260), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n266), .A2(G244), .A3(G1698), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n266), .A2(G238), .A3(new_n270), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n616), .A3(new_n490), .ZN(new_n617));
  AOI211_X1 g0417(.A(new_n285), .B(new_n614), .C1(new_n617), .C2(new_n274), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n610), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n274), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n613), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(G200), .ZN(new_n622));
  XOR2_X1   g0422(.A(new_n446), .B(KEYINPUT86), .Z(new_n623));
  NAND2_X1  g0423(.A1(new_n601), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n614), .B1(new_n617), .B2(new_n274), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n624), .A2(new_n609), .B1(new_n625), .B2(new_n338), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n621), .A2(new_n359), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n619), .A2(new_n622), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT87), .B1(new_n600), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n562), .A2(new_n563), .ZN(new_n630));
  AOI21_X1  g0430(.A(KEYINPUT85), .B1(new_n630), .B2(new_n582), .ZN(new_n631));
  AOI211_X1 g0431(.A(new_n593), .B(new_n551), .C1(new_n562), .C2(new_n563), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n599), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n564), .A2(new_n578), .A3(new_n580), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n633), .A2(KEYINPUT87), .A3(new_n628), .A4(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n516), .B(new_n548), .C1(new_n629), .C2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n464), .A2(new_n637), .ZN(G372));
  NAND2_X1  g0438(.A1(new_n624), .A2(new_n609), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n625), .A2(new_n338), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT89), .ZN(new_n642));
  XNOR2_X1  g0442(.A(new_n613), .B(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(G169), .B1(new_n643), .B2(new_n620), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n609), .B(new_n602), .C1(new_n621), .C2(new_n285), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n257), .B1(new_n643), .B2(new_n620), .ZN(new_n646));
  OAI22_X1  g0446(.A1(new_n641), .A2(new_n644), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n647), .A2(new_n515), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n633), .A2(new_n634), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT90), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n633), .A2(new_n648), .A3(KEYINPUT90), .A4(new_n634), .ZN(new_n652));
  INV_X1    g0452(.A(new_n508), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n653), .A2(new_n546), .A3(new_n535), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n651), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n646), .ZN(new_n656));
  INV_X1    g0456(.A(new_n644), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n619), .A2(new_n656), .B1(new_n626), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n658), .A2(new_n599), .A3(new_n659), .A4(new_n592), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n626), .A2(new_n657), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI211_X1 g0462(.A(new_n628), .B(new_n599), .C1(new_n631), .C2(new_n632), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n662), .B1(KEYINPUT26), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n655), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n463), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n433), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n426), .B1(new_n667), .B2(new_n456), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n668), .A2(new_n336), .A3(new_n347), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n344), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n391), .A2(new_n399), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n377), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT91), .ZN(G369));
  NAND3_X1  g0474(.A1(new_n276), .A2(new_n232), .A3(G13), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(KEYINPUT27), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n537), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n680), .B1(new_n545), .B2(new_n547), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n546), .A2(new_n535), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(new_n680), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G330), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n516), .B1(new_n507), .B2(new_n679), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(new_n653), .B2(new_n679), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n682), .A2(new_n679), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT92), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g0492(.A(new_n679), .B(KEYINPUT93), .Z(new_n693));
  NAND2_X1  g0493(.A1(new_n508), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n689), .A2(new_n692), .A3(new_n694), .ZN(G399));
  NOR2_X1   g0495(.A1(new_n225), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n229), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n663), .A2(KEYINPUT94), .A3(new_n659), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n599), .A2(new_n592), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(KEYINPUT26), .A3(new_n658), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(KEYINPUT94), .B1(new_n663), .B2(new_n659), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n600), .A2(new_n648), .A3(new_n654), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(new_n661), .ZN(new_n709));
  OAI211_X1 g0509(.A(KEYINPUT29), .B(new_n679), .C1(new_n707), .C2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n693), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(new_n655), .B2(new_n664), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n710), .B1(KEYINPUT29), .B2(new_n712), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n508), .A2(new_n515), .A3(new_n711), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n548), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n633), .A2(new_n628), .A3(new_n634), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT87), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n715), .B1(new_n718), .B2(new_n635), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n481), .A2(new_n621), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n526), .A2(new_n531), .A3(G179), .A4(new_n480), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n720), .A2(new_n722), .A3(new_n579), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(KEYINPUT30), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT30), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n721), .A2(new_n481), .A3(new_n621), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(new_n579), .ZN(new_n727));
  AOI21_X1  g0527(.A(G179), .B1(new_n643), .B2(new_n620), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n728), .A2(new_n481), .A3(new_n532), .ZN(new_n729));
  OAI22_X1  g0529(.A1(new_n724), .A2(new_n727), .B1(new_n598), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n711), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT31), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n729), .A2(new_n598), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n723), .A2(KEYINPUT30), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n726), .A2(new_n725), .A3(new_n579), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n733), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n732), .B1(new_n736), .B2(new_n679), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n731), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(G330), .B1(new_n719), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n713), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n701), .B1(new_n741), .B2(G1), .ZN(G364));
  NAND2_X1  g0542(.A1(new_n232), .A2(G13), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT95), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G45), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G1), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n696), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n686), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n684), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n748), .B1(G330), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n225), .A2(new_n292), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G355), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(G116), .B2(new_n224), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n225), .A2(new_n266), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n755), .B1(new_n465), .B2(new_n230), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n255), .A2(G45), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G13), .A2(G33), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(G20), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n231), .B1(G20), .B2(new_n359), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n747), .B1(new_n758), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n257), .A2(G190), .ZN(new_n766));
  OAI21_X1  g0566(.A(G20), .B1(new_n766), .B2(G179), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT96), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G97), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n232), .A2(new_n338), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(G190), .A3(G200), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n232), .A2(G179), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n776), .A2(new_n285), .A3(G200), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n775), .A2(new_n202), .B1(new_n777), .B2(new_n436), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n774), .A2(new_n285), .A3(G200), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n776), .A2(G190), .A3(G200), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n779), .A2(new_n298), .B1(new_n780), .B2(new_n212), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G190), .A2(G200), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n776), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G159), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT32), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n766), .A2(new_n232), .A3(new_n338), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n266), .B1(new_n789), .B2(new_n297), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n774), .A2(new_n783), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n790), .B1(G77), .B2(new_n792), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n773), .A2(new_n782), .A3(new_n787), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n792), .A2(G311), .ZN(new_n795));
  INV_X1    g0595(.A(new_n775), .ZN(new_n796));
  INV_X1    g0596(.A(new_n780), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G326), .A2(new_n796), .B1(new_n797), .B2(G303), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n266), .B1(new_n788), .B2(G322), .ZN(new_n799));
  INV_X1    g0599(.A(new_n779), .ZN(new_n800));
  INV_X1    g0600(.A(G317), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(KEYINPUT33), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n801), .A2(KEYINPUT33), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n800), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  AND4_X1   g0604(.A1(new_n795), .A2(new_n798), .A3(new_n799), .A4(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G294), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n805), .B1(new_n806), .B2(new_n771), .ZN(new_n807));
  INV_X1    g0607(.A(G283), .ZN(new_n808));
  INV_X1    g0608(.A(G329), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n777), .A2(new_n808), .B1(new_n784), .B2(new_n809), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT97), .Z(new_n811));
  OAI21_X1  g0611(.A(new_n794), .B1(new_n807), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n765), .B1(new_n812), .B2(new_n762), .ZN(new_n813));
  INV_X1    g0613(.A(new_n761), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n749), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n750), .A2(new_n815), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT98), .Z(G396));
  INV_X1    g0617(.A(new_n679), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n456), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n450), .A2(new_n818), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n453), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n819), .B1(new_n821), .B2(new_n456), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n712), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n665), .A2(new_n693), .A3(new_n822), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n747), .B1(new_n825), .B2(new_n739), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n739), .B2(new_n825), .ZN(new_n827));
  INV_X1    g0627(.A(new_n747), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n762), .A2(new_n759), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n828), .B1(new_n352), .B2(new_n829), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n775), .A2(new_n529), .B1(new_n780), .B2(new_n436), .ZN(new_n831));
  INV_X1    g0631(.A(G311), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n292), .B1(new_n784), .B2(new_n832), .C1(new_n789), .C2(new_n806), .ZN(new_n833));
  INV_X1    g0633(.A(new_n777), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n831), .B(new_n833), .C1(G87), .C2(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n800), .A2(G283), .B1(new_n792), .B2(G116), .ZN(new_n836));
  OR2_X1    g0636(.A1(new_n836), .A2(KEYINPUT99), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(KEYINPUT99), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n835), .A2(new_n773), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n792), .A2(G159), .B1(new_n788), .B2(G143), .ZN(new_n840));
  INV_X1    g0640(.A(G137), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n840), .B1(new_n841), .B2(new_n775), .C1(new_n366), .C2(new_n779), .ZN(new_n842));
  XOR2_X1   g0642(.A(new_n842), .B(KEYINPUT34), .Z(new_n843));
  NAND2_X1  g0643(.A1(new_n834), .A2(G68), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n844), .B1(new_n202), .B2(new_n780), .C1(new_n771), .C2(new_n297), .ZN(new_n845));
  INV_X1    g0645(.A(new_n784), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n292), .B1(new_n846), .B2(G132), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT100), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n839), .B1(new_n843), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n850), .A2(KEYINPUT101), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(KEYINPUT101), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n762), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n830), .B1(new_n822), .B2(new_n760), .C1(new_n851), .C2(new_n853), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n827), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(G384));
  NOR2_X1   g0656(.A1(new_n744), .A2(new_n276), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT40), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT103), .ZN(new_n859));
  AND3_X1   g0659(.A1(new_n317), .A2(new_n859), .A3(new_n323), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n859), .B1(new_n317), .B2(new_n323), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n678), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n340), .B1(new_n860), .B2(new_n861), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n325), .B1(new_n291), .B2(new_n324), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n333), .A2(KEYINPUT79), .A3(new_n334), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n862), .A2(new_n863), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT37), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT37), .B1(new_n340), .B2(new_n324), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n324), .A2(new_n678), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n864), .A2(new_n868), .A3(new_n865), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n862), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n348), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT38), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n871), .A2(new_n873), .A3(KEYINPUT38), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n434), .B1(new_n409), .B2(new_n818), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n409), .A2(new_n818), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(new_n426), .B2(new_n433), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n822), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n715), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n629), .B2(new_n636), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n730), .A2(new_n818), .B1(KEYINPUT105), .B2(new_n732), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n732), .A2(KEYINPUT105), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n736), .A2(new_n679), .A3(new_n886), .ZN(new_n887));
  OR2_X1    g0687(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n884), .A2(KEYINPUT106), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT106), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n885), .A2(new_n887), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n890), .B1(new_n719), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n882), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT107), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n878), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI211_X1 g0695(.A(KEYINPUT107), .B(new_n882), .C1(new_n889), .C2(new_n892), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n858), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT104), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n877), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n871), .A2(new_n873), .A3(KEYINPUT104), .A4(KEYINPUT38), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n870), .A2(new_n875), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n348), .A2(new_n324), .A3(new_n678), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n340), .A2(new_n324), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n345), .A2(new_n904), .A3(new_n869), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n905), .A2(KEYINPUT37), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n902), .B1(new_n903), .B2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n901), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(KEYINPUT40), .A3(new_n893), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n897), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n889), .A2(new_n892), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n463), .A2(new_n912), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n911), .A2(new_n913), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n914), .A2(new_n915), .A3(new_n685), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n672), .B1(new_n464), .B2(new_n713), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n344), .A2(new_n678), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n434), .B(new_n880), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n819), .B(KEYINPUT102), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n920), .B1(new_n824), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n919), .B1(new_n922), .B2(new_n878), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n426), .A2(new_n818), .ZN(new_n924));
  INV_X1    g0724(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n876), .A2(KEYINPUT39), .A3(new_n877), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n907), .B1(new_n899), .B2(new_n900), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n925), .B(new_n926), .C1(new_n927), .C2(KEYINPUT39), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n923), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n918), .B(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n857), .B1(new_n917), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n930), .B2(new_n917), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n587), .A2(KEYINPUT35), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n587), .A2(KEYINPUT35), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n933), .A2(new_n934), .A3(G116), .A4(new_n233), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT36), .ZN(new_n936));
  NOR3_X1   g0736(.A1(new_n229), .A2(new_n352), .A3(new_n299), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n298), .A2(G50), .ZN(new_n938));
  OAI211_X1 g0738(.A(G1), .B(new_n318), .C1(new_n937), .C2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n932), .A2(new_n936), .A3(new_n939), .ZN(G367));
  NAND2_X1  g0740(.A1(new_n610), .A2(new_n818), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n658), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n661), .B2(new_n941), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n600), .B1(new_n564), .B2(new_n693), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n703), .A2(new_n711), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n947), .A2(new_n688), .A3(new_n691), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(KEYINPUT42), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n947), .A2(new_n508), .B1(new_n599), .B2(new_n596), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n949), .B1(new_n711), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n948), .A2(KEYINPUT42), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n944), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n943), .A2(KEYINPUT43), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n953), .B(new_n954), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n945), .A2(new_n946), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n689), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n955), .B(new_n957), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n696), .B(KEYINPUT41), .Z(new_n959));
  INV_X1    g0759(.A(KEYINPUT108), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n692), .A2(new_n694), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n960), .B1(new_n961), .B2(new_n956), .ZN(new_n962));
  AOI211_X1 g0762(.A(KEYINPUT108), .B(new_n947), .C1(new_n692), .C2(new_n694), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT44), .ZN(new_n964));
  OR3_X1    g0764(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n961), .A2(new_n956), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT45), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n964), .B1(new_n962), .B2(new_n963), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n965), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n689), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n686), .A2(new_n688), .ZN(new_n972));
  AND3_X1   g0772(.A1(new_n972), .A2(new_n689), .A3(new_n691), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n691), .B1(new_n972), .B2(new_n689), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n741), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n965), .A2(new_n967), .A3(new_n689), .A4(new_n968), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n971), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n959), .B1(new_n979), .B2(new_n741), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n958), .B1(new_n980), .B2(new_n746), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n247), .A2(new_n755), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n763), .B1(new_n224), .B2(new_n446), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n747), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n791), .A2(new_n808), .B1(new_n784), .B2(new_n801), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n292), .B1(new_n789), .B2(new_n529), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n780), .A2(new_n518), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n985), .B(new_n986), .C1(KEYINPUT46), .C2(new_n987), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(KEYINPUT46), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n772), .A2(G107), .ZN(new_n990));
  OAI22_X1  g0790(.A1(new_n779), .A2(new_n806), .B1(new_n777), .B2(new_n214), .ZN(new_n991));
  XOR2_X1   g0791(.A(KEYINPUT109), .B(G311), .Z(new_n992));
  AOI21_X1  g0792(.A(new_n991), .B1(new_n796), .B2(new_n992), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n988), .A2(new_n989), .A3(new_n990), .A4(new_n993), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n779), .A2(new_n785), .B1(new_n780), .B2(new_n297), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(G143), .B2(new_n796), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n846), .A2(G137), .B1(new_n788), .B2(G150), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n996), .B(new_n997), .C1(new_n202), .C2(new_n791), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n772), .A2(G68), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT110), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n777), .A2(new_n352), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1000), .B1(new_n1001), .B2(new_n292), .ZN(new_n1002));
  OAI211_X1 g0802(.A(KEYINPUT110), .B(new_n266), .C1(new_n777), .C2(new_n352), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n999), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n994), .B1(new_n998), .B2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT47), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n984), .B1(new_n1006), .B2(new_n762), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n814), .B2(new_n943), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n981), .A2(new_n1008), .ZN(G387));
  NOR2_X1   g0809(.A1(new_n977), .A2(new_n697), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n741), .B2(new_n975), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n975), .A2(new_n746), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n762), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n266), .B1(new_n846), .B2(G326), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n518), .B2(new_n777), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n792), .A2(G303), .B1(new_n788), .B2(G317), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT112), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G322), .A2(new_n796), .B1(new_n800), .B2(new_n992), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT113), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n1020), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1021), .A2(KEYINPUT48), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(KEYINPUT48), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n771), .A2(new_n808), .B1(new_n806), .B2(new_n780), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1015), .B1(new_n1025), .B2(KEYINPUT49), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(KEYINPUT49), .B2(new_n1025), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n292), .B1(new_n846), .B2(G150), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n352), .B2(new_n780), .C1(new_n214), .C2(new_n777), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT111), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n772), .A2(new_n623), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n792), .A2(G68), .B1(new_n788), .B2(G50), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n321), .B2(new_n779), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G159), .B2(new_n796), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1030), .A2(new_n1031), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1013), .B1(new_n1027), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n698), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1037), .A2(new_n751), .B1(new_n436), .B2(new_n225), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n243), .A2(new_n465), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n321), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n202), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1041), .B(KEYINPUT50), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n698), .B(new_n465), .C1(new_n298), .C2(new_n352), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n754), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1038), .B1(new_n1039), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n828), .B1(new_n1045), .B2(new_n763), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n688), .B2(new_n814), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1012), .B1(new_n1036), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1011), .A2(new_n1049), .ZN(G393));
  NAND2_X1  g0850(.A1(new_n971), .A2(new_n978), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n746), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n956), .A2(new_n761), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n252), .A2(new_n754), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n763), .B1(new_n214), .B2(new_n224), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n747), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n772), .A2(G77), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n792), .A2(new_n1040), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n292), .B1(new_n846), .B2(G143), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n298), .A2(new_n780), .B1(new_n777), .B2(new_n212), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(G50), .B2(new_n800), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .A4(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n796), .A2(G150), .B1(G159), .B2(new_n788), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT51), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n791), .A2(new_n806), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n266), .B(new_n1066), .C1(G322), .C2(new_n846), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n436), .A2(new_n777), .B1(new_n780), .B2(new_n808), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(G303), .B2(new_n800), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1067), .B(new_n1069), .C1(new_n518), .C2(new_n771), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n796), .A2(G317), .B1(G311), .B2(new_n788), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT52), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n1063), .A2(new_n1065), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1057), .B1(new_n762), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1053), .B1(new_n1054), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1051), .A2(new_n976), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1076), .A2(new_n696), .A3(new_n979), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1077), .ZN(G390));
  NAND2_X1  g0878(.A1(new_n821), .A2(new_n456), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n679), .B(new_n1079), .C1(new_n707), .C2(new_n709), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n819), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n920), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1084), .A2(new_n909), .A3(new_n924), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n926), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT39), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1086), .B1(new_n909), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n922), .A2(new_n925), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1085), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n685), .B1(new_n889), .B2(new_n892), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n882), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g0895(.A(G330), .B(new_n822), .C1(new_n719), .C2(new_n738), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1096), .A2(new_n920), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1085), .B(new_n1098), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1095), .A2(new_n746), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n828), .B1(new_n321), .B2(new_n829), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT115), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n788), .A2(G132), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(KEYINPUT54), .B(G143), .ZN(new_n1104));
  INV_X1    g0904(.A(G128), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1103), .B1(new_n791), .B2(new_n1104), .C1(new_n1105), .C2(new_n775), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n797), .A2(G150), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT53), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1106), .B(new_n1108), .C1(G137), .C2(new_n800), .ZN(new_n1109));
  INV_X1    g0909(.A(G125), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n266), .B1(new_n784), .B2(new_n1110), .C1(new_n202), .C2(new_n777), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT116), .Z(new_n1112));
  OAI211_X1 g0912(.A(new_n1109), .B(new_n1112), .C1(new_n785), .C2(new_n771), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1113), .A2(KEYINPUT117), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1113), .A2(KEYINPUT117), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n789), .A2(new_n518), .B1(new_n791), .B2(new_n214), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n844), .B1(new_n436), .B2(new_n779), .C1(new_n808), .C2(new_n775), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n1116), .B(new_n1117), .C1(G294), .C2(new_n846), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n292), .B1(new_n780), .B2(new_n212), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT118), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1118), .A2(new_n1058), .A3(new_n1120), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1114), .A2(new_n1115), .A3(new_n1121), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1102), .B1(new_n1122), .B2(new_n1013), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n926), .B1(new_n927), .B2(KEYINPUT39), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1123), .B1(new_n1124), .B2(new_n759), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT119), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1100), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1096), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1093), .B1(new_n1083), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n824), .A2(new_n921), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1083), .B1(new_n1091), .B2(new_n822), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n1080), .B(new_n1081), .C1(new_n1096), .C2(new_n920), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n1132), .A2(new_n1133), .A3(KEYINPUT114), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT114), .ZN(new_n1135));
  AOI21_X1  g0935(.A(KEYINPUT106), .B1(new_n884), .B2(new_n888), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n719), .A2(new_n890), .A3(new_n891), .ZN(new_n1137));
  OAI211_X1 g0937(.A(G330), .B(new_n822), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n920), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1133), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1135), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1131), .B1(new_n1134), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n463), .A2(new_n1091), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1143), .B(new_n672), .C1(new_n464), .C2(new_n713), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  OR2_X1    g0946(.A1(new_n922), .A2(new_n925), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n927), .A2(new_n925), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n1147), .A2(new_n1124), .B1(new_n1084), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1099), .B1(new_n1149), .B2(new_n1093), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n697), .B1(new_n1146), .B2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1142), .A2(new_n1099), .A3(new_n1095), .A4(new_n1145), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1127), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(G378));
  OAI22_X1  g0954(.A1(new_n775), .A2(new_n1110), .B1(new_n780), .B2(new_n1104), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n800), .A2(G132), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1156), .B1(new_n1105), .B2(new_n789), .C1(new_n841), .C2(new_n791), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1155), .B(new_n1157), .C1(G150), .C2(new_n772), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT59), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1161));
  AOI211_X1 g0961(.A(G33), .B(G41), .C1(new_n846), .C2(G124), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n785), .B2(new_n777), .ZN(new_n1163));
  NOR3_X1   g0963(.A1(new_n1160), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n777), .A2(new_n297), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n214), .A2(new_n779), .B1(new_n775), .B2(new_n518), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1165), .B(new_n1166), .C1(G77), .C2(new_n797), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n266), .A2(G41), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1168), .B1(new_n808), .B2(new_n784), .C1(new_n789), .C2(new_n436), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n623), .B2(new_n792), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1167), .A2(new_n1170), .A3(new_n999), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT58), .ZN(new_n1172));
  OR2_X1    g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1174));
  AOI211_X1 g0974(.A(G50), .B(new_n1168), .C1(new_n258), .C2(new_n259), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT120), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1173), .A2(new_n1174), .A3(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n762), .B1(new_n1164), .B2(new_n1177), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT121), .Z(new_n1179));
  AOI211_X1 g0979(.A(new_n828), .B(new_n1179), .C1(new_n202), .C2(new_n829), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n375), .A2(new_n678), .ZN(new_n1181));
  XOR2_X1   g0981(.A(new_n400), .B(new_n1181), .Z(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1182), .B(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1180), .B1(new_n1184), .B2(new_n760), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT122), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n927), .A2(new_n858), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n685), .B1(new_n1187), .B2(new_n893), .ZN(new_n1188));
  AND3_X1   g0988(.A1(new_n897), .A2(new_n929), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n929), .B1(new_n897), .B2(new_n1188), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1184), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  AND2_X1   g0991(.A1(new_n923), .A2(new_n928), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n878), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1092), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1193), .B1(new_n1194), .B2(KEYINPUT107), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n893), .A2(new_n894), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT40), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n910), .A2(G330), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1192), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1184), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n897), .A2(new_n929), .A3(new_n1188), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1191), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1186), .B1(new_n746), .B2(new_n1203), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1202), .A2(new_n1191), .B1(new_n1152), .B2(new_n1145), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n696), .B1(new_n1205), .B2(KEYINPUT57), .ZN(new_n1206));
  OAI21_X1  g1006(.A(KEYINPUT114), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1139), .A2(new_n1135), .A3(new_n1140), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1207), .A2(new_n1208), .B1(new_n1130), .B2(new_n1129), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1145), .B1(new_n1150), .B2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1203), .A2(KEYINPUT57), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1204), .B1(new_n1206), .B2(new_n1212), .ZN(G375));
  NAND2_X1  g1013(.A1(new_n920), .A2(new_n759), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n779), .A2(new_n1104), .B1(new_n780), .B2(new_n785), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n1165), .B(new_n1215), .C1(G132), .C2(new_n796), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n791), .A2(new_n366), .B1(new_n784), .B2(new_n1105), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n292), .B(new_n1217), .C1(G137), .C2(new_n788), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1216), .B(new_n1218), .C1(new_n202), .C2(new_n771), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n775), .A2(new_n806), .B1(new_n780), .B2(new_n214), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1001), .B(new_n1220), .C1(G116), .C2(new_n800), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n266), .B1(new_n846), .B2(G303), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n792), .A2(G107), .B1(new_n788), .B2(G283), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1221), .A2(new_n1031), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1013), .B1(new_n1219), .B2(new_n1224), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n828), .B(new_n1225), .C1(new_n298), .C2(new_n829), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n1142), .A2(new_n746), .B1(new_n1214), .B2(new_n1226), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1209), .A2(new_n1144), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1228), .A2(new_n959), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1144), .B(new_n1131), .C1(new_n1134), .C2(new_n1141), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1227), .B1(new_n1229), .B2(new_n1231), .ZN(G381));
  INV_X1    g1032(.A(G390), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(G393), .A2(G396), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1233), .A2(new_n855), .A3(new_n1234), .ZN(new_n1235));
  OR3_X1    g1035(.A1(new_n1235), .A2(G387), .A3(G381), .ZN(new_n1236));
  OR3_X1    g1036(.A1(new_n1236), .A2(G378), .A3(G375), .ZN(G407));
  INV_X1    g1037(.A(G343), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(G213), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1153), .A2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(G407), .B(G213), .C1(G375), .C2(new_n1241), .ZN(G409));
  NAND2_X1  g1042(.A1(new_n1233), .A2(G387), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(G390), .A2(new_n981), .A3(new_n1008), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  AND2_X1   g1045(.A1(G393), .A2(G396), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1245), .B1(new_n1234), .B2(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1234), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1243), .A2(new_n1248), .A3(new_n1244), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1250));
  OAI211_X1 g1050(.A(G378), .B(new_n1204), .C1(new_n1206), .C2(new_n1212), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT123), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1191), .A2(new_n1252), .A3(new_n1202), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1252), .B1(new_n1191), .B2(new_n1202), .ZN(new_n1254));
  NOR3_X1   g1054(.A1(new_n1253), .A2(new_n1254), .A3(new_n1052), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1186), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1200), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1210), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1256), .B1(new_n1259), .B2(new_n959), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1153), .B1(new_n1255), .B2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1251), .A2(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1228), .A2(new_n697), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT124), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT60), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1264), .B(new_n1265), .C1(new_n1209), .C2(new_n1144), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT60), .B1(new_n1230), .B2(KEYINPUT124), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1263), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1268), .A2(G384), .A3(new_n1227), .ZN(new_n1269));
  AOI21_X1  g1069(.A(G384), .B1(new_n1268), .B2(new_n1227), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1262), .A2(new_n1239), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT62), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1240), .B1(new_n1251), .B2(new_n1261), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1275), .A2(KEYINPUT62), .A3(new_n1271), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1274), .A2(KEYINPUT125), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1262), .A2(new_n1239), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1240), .A2(G2897), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1146), .A2(new_n696), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1230), .A2(KEYINPUT124), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1265), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1230), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1282), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1227), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n855), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1268), .A2(G384), .A3(new_n1227), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1288), .A2(new_n1289), .A3(new_n1279), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1281), .A2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT61), .B1(new_n1278), .B2(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1292), .B1(new_n1274), .B2(KEYINPUT125), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1250), .B1(new_n1277), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT126), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT61), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1281), .A2(new_n1290), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT63), .ZN(new_n1298));
  OAI221_X1 g1098(.A(new_n1296), .B1(new_n1275), .B2(new_n1297), .C1(new_n1272), .C2(new_n1298), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1272), .A2(new_n1298), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  OR2_X1    g1102(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1294), .A2(new_n1295), .A3(new_n1303), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1296), .B1(new_n1275), .B2(new_n1297), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT125), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT62), .B1(new_n1275), .B2(new_n1271), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1305), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1274), .A2(KEYINPUT125), .A3(new_n1276), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1300), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1311));
  OAI21_X1  g1111(.A(KEYINPUT126), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1304), .A2(new_n1312), .ZN(G405));
  NAND2_X1  g1113(.A1(G375), .A2(new_n1153), .ZN(new_n1314));
  AND2_X1   g1114(.A1(new_n1314), .A2(new_n1251), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1300), .A2(new_n1271), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT127), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1250), .B1(new_n1270), .B2(new_n1269), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1317), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1318), .B1(new_n1317), .B2(new_n1319), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1316), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1317), .A2(new_n1319), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(KEYINPUT127), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1317), .A2(new_n1318), .A3(new_n1319), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1324), .A2(new_n1315), .A3(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1322), .A2(new_n1326), .ZN(G402));
endmodule


