//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 0 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n187));
  XNOR2_X1  g001(.A(G110), .B(G140), .ZN(new_n188));
  OR2_X1    g002(.A1(new_n188), .A2(KEYINPUT77), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT78), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(KEYINPUT77), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(new_n190), .A3(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G227), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G953), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n188), .A2(KEYINPUT77), .ZN(new_n195));
  INV_X1    g009(.A(G140), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G110), .ZN(new_n197));
  INV_X1    g011(.A(G110), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G140), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n197), .A2(new_n199), .A3(KEYINPUT77), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT78), .B1(new_n195), .B2(new_n200), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n192), .A2(new_n194), .A3(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n194), .B1(new_n192), .B2(new_n201), .ZN(new_n203));
  OR2_X1    g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT11), .ZN(new_n205));
  INV_X1    g019(.A(G134), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(G137), .ZN(new_n207));
  INV_X1    g021(.A(G137), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT11), .A3(G134), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(G137), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G131), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n207), .A2(new_n209), .A3(new_n213), .A4(new_n210), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G104), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT3), .B1(new_n217), .B2(G107), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n219));
  INV_X1    g033(.A(G107), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G104), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n217), .A2(G107), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n218), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n223), .A2(new_n224), .A3(G101), .ZN(new_n225));
  INV_X1    g039(.A(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G143), .ZN(new_n227));
  INV_X1    g041(.A(G143), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G146), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n227), .A2(new_n229), .A3(KEYINPUT0), .A4(G128), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n228), .A2(G146), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n226), .A2(G143), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT0), .B(G128), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n230), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n225), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n223), .A2(G101), .ZN(new_n237));
  INV_X1    g051(.A(G101), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n218), .A2(new_n221), .A3(new_n238), .A4(new_n222), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n237), .A2(KEYINPUT4), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n236), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT10), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT79), .ZN(new_n243));
  XNOR2_X1  g057(.A(G104), .B(G107), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n243), .B1(new_n244), .B2(new_n238), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n217), .A2(G107), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n220), .A2(G104), .ZN(new_n247));
  OAI211_X1 g061(.A(KEYINPUT79), .B(G101), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n245), .A2(new_n239), .A3(new_n248), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT1), .B1(new_n228), .B2(G146), .ZN(new_n250));
  OAI211_X1 g064(.A(G128), .B(new_n250), .C1(new_n231), .C2(new_n232), .ZN(new_n251));
  INV_X1    g065(.A(G128), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n227), .B(new_n229), .C1(KEYINPUT1), .C2(new_n252), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n242), .B1(new_n249), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n245), .A2(new_n239), .A3(new_n248), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n251), .A2(new_n253), .ZN(new_n257));
  NOR3_X1   g071(.A1(new_n256), .A2(KEYINPUT10), .A3(new_n257), .ZN(new_n258));
  OAI211_X1 g072(.A(new_n216), .B(new_n241), .C1(new_n255), .C2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n204), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT80), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n241), .B1(new_n255), .B2(new_n258), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n215), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n204), .A2(new_n259), .A3(KEYINPUT80), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n249), .A2(new_n254), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n256), .A2(new_n257), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT12), .B1(new_n269), .B2(new_n215), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT12), .ZN(new_n271));
  AOI211_X1 g085(.A(new_n271), .B(new_n216), .C1(new_n267), .C2(new_n268), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n259), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n202), .A2(new_n203), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI21_X1  g089(.A(G902), .B1(new_n266), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G469), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n187), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n249), .A2(new_n242), .A3(new_n254), .ZN(new_n279));
  OAI21_X1  g093(.A(KEYINPUT10), .B1(new_n256), .B2(new_n257), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n279), .A2(new_n280), .B1(new_n236), .B2(new_n240), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n274), .B1(new_n281), .B2(new_n216), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n282), .A2(KEYINPUT80), .B1(new_n215), .B2(new_n263), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n283), .A2(new_n262), .B1(new_n273), .B2(new_n274), .ZN(new_n284));
  OAI211_X1 g098(.A(KEYINPUT81), .B(G469), .C1(new_n284), .C2(G902), .ZN(new_n285));
  INV_X1    g099(.A(G902), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n259), .B(new_n204), .C1(new_n270), .C2(new_n272), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n204), .B1(new_n264), .B2(new_n259), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT82), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n287), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI211_X1 g104(.A(KEYINPUT82), .B(new_n204), .C1(new_n264), .C2(new_n259), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n277), .B(new_n286), .C1(new_n290), .C2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n278), .A2(new_n285), .A3(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(G214), .B1(G237), .B2(G902), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n223), .A2(new_n224), .A3(G101), .ZN(new_n296));
  XNOR2_X1  g110(.A(KEYINPUT2), .B(G113), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT64), .ZN(new_n299));
  INV_X1    g113(.A(G119), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n299), .B1(new_n300), .B2(G116), .ZN(new_n301));
  INV_X1    g115(.A(G116), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(KEYINPUT64), .A3(G119), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n300), .A2(G116), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n298), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n298), .B1(new_n305), .B2(new_n304), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n296), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n240), .ZN(new_n310));
  OAI21_X1  g124(.A(G113), .B1(new_n305), .B2(KEYINPUT5), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n304), .A2(new_n305), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT5), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n306), .A2(new_n239), .A3(new_n248), .A4(new_n245), .ZN(new_n317));
  OAI22_X1  g131(.A1(new_n309), .A2(new_n310), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G110), .B(G122), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n319), .B(KEYINPUT83), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  OAI221_X1 g136(.A(new_n320), .B1(new_n316), .B2(new_n317), .C1(new_n309), .C2(new_n310), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n323), .A3(KEYINPUT6), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT6), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n318), .A2(new_n325), .A3(new_n321), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT72), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(KEYINPUT72), .A2(G125), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n230), .B(new_n331), .C1(new_n233), .C2(new_n234), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n332), .B1(new_n257), .B2(new_n331), .ZN(new_n333));
  INV_X1    g147(.A(G224), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(G953), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n335), .B(KEYINPUT84), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n333), .B(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n324), .A2(new_n326), .A3(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT7), .B1(new_n334), .B2(G953), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n333), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n332), .B(new_n339), .C1(new_n257), .C2(new_n331), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n313), .A2(new_n297), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n225), .B1(new_n344), .B2(new_n306), .ZN(new_n345));
  INV_X1    g159(.A(new_n317), .ZN(new_n346));
  AOI22_X1  g160(.A1(new_n240), .A2(new_n345), .B1(new_n346), .B2(new_n315), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n343), .B1(new_n347), .B2(new_n320), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n320), .B(KEYINPUT8), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n311), .B(KEYINPUT85), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n313), .A2(new_n314), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n352), .A2(new_n317), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n249), .B1(new_n306), .B2(new_n315), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n349), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(G902), .B1(new_n348), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(G210), .B1(G237), .B2(G902), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n338), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n357), .B1(new_n338), .B2(new_n356), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n295), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(KEYINPUT9), .B(G234), .ZN(new_n363));
  OAI21_X1  g177(.A(G221), .B1(new_n363), .B2(G902), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n293), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT68), .ZN(new_n366));
  NOR2_X1   g180(.A1(G472), .A2(G902), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT31), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n307), .A2(new_n308), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n206), .A2(G137), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n208), .A2(G134), .ZN(new_n372));
  OAI21_X1  g186(.A(G131), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n214), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT65), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n254), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n235), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n215), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n251), .A2(new_n214), .A3(new_n373), .A4(new_n253), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT65), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n376), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT30), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT30), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n378), .A2(new_n383), .A3(new_n379), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n370), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n376), .A2(new_n370), .A3(new_n378), .A4(new_n380), .ZN(new_n386));
  XOR2_X1   g200(.A(KEYINPUT66), .B(KEYINPUT27), .Z(new_n387));
  NOR2_X1   g201(.A1(G237), .A2(G953), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G210), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n387), .B(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT26), .B(G101), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n390), .B(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n369), .B1(new_n385), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n393), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n378), .A2(new_n383), .A3(new_n379), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n396), .B1(KEYINPUT30), .B2(new_n381), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n395), .B(KEYINPUT31), .C1(new_n397), .C2(new_n370), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n370), .A2(new_n378), .A3(new_n379), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT28), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n378), .A2(new_n379), .ZN(new_n403));
  INV_X1    g217(.A(new_n370), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n402), .B(new_n405), .C1(new_n401), .C2(new_n386), .ZN(new_n406));
  INV_X1    g220(.A(new_n392), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n368), .B1(new_n399), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT67), .B(KEYINPUT32), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n366), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n410), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n394), .A2(new_n398), .B1(new_n407), .B2(new_n406), .ZN(new_n413));
  OAI211_X1 g227(.A(KEYINPUT68), .B(new_n412), .C1(new_n413), .C2(new_n368), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n381), .B(new_n370), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n402), .B1(new_n416), .B2(new_n401), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n392), .A2(KEYINPUT29), .ZN(new_n418));
  INV_X1    g232(.A(new_n386), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n385), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n420), .A2(new_n392), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT29), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n406), .B2(new_n407), .ZN(new_n423));
  OAI221_X1 g237(.A(new_n286), .B1(new_n417), .B2(new_n418), .C1(new_n421), .C2(new_n423), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n424), .A2(G472), .B1(new_n409), .B2(KEYINPUT32), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n415), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT25), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT22), .B(G137), .ZN(new_n428));
  INV_X1    g242(.A(G953), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n429), .A2(G221), .A3(G234), .ZN(new_n430));
  XOR2_X1   g244(.A(new_n428), .B(new_n430), .Z(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT73), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT24), .B(G110), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT70), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n300), .A2(G128), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n252), .A2(G119), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n252), .A2(G119), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n300), .A2(G128), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT70), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n435), .B1(new_n439), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT23), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(new_n300), .B2(G128), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n252), .A2(KEYINPUT23), .A3(G119), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n445), .A2(new_n446), .A3(new_n198), .A4(new_n441), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n433), .B1(new_n443), .B2(new_n448), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT70), .ZN(new_n450));
  AOI21_X1  g264(.A(KEYINPUT70), .B1(new_n440), .B2(new_n441), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n434), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n447), .A3(KEYINPUT73), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n329), .A2(G140), .A3(new_n330), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT71), .B1(new_n328), .B2(G140), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT71), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(new_n196), .A3(G125), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n454), .A2(KEYINPUT16), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT16), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n331), .A2(new_n459), .A3(new_n196), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(G146), .A3(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(G125), .B(G140), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n226), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n449), .A2(new_n453), .A3(new_n461), .A4(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT74), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n450), .A2(new_n451), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n445), .A2(new_n441), .A3(new_n446), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n466), .A2(new_n435), .B1(G110), .B2(new_n467), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n458), .A2(G146), .A3(new_n460), .ZN(new_n469));
  AOI21_X1  g283(.A(G146), .B1(new_n458), .B2(new_n460), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AND3_X1   g285(.A1(new_n464), .A2(new_n465), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n465), .B1(new_n464), .B2(new_n471), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n432), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n464), .A2(new_n471), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n431), .ZN(new_n476));
  AOI21_X1  g290(.A(G902), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  OAI211_X1 g291(.A(KEYINPUT76), .B(new_n427), .C1(new_n477), .C2(KEYINPUT75), .ZN(new_n478));
  NAND2_X1  g292(.A1(G217), .A2(G902), .ZN(new_n479));
  INV_X1    g293(.A(G217), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n479), .B1(new_n480), .B2(G234), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT69), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT76), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n475), .A2(KEYINPUT74), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n464), .A2(new_n465), .A3(new_n471), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n431), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n476), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n286), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT75), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n483), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT25), .B1(new_n477), .B2(KEYINPUT76), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n478), .B(new_n482), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n474), .A2(new_n476), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n482), .A2(G902), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n492), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(G475), .A2(G902), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(G113), .B(G122), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(new_n217), .ZN(new_n500));
  AND2_X1   g314(.A1(KEYINPUT72), .A2(G125), .ZN(new_n501));
  NOR2_X1   g315(.A1(KEYINPUT72), .A2(G125), .ZN(new_n502));
  NOR3_X1   g316(.A1(new_n501), .A2(new_n502), .A3(new_n196), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n455), .A2(new_n457), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT86), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT86), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n454), .A2(new_n506), .A3(new_n455), .A4(new_n457), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n505), .A2(KEYINPUT19), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT19), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n462), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n226), .A3(new_n510), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n388), .A2(G143), .A3(G214), .ZN(new_n512));
  AOI21_X1  g326(.A(G143), .B1(new_n388), .B2(G214), .ZN(new_n513));
  OAI21_X1  g327(.A(G131), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(G237), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(new_n429), .A3(G214), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n228), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n388), .A2(G143), .A3(G214), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(new_n213), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n461), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n511), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n505), .A2(G146), .A3(new_n507), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n463), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n517), .A2(new_n518), .ZN(new_n525));
  NAND2_X1  g339(.A1(KEYINPUT18), .A2(G131), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n525), .B(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n500), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n469), .A2(new_n470), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n514), .A2(new_n531), .A3(new_n519), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n525), .A2(KEYINPUT17), .A3(G131), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n530), .A2(new_n534), .B1(new_n524), .B2(new_n527), .ZN(new_n535));
  AOI22_X1  g349(.A1(new_n529), .A2(KEYINPUT87), .B1(new_n500), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT87), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n511), .A2(new_n521), .B1(new_n524), .B2(new_n527), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n537), .B1(new_n538), .B2(new_n500), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n498), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT20), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT88), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n522), .A2(new_n528), .ZN(new_n543));
  INV_X1    g357(.A(new_n500), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(KEYINPUT87), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n535), .A2(new_n500), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n539), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(new_n497), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT88), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT20), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n547), .A2(new_n541), .A3(new_n497), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT89), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT89), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n540), .A2(new_n553), .A3(new_n541), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n542), .A2(new_n550), .A3(new_n552), .A4(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G475), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n535), .B(new_n500), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n556), .B1(new_n557), .B2(new_n286), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n228), .A2(G128), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n252), .A2(G143), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(new_n206), .ZN(new_n563));
  XNOR2_X1  g377(.A(G116), .B(G122), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n220), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n302), .A2(KEYINPUT14), .A3(G122), .ZN(new_n566));
  INV_X1    g380(.A(new_n564), .ZN(new_n567));
  OAI211_X1 g381(.A(G107), .B(new_n566), .C1(new_n567), .C2(KEYINPUT14), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n563), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n560), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n570), .A2(KEYINPUT13), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n561), .B1(new_n570), .B2(KEYINPUT13), .ZN(new_n572));
  OAI21_X1  g386(.A(G134), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n562), .A2(new_n206), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n564), .B(new_n220), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n569), .A2(new_n576), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n363), .A2(new_n480), .A3(G953), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(KEYINPUT90), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n579), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(new_n576), .A3(new_n569), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT91), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n581), .A2(KEYINPUT91), .A3(new_n576), .A4(new_n569), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n585), .A3(new_n286), .ZN(new_n586));
  INV_X1    g400(.A(G478), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(KEYINPUT15), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n588), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n584), .A2(new_n585), .A3(new_n286), .A4(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(G952), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(G953), .ZN(new_n593));
  NAND2_X1  g407(.A1(G234), .A2(G237), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(G898), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n429), .B1(KEYINPUT21), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n597), .B1(KEYINPUT21), .B2(new_n596), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n594), .A2(G902), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n595), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n589), .A2(new_n591), .A3(new_n600), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n555), .A2(new_n559), .A3(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n365), .A2(new_n426), .A3(new_n496), .A4(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n584), .A2(new_n585), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n580), .A2(new_n582), .A3(KEYINPUT33), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n587), .A2(G902), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n609), .A2(new_n610), .B1(new_n587), .B2(new_n586), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n555), .B2(new_n559), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT92), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n293), .A2(new_n364), .ZN(new_n615));
  INV_X1    g429(.A(new_n409), .ZN(new_n616));
  OAI21_X1  g430(.A(G472), .B1(new_n413), .B2(G902), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n294), .B(new_n600), .C1(new_n358), .C2(new_n360), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  AND4_X1   g434(.A1(new_n492), .A2(new_n618), .A3(new_n495), .A4(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n614), .A2(new_n615), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT34), .B(G104), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  NAND2_X1  g438(.A1(new_n589), .A2(new_n591), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n549), .B1(new_n548), .B2(KEYINPUT20), .ZN(new_n626));
  AOI211_X1 g440(.A(KEYINPUT88), .B(new_n541), .C1(new_n547), .C2(new_n497), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n558), .B1(new_n628), .B2(new_n551), .ZN(new_n629));
  AND4_X1   g443(.A1(new_n615), .A2(new_n621), .A3(new_n625), .A4(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT35), .B(G107), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  NOR2_X1   g446(.A1(new_n472), .A2(new_n473), .ZN(new_n633));
  OR2_X1    g447(.A1(new_n432), .A2(KEYINPUT36), .ZN(new_n634));
  XOR2_X1   g448(.A(new_n633), .B(new_n634), .Z(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n494), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n492), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n365), .A2(new_n602), .A3(new_n618), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT37), .B(G110), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT93), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n638), .B(new_n640), .ZN(G12));
  AOI22_X1  g455(.A1(new_n415), .A2(new_n425), .B1(new_n492), .B2(new_n636), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n542), .A2(new_n550), .A3(new_n551), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n599), .A2(G900), .A3(new_n429), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT94), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n595), .B(KEYINPUT95), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AND4_X1   g461(.A1(new_n559), .A2(new_n643), .A3(new_n625), .A4(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n365), .A2(new_n642), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G128), .ZN(G30));
  XNOR2_X1  g464(.A(new_n647), .B(KEYINPUT39), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n615), .A2(new_n651), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n652), .A2(KEYINPUT40), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n359), .A2(new_n361), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT38), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n294), .A3(new_n625), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n553), .B1(new_n540), .B2(new_n541), .ZN(new_n657));
  AND4_X1   g471(.A1(new_n553), .A2(new_n547), .A3(new_n541), .A4(new_n497), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n558), .B1(new_n628), .B2(new_n659), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n656), .A2(new_n660), .A3(new_n637), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n652), .A2(KEYINPUT40), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n416), .A2(new_n407), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n663), .B1(new_n420), .B2(new_n407), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT96), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT96), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n666), .B(new_n663), .C1(new_n420), .C2(new_n407), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n665), .A2(new_n286), .A3(new_n667), .ZN(new_n668));
  AOI22_X1  g482(.A1(new_n668), .A2(G472), .B1(new_n409), .B2(KEYINPUT32), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n415), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n653), .A2(new_n661), .A3(new_n662), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G143), .ZN(G45));
  INV_X1    g486(.A(new_n647), .ZN(new_n673));
  AOI211_X1 g487(.A(new_n611), .B(new_n673), .C1(new_n555), .C2(new_n559), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n365), .A2(new_n642), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G146), .ZN(G48));
  NOR2_X1   g490(.A1(new_n612), .A2(new_n613), .ZN(new_n677));
  AOI211_X1 g491(.A(KEYINPUT92), .B(new_n611), .C1(new_n555), .C2(new_n559), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n620), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n286), .B1(new_n290), .B2(new_n291), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(G469), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT97), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n681), .A2(new_n682), .A3(new_n364), .A4(new_n292), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n681), .A2(new_n364), .A3(new_n292), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT97), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n496), .A2(new_n426), .A3(new_n683), .A4(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n679), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT41), .B(G113), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT98), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n687), .B(new_n689), .ZN(G15));
  NAND3_X1  g504(.A1(new_n629), .A2(new_n625), .A3(new_n620), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G116), .ZN(G18));
  NAND3_X1  g507(.A1(new_n685), .A2(new_n362), .A3(new_n683), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(new_n602), .A3(new_n642), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  INV_X1    g511(.A(KEYINPUT100), .ZN(new_n698));
  OAI211_X1 g512(.A(new_n294), .B(new_n625), .C1(new_n358), .C2(new_n360), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n698), .B1(new_n660), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n555), .A2(new_n559), .ZN(new_n701));
  INV_X1    g515(.A(new_n699), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n701), .A2(KEYINPUT100), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n685), .A2(new_n683), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n492), .A2(new_n495), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT99), .ZN(new_n708));
  AOI22_X1  g522(.A1(new_n394), .A2(new_n398), .B1(new_n417), .B2(new_n407), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n708), .B1(new_n709), .B2(new_n368), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n417), .A2(new_n407), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n399), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(KEYINPUT99), .A3(new_n367), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n710), .A2(new_n713), .A3(new_n617), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n707), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n704), .A2(new_n600), .A3(new_n706), .A4(new_n715), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT101), .B(G122), .Z(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G24));
  NAND2_X1  g532(.A1(new_n612), .A2(new_n647), .ZN(new_n719));
  INV_X1    g533(.A(new_n714), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n637), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n694), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n328), .ZN(G27));
  NAND2_X1  g537(.A1(new_n496), .A2(new_n426), .ZN(new_n724));
  INV_X1    g538(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n719), .A2(KEYINPUT42), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n654), .A2(new_n295), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n256), .A2(new_n257), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n256), .A2(new_n257), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n215), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n271), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n269), .A2(KEYINPUT12), .A3(new_n215), .ZN(new_n732));
  AOI22_X1  g546(.A1(new_n731), .A2(new_n732), .B1(new_n216), .B2(new_n281), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT102), .B1(new_n733), .B2(new_n204), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT102), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n273), .A2(new_n735), .A3(new_n274), .ZN(new_n736));
  AOI22_X1  g550(.A1(new_n734), .A2(new_n736), .B1(new_n283), .B2(new_n262), .ZN(new_n737));
  OAI21_X1  g551(.A(G469), .B1(new_n737), .B2(G902), .ZN(new_n738));
  AOI21_X1  g552(.A(KEYINPUT103), .B1(new_n738), .B2(new_n292), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n733), .A2(KEYINPUT102), .A3(new_n204), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n735), .B1(new_n273), .B2(new_n274), .ZN(new_n741));
  OAI211_X1 g555(.A(G469), .B(new_n266), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(G469), .A2(G902), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n292), .A2(new_n742), .A3(KEYINPUT103), .A4(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n364), .B(new_n727), .C1(new_n739), .C2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(KEYINPUT104), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT104), .ZN(new_n748));
  INV_X1    g562(.A(new_n364), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n292), .A2(new_n742), .A3(new_n743), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT103), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n749), .B1(new_n752), .B2(new_n744), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n748), .B1(new_n753), .B2(new_n727), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n725), .B(new_n726), .C1(new_n747), .C2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n425), .B1(KEYINPUT32), .B2(new_n409), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n674), .A2(new_n496), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n746), .A2(KEYINPUT104), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n753), .A2(new_n748), .A3(new_n727), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n755), .B1(new_n756), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n213), .ZN(G33));
  OAI211_X1 g577(.A(new_n725), .B(new_n648), .C1(new_n747), .C2(new_n754), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  NAND2_X1  g579(.A1(new_n737), .A2(KEYINPUT45), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n766), .B(G469), .C1(KEYINPUT45), .C2(new_n284), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n743), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT46), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n767), .A2(KEYINPUT46), .A3(new_n743), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(new_n292), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n364), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n774), .A2(new_n651), .A3(new_n727), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n618), .B1(new_n492), .B2(new_n636), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n776), .B(KEYINPUT105), .Z(new_n777));
  NOR2_X1   g591(.A1(new_n701), .A2(new_n611), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT43), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT44), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n775), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n782), .B1(new_n781), .B2(new_n780), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  NAND2_X1  g598(.A1(new_n774), .A2(KEYINPUT47), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n773), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(new_n727), .ZN(new_n789));
  NOR4_X1   g603(.A1(new_n719), .A2(new_n496), .A3(new_n426), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT106), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT100), .B1(new_n701), .B2(new_n702), .ZN(new_n795));
  AOI211_X1 g609(.A(new_n698), .B(new_n699), .C1(new_n555), .C2(new_n559), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n492), .A2(new_n636), .A3(new_n647), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n753), .A2(new_n798), .A3(new_n670), .ZN(new_n799));
  OAI21_X1  g613(.A(KEYINPUT107), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT107), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n492), .A2(new_n636), .A3(new_n647), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(new_n415), .B2(new_n669), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n704), .A2(new_n801), .A3(new_n753), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n365), .B(new_n642), .C1(new_n674), .C2(new_n648), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n722), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n805), .A2(KEYINPUT52), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT52), .B1(new_n805), .B2(new_n808), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n719), .A2(new_n721), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n812), .B1(new_n747), .B2(new_n754), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n789), .A2(new_n625), .A3(new_n673), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(new_n642), .A3(new_n615), .A4(new_n629), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n764), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n758), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(new_n747), .B2(new_n754), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n724), .B1(new_n759), .B2(new_n760), .ZN(new_n819));
  AOI22_X1  g633(.A1(new_n818), .A2(KEYINPUT42), .B1(new_n819), .B2(new_n726), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n715), .A2(new_n600), .A3(new_n683), .A4(new_n685), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n797), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n426), .A2(new_n602), .A3(new_n637), .ZN(new_n823));
  OAI22_X1  g637(.A1(new_n686), .A2(new_n691), .B1(new_n823), .B2(new_n694), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n687), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n555), .A2(new_n559), .A3(new_n625), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(new_n660), .B2(new_n611), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n621), .A2(new_n827), .A3(new_n615), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n828), .A2(new_n603), .A3(new_n638), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n816), .A2(new_n820), .A3(new_n825), .A4(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n794), .B1(new_n811), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT109), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n829), .A2(new_n764), .A3(new_n813), .A4(new_n815), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT110), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n805), .A2(new_n808), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT52), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n805), .A2(new_n808), .A3(KEYINPUT52), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n794), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n614), .A2(new_n725), .A3(new_n620), .A4(new_n706), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n716), .A3(new_n692), .A4(new_n696), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT111), .B1(new_n762), .B2(new_n843), .ZN(new_n844));
  OR3_X1    g658(.A1(new_n762), .A2(new_n843), .A3(KEYINPUT111), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n836), .A2(new_n841), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT109), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n847), .B(new_n794), .C1(new_n811), .C2(new_n830), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n832), .A2(new_n833), .A3(new_n846), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n839), .A2(new_n840), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n834), .A2(new_n762), .A3(new_n843), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n850), .A2(new_n851), .A3(KEYINPUT53), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n831), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT108), .B1(new_n853), .B2(KEYINPUT54), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT108), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n855), .B(new_n833), .C1(new_n831), .C2(new_n852), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n849), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT112), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g673(.A(KEYINPUT112), .B(new_n849), .C1(new_n854), .C2(new_n856), .ZN(new_n860));
  INV_X1    g674(.A(new_n646), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n779), .A2(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n862), .A2(new_n715), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n705), .A2(new_n294), .A3(new_n655), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT50), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n865), .B(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n705), .A2(new_n789), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n862), .A2(new_n637), .A3(new_n720), .A4(new_n868), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n670), .A2(new_n707), .A3(new_n595), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n868), .A2(new_n870), .A3(new_n660), .A4(new_n611), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT51), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n863), .A2(new_n727), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n681), .A2(new_n749), .A3(new_n292), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n785), .A2(new_n787), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n872), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n867), .A2(new_n869), .A3(new_n871), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n757), .A2(new_n496), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n862), .A2(new_n879), .A3(new_n868), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT48), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n614), .A2(new_n868), .A3(new_n870), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n593), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n863), .B2(new_n695), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT114), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n881), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n885), .B1(new_n881), .B2(new_n884), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n877), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n865), .B(KEYINPUT50), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n869), .A2(new_n871), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n874), .B(KEYINPUT113), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n873), .B1(new_n788), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT51), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n859), .A2(new_n860), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n592), .A2(new_n429), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n681), .A2(new_n292), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n899), .A2(KEYINPUT49), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(KEYINPUT49), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n364), .A2(new_n294), .ZN(new_n902));
  NOR4_X1   g716(.A1(new_n655), .A2(new_n900), .A3(new_n901), .A4(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n670), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n903), .A2(new_n496), .A3(new_n904), .A4(new_n778), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n898), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT115), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n898), .A2(KEYINPUT115), .A3(new_n905), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(G75));
  NAND3_X1  g724(.A1(new_n832), .A2(new_n846), .A3(new_n848), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n911), .A2(G210), .A3(G902), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT117), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT56), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n324), .A2(new_n326), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(KEYINPUT116), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n337), .B(KEYINPUT55), .Z(new_n918));
  XOR2_X1   g732(.A(new_n917), .B(new_n918), .Z(new_n919));
  NAND3_X1  g733(.A1(new_n914), .A2(new_n915), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n920), .B1(new_n913), .B2(new_n912), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n919), .B1(new_n912), .B2(new_n915), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n429), .A2(G952), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(G51));
  NAND2_X1  g738(.A1(new_n911), .A2(KEYINPUT54), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(new_n849), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n743), .B(KEYINPUT57), .ZN(new_n928));
  OAI22_X1  g742(.A1(new_n927), .A2(new_n928), .B1(new_n291), .B2(new_n290), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n911), .A2(G902), .ZN(new_n930));
  OR2_X1    g744(.A1(new_n930), .A2(new_n767), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n923), .B1(new_n929), .B2(new_n931), .ZN(G54));
  INV_X1    g746(.A(new_n923), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT58), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n930), .A2(new_n934), .A3(new_n556), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n933), .B1(new_n935), .B2(new_n547), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n936), .B1(new_n547), .B2(new_n935), .ZN(G60));
  NAND2_X1  g751(.A1(new_n859), .A2(new_n860), .ZN(new_n938));
  XNOR2_X1  g752(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n939));
  NAND2_X1  g753(.A1(G478), .A2(G902), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(new_n608), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT120), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n609), .A2(new_n941), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n926), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT119), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT119), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n926), .A2(new_n949), .A3(new_n946), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n923), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n943), .A2(new_n944), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n609), .B1(new_n938), .B2(new_n941), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n949), .B1(new_n926), .B2(new_n946), .ZN(new_n954));
  AOI211_X1 g768(.A(KEYINPUT119), .B(new_n945), .C1(new_n925), .C2(new_n849), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n933), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(KEYINPUT120), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n952), .A2(new_n957), .ZN(G63));
  INV_X1    g772(.A(KEYINPUT122), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n933), .B1(new_n959), .B2(KEYINPUT61), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n479), .B(KEYINPUT60), .Z(new_n961));
  NAND2_X1  g775(.A1(new_n911), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n493), .B(KEYINPUT121), .Z(new_n963));
  AOI21_X1  g777(.A(new_n960), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n635), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n964), .B1(new_n965), .B2(new_n962), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n959), .A2(KEYINPUT61), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n966), .B(new_n967), .ZN(G66));
  OAI21_X1  g782(.A(new_n598), .B1(G224), .B2(new_n429), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT123), .Z(new_n970));
  AND2_X1   g784(.A1(new_n825), .A2(new_n829), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n970), .B1(new_n971), .B2(G953), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n917), .B1(G898), .B2(new_n429), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT124), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT125), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n972), .B(new_n975), .ZN(G69));
  NAND2_X1  g790(.A1(new_n508), .A2(new_n510), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n397), .B(new_n977), .Z(new_n978));
  NAND2_X1  g792(.A1(new_n792), .A2(new_n783), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n671), .A2(new_n808), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(KEYINPUT62), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n981), .A2(KEYINPUT62), .ZN(new_n983));
  INV_X1    g797(.A(new_n827), .ZN(new_n984));
  NOR4_X1   g798(.A1(new_n984), .A2(new_n652), .A3(new_n724), .A4(new_n789), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n980), .A2(new_n982), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n978), .B1(new_n987), .B2(G953), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n429), .A2(G900), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n774), .A2(new_n651), .A3(new_n704), .A4(new_n879), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n820), .A2(new_n990), .A3(new_n764), .A4(new_n808), .ZN(new_n991));
  OR3_X1    g805(.A1(new_n979), .A2(KEYINPUT126), .A3(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(KEYINPUT126), .B1(new_n979), .B2(new_n991), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n989), .B1(new_n994), .B2(new_n429), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n988), .B1(new_n995), .B2(new_n978), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n429), .B1(G227), .B2(G900), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(G72));
  NAND2_X1  g812(.A1(new_n987), .A2(new_n971), .ZN(new_n999));
  NAND2_X1  g813(.A1(G472), .A2(G902), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT63), .Z(new_n1001));
  AOI211_X1 g815(.A(new_n407), .B(new_n420), .C1(new_n999), .C2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n420), .A2(new_n407), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n992), .A2(new_n971), .A3(new_n993), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1003), .B1(new_n1004), .B2(new_n1001), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n385), .A2(new_n393), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1001), .B1(new_n421), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1007), .B1(new_n831), .B2(new_n852), .ZN(new_n1008));
  NOR4_X1   g822(.A1(new_n1002), .A2(new_n923), .A3(new_n1005), .A4(new_n1008), .ZN(G57));
endmodule


