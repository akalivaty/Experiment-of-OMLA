//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 1 0 1 1 1 1 1 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G119), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G128), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT24), .B(G110), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n194));
  NOR3_X1   g008(.A1(new_n194), .A2(new_n189), .A3(G128), .ZN(new_n195));
  OR2_X1    g009(.A1(new_n195), .A2(KEYINPUT71), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT72), .ZN(new_n197));
  AOI22_X1  g011(.A1(new_n197), .A2(new_n194), .B1(new_n187), .B2(G119), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n198), .B1(new_n197), .B2(new_n194), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n195), .A2(KEYINPUT71), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n196), .A2(new_n199), .A3(new_n190), .A4(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n193), .B1(new_n201), .B2(G110), .ZN(new_n202));
  XNOR2_X1  g016(.A(G125), .B(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT16), .ZN(new_n205));
  INV_X1    g019(.A(G140), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G125), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(G146), .A3(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n203), .A2(new_n209), .ZN(new_n210));
  AND2_X1   g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n191), .A2(new_n192), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n212), .B1(new_n201), .B2(G110), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n206), .A2(G125), .ZN(new_n214));
  INV_X1    g028(.A(G125), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G140), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n207), .B1(new_n217), .B2(new_n205), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(new_n209), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n208), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n202), .A2(new_n211), .B1(new_n213), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT22), .B(G137), .ZN(new_n222));
  INV_X1    g036(.A(G953), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(G221), .A3(G234), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n222), .B(new_n224), .ZN(new_n225));
  XOR2_X1   g039(.A(new_n225), .B(KEYINPUT73), .Z(new_n226));
  OR2_X1    g040(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n221), .A2(new_n225), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G902), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(KEYINPUT25), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n233), .B1(new_n229), .B2(G902), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G217), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n236), .B1(G234), .B2(new_n231), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n237), .A2(G902), .ZN(new_n238));
  XOR2_X1   g052(.A(new_n238), .B(KEYINPUT74), .Z(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n235), .A2(new_n237), .B1(new_n240), .B2(new_n230), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT28), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n209), .A2(G143), .ZN(new_n244));
  INV_X1    g058(.A(G143), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G146), .ZN(new_n246));
  OR2_X1    g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  NAND2_X1  g061(.A1(KEYINPUT0), .A2(G128), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n244), .A2(new_n246), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n244), .A2(new_n246), .A3(new_n248), .ZN(new_n250));
  OR2_X1    g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G134), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT11), .B1(new_n252), .B2(G137), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n254));
  INV_X1    g068(.A(G137), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(G134), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G131), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT65), .B1(new_n255), .B2(G134), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT65), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(new_n252), .A3(G137), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n257), .A2(new_n258), .A3(new_n259), .A4(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n259), .A2(new_n261), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n258), .B1(new_n264), .B2(new_n257), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n251), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n187), .A2(KEYINPUT1), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(new_n244), .A3(new_n246), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n187), .B1(new_n244), .B2(KEYINPUT1), .ZN(new_n269));
  XNOR2_X1  g083(.A(G143), .B(G146), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n252), .A2(G137), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n255), .A2(G134), .ZN(new_n273));
  OAI21_X1  g087(.A(G131), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n262), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n266), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(KEYINPUT2), .A2(G113), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT66), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT66), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n279), .B1(KEYINPUT2), .B2(G113), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(KEYINPUT2), .A2(G113), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(G116), .B(G119), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n281), .A2(new_n282), .A3(new_n284), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n243), .B1(new_n276), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(G237), .A2(G953), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G210), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n291), .B(KEYINPUT27), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT26), .B(G101), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT29), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT67), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n262), .A2(new_n271), .A3(new_n298), .A4(new_n274), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n249), .A2(new_n250), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n257), .A2(new_n259), .A3(new_n261), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G131), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n301), .B1(new_n303), .B2(new_n262), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n300), .A2(new_n304), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n286), .A2(new_n287), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n275), .A2(KEYINPUT67), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n305), .A2(KEYINPUT68), .A3(new_n306), .A4(new_n307), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n307), .A2(new_n266), .A3(new_n306), .A4(new_n299), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT68), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n305), .A2(new_n307), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n308), .A2(new_n311), .B1(new_n312), .B2(new_n288), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n289), .B(new_n297), .C1(new_n313), .C2(new_n243), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT70), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n312), .A2(new_n288), .ZN(new_n316));
  AND2_X1   g130(.A1(new_n309), .A2(new_n310), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n309), .A2(new_n310), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT28), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT70), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n320), .A2(new_n321), .A3(new_n289), .A4(new_n297), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n315), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n308), .A2(new_n311), .A3(KEYINPUT28), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n276), .A2(new_n288), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n324), .A2(new_n294), .A3(new_n325), .A4(new_n289), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n296), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n307), .A2(new_n266), .A3(new_n299), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT64), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n329), .B1(new_n266), .B2(new_n275), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT30), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT30), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n276), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n288), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n308), .A2(new_n311), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n294), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n231), .B1(new_n327), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(G472), .B1(new_n323), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n334), .A2(new_n294), .A3(new_n335), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(KEYINPUT31), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n324), .A2(new_n325), .A3(new_n289), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n295), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT31), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n334), .A2(new_n343), .A3(new_n294), .A4(new_n335), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n340), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(G472), .A2(G902), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(KEYINPUT32), .A3(new_n346), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n338), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n346), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT69), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT32), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT69), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n345), .A2(new_n352), .A3(new_n346), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n350), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n242), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT9), .B(G234), .ZN(new_n356));
  OAI21_X1  g170(.A(G221), .B1(new_n356), .B2(G902), .ZN(new_n357));
  INV_X1    g171(.A(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G101), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT75), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT3), .ZN(new_n361));
  INV_X1    g175(.A(G104), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n360), .A2(new_n361), .B1(new_n362), .B2(G107), .ZN(new_n363));
  NAND2_X1  g177(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n364));
  NOR3_X1   g178(.A1(new_n364), .A2(new_n362), .A3(G107), .ZN(new_n365));
  INV_X1    g179(.A(G107), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n366), .A2(G104), .B1(KEYINPUT75), .B2(KEYINPUT3), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n359), .B(new_n363), .C1(new_n365), .C2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n362), .A2(G107), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n366), .A2(G104), .ZN(new_n370));
  OAI21_X1  g184(.A(G101), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT78), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n368), .A2(new_n374), .A3(new_n371), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  OR2_X1    g190(.A1(new_n269), .A2(new_n270), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n377), .A2(new_n268), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n270), .ZN(new_n380));
  OAI211_X1 g194(.A(KEYINPUT76), .B(KEYINPUT1), .C1(new_n245), .C2(G146), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G128), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT76), .B1(new_n244), .B2(KEYINPUT1), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n380), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT77), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT77), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n386), .B(new_n380), .C1(new_n382), .C2(new_n383), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n268), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n372), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n379), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n263), .A2(new_n265), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(KEYINPUT12), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT12), .ZN(new_n395));
  AOI211_X1 g209(.A(new_n395), .B(new_n392), .C1(new_n379), .C2(new_n390), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G110), .B(G140), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n223), .A2(G227), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n399), .B(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT10), .B1(new_n388), .B2(new_n389), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n363), .B1(new_n365), .B2(new_n367), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G101), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(KEYINPUT4), .A3(new_n368), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n403), .A2(new_n406), .A3(G101), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n405), .A2(new_n251), .A3(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n402), .A2(new_n408), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n271), .A2(KEYINPUT10), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n373), .A2(new_n410), .A3(new_n375), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT79), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT79), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n373), .A2(new_n410), .A3(new_n413), .A4(new_n375), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n409), .A2(new_n415), .A3(new_n392), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT80), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT80), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n409), .A2(new_n415), .A3(new_n418), .A4(new_n392), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n401), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT81), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n398), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI211_X1 g236(.A(KEYINPUT81), .B(new_n401), .C1(new_n417), .C2(new_n419), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n417), .A2(new_n419), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n409), .A2(new_n415), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n393), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n401), .ZN(new_n428));
  OAI22_X1  g242(.A1(new_n422), .A2(new_n423), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G469), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n430), .A3(new_n231), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n430), .A2(new_n231), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n424), .A2(new_n398), .ZN(new_n433));
  AOI22_X1  g247(.A1(new_n433), .A2(new_n401), .B1(new_n420), .B2(new_n426), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n432), .B1(new_n434), .B2(G469), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n358), .B1(new_n431), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G237), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(new_n223), .A3(G214), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n245), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n290), .A2(G143), .A3(G214), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(KEYINPUT18), .A2(G131), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n217), .A2(G146), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n442), .A2(new_n443), .B1(new_n210), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n443), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n441), .A2(KEYINPUT85), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(KEYINPUT85), .B1(new_n441), .B2(new_n446), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n445), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n218), .A2(new_n209), .ZN(new_n451));
  AOI21_X1  g265(.A(G146), .B1(new_n204), .B2(new_n207), .ZN(new_n452));
  OAI21_X1  g266(.A(KEYINPUT87), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT87), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n219), .A2(new_n454), .A3(new_n208), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n441), .A2(KEYINPUT17), .A3(G131), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n441), .A2(G131), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n439), .A2(new_n258), .A3(new_n440), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n457), .B1(new_n460), .B2(KEYINPUT17), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n450), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(G113), .B(G122), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(new_n362), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n464), .B(new_n450), .C1(new_n456), .C2(new_n461), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n231), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(G475), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT20), .ZN(new_n471));
  NOR2_X1   g285(.A1(G475), .A2(G902), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT86), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n444), .A2(new_n210), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n474), .B1(new_n441), .B2(new_n446), .ZN(new_n475));
  INV_X1    g289(.A(new_n449), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n475), .B1(new_n476), .B2(new_n447), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n203), .A2(KEYINPUT19), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n203), .A2(KEYINPUT19), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n209), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n460), .A2(new_n481), .A3(new_n208), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n473), .B(new_n465), .C1(new_n477), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n467), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT19), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n217), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(G146), .B1(new_n486), .B2(new_n478), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n451), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n460), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n450), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n473), .B1(new_n490), .B2(new_n465), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n471), .B(new_n472), .C1(new_n484), .C2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n476), .A2(new_n447), .ZN(new_n494));
  AOI22_X1  g308(.A1(new_n494), .A2(new_n445), .B1(new_n488), .B2(new_n460), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT86), .B1(new_n495), .B2(new_n464), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(new_n467), .A3(new_n483), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n471), .B1(new_n497), .B2(new_n472), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n470), .B1(new_n493), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G952), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n500), .A2(G953), .ZN(new_n501));
  INV_X1    g315(.A(G234), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n501), .B1(new_n502), .B2(new_n437), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AOI211_X1 g318(.A(new_n231), .B(new_n223), .C1(G234), .C2(G237), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT21), .B(G898), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n356), .A2(new_n236), .A3(G953), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G116), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G122), .ZN(new_n511));
  INV_X1    g325(.A(G122), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G116), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(new_n513), .A3(new_n366), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n245), .A2(G128), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n187), .A2(G143), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n515), .A2(new_n516), .A3(new_n252), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n252), .B1(new_n515), .B2(new_n516), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n514), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT14), .B1(new_n512), .B2(G116), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n512), .A2(G116), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT89), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT14), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n510), .B2(G122), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT89), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n511), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT90), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n527), .B1(new_n511), .B2(KEYINPUT14), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n521), .A2(KEYINPUT90), .A3(new_n523), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n522), .A2(new_n526), .A3(new_n528), .A4(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n519), .B1(G107), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n515), .A2(new_n516), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT13), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n516), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n532), .A2(new_n534), .A3(G134), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n515), .B(new_n516), .C1(new_n533), .C2(new_n252), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT88), .ZN(new_n538));
  INV_X1    g352(.A(new_n514), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n366), .B1(new_n511), .B2(new_n513), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n511), .A2(new_n513), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G107), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(KEYINPUT88), .A3(new_n514), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n537), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n509), .B1(new_n531), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n530), .A2(G107), .ZN(new_n547));
  INV_X1    g361(.A(new_n519), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n535), .A2(new_n536), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n539), .A2(new_n538), .A3(new_n540), .ZN(new_n551));
  AOI21_X1  g365(.A(KEYINPUT88), .B1(new_n543), .B2(new_n514), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n549), .A2(new_n553), .A3(new_n508), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n546), .A2(new_n554), .A3(KEYINPUT91), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n549), .A2(new_n553), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT91), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n556), .A2(new_n557), .A3(new_n509), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(new_n231), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(G478), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n560), .A2(KEYINPUT15), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n559), .B(new_n561), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n499), .A2(new_n507), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(G214), .B1(G237), .B2(G902), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT5), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(new_n189), .A3(G116), .ZN(new_n567));
  OAI211_X1 g381(.A(G113), .B(new_n567), .C1(new_n285), .C2(new_n566), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n373), .A2(new_n287), .A3(new_n375), .A4(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n405), .A2(new_n288), .A3(new_n407), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(G110), .B(G122), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n574), .A2(KEYINPUT6), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n301), .A2(G125), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(G125), .B2(new_n271), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n223), .A2(G224), .ZN(new_n579));
  XOR2_X1   g393(.A(new_n579), .B(KEYINPUT82), .Z(new_n580));
  XNOR2_X1  g394(.A(new_n578), .B(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT6), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n571), .A2(new_n582), .A3(new_n573), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n576), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT84), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n579), .A2(KEYINPUT7), .ZN(new_n586));
  OAI221_X1 g400(.A(new_n577), .B1(new_n585), .B2(new_n586), .C1(G125), .C2(new_n271), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n586), .B1(new_n577), .B2(new_n585), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n578), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n575), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  XOR2_X1   g404(.A(new_n572), .B(KEYINPUT8), .Z(new_n591));
  NAND2_X1  g405(.A1(new_n568), .A2(new_n287), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n372), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n591), .B1(new_n569), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(KEYINPUT83), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT83), .ZN(new_n596));
  AOI211_X1 g410(.A(new_n596), .B(new_n591), .C1(new_n569), .C2(new_n593), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n590), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n584), .A2(new_n598), .A3(new_n231), .ZN(new_n599));
  OAI21_X1  g413(.A(G210), .B1(G237), .B2(G902), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n584), .A2(new_n598), .A3(new_n231), .A4(new_n600), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n565), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n563), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n355), .A2(new_n436), .A3(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  INV_X1    g422(.A(new_n436), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n345), .A2(new_n231), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(KEYINPUT92), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT92), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n345), .A2(new_n612), .A3(new_n231), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n611), .A2(G472), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n353), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n352), .B1(new_n345), .B2(new_n346), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n609), .A2(new_n618), .A3(new_n242), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT33), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n555), .A2(new_n620), .A3(new_n558), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n560), .A2(G902), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT93), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n620), .B1(new_n556), .B2(new_n509), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n623), .B1(new_n624), .B2(new_n554), .ZN(new_n625));
  AND4_X1   g439(.A1(new_n623), .A2(new_n546), .A3(new_n554), .A4(KEYINPUT33), .ZN(new_n626));
  OAI211_X1 g440(.A(new_n621), .B(new_n622), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT94), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n624), .A2(new_n623), .A3(new_n554), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n546), .A2(new_n554), .A3(KEYINPUT33), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(KEYINPUT93), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n633), .A2(KEYINPUT94), .A3(new_n621), .A4(new_n622), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n629), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT95), .B(G478), .Z(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n559), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT96), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n635), .A2(KEYINPUT97), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT97), .B1(new_n635), .B2(new_n640), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n499), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n602), .A2(new_n603), .ZN(new_n644));
  INV_X1    g458(.A(new_n507), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(new_n564), .A3(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n619), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT34), .B(G104), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G6));
  OAI21_X1  g464(.A(new_n470), .B1(KEYINPUT98), .B2(new_n492), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n493), .A2(new_n498), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n651), .B1(KEYINPUT98), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n562), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n646), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n619), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT35), .B(G107), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G9));
  AOI211_X1 g472(.A(new_n358), .B(new_n605), .C1(new_n431), .C2(new_n435), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT36), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n226), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n221), .B(new_n661), .ZN(new_n662));
  AOI22_X1  g476(.A1(new_n235), .A2(new_n237), .B1(new_n240), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n614), .A2(new_n617), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT37), .B(G110), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  AOI21_X1  g482(.A(new_n663), .B1(new_n348), .B2(new_n354), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT99), .B(G900), .Z(new_n670));
  NAND2_X1  g484(.A1(new_n505), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n654), .B1(new_n503), .B2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n669), .A2(new_n436), .A3(new_n604), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  NAND2_X1  g488(.A1(new_n671), .A2(new_n503), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT39), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n609), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n679), .A2(KEYINPUT40), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(KEYINPUT40), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n231), .B1(new_n319), .B2(new_n294), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n295), .B1(new_n334), .B2(new_n335), .ZN(new_n683));
  OAI21_X1  g497(.A(G472), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n347), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n354), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n663), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n644), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n499), .A2(new_n562), .ZN(new_n691));
  NOR4_X1   g505(.A1(new_n687), .A2(new_n565), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n680), .A2(new_n681), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G143), .ZN(G45));
  OAI211_X1 g508(.A(new_n499), .B(new_n675), .C1(new_n641), .C2(new_n642), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT101), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n635), .A2(new_n640), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT97), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n635), .A2(new_n640), .A3(KEYINPUT97), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n702), .A2(KEYINPUT101), .A3(new_n499), .A4(new_n675), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT102), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n697), .A2(new_n703), .A3(new_n704), .A4(new_n604), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n705), .A2(new_n436), .A3(new_n669), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n697), .A2(new_n703), .A3(new_n604), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT102), .ZN(new_n708));
  AOI21_X1  g522(.A(KEYINPUT103), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n669), .A2(new_n436), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n708), .A2(new_n710), .A3(KEYINPUT103), .A4(new_n705), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n209), .ZN(G48));
  AND3_X1   g528(.A1(new_n429), .A2(new_n430), .A3(new_n231), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n430), .B1(new_n429), .B2(new_n231), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n715), .A2(new_n716), .A3(new_n358), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n355), .A3(new_n647), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT41), .B(G113), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G15));
  NAND3_X1  g534(.A1(new_n717), .A2(new_n355), .A3(new_n655), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G116), .ZN(G18));
  NAND3_X1  g536(.A1(new_n717), .A2(new_n669), .A3(new_n606), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G119), .ZN(G21));
  NOR2_X1   g538(.A1(new_n646), .A2(new_n691), .ZN(new_n725));
  INV_X1    g539(.A(new_n289), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n726), .B1(new_n319), .B2(KEYINPUT28), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n340), .B(new_n344), .C1(new_n727), .C2(new_n294), .ZN(new_n728));
  AOI22_X1  g542(.A1(new_n610), .A2(G472), .B1(new_n346), .B2(new_n728), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n725), .A2(new_n729), .A3(new_n241), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n717), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G122), .ZN(G24));
  NAND2_X1  g546(.A1(new_n717), .A2(new_n604), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n697), .A2(new_n703), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n728), .A2(new_n346), .ZN(new_n736));
  INV_X1    g550(.A(G472), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n737), .B1(new_n345), .B2(new_n231), .ZN(new_n738));
  NOR3_X1   g552(.A1(new_n736), .A2(new_n663), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n734), .A2(new_n735), .A3(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  INV_X1    g555(.A(new_n347), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT32), .B1(new_n345), .B2(new_n346), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT104), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n743), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT104), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n746), .A3(new_n347), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n744), .A2(new_n747), .A3(new_n338), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n241), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n602), .A2(new_n603), .A3(new_n357), .A4(new_n564), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n750), .B1(new_n431), .B2(new_n435), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n697), .A3(new_n703), .ZN(new_n752));
  OAI21_X1  g566(.A(KEYINPUT42), .B1(new_n749), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT42), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n735), .A2(new_n754), .A3(new_n355), .A4(new_n751), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G131), .ZN(G33));
  NAND2_X1  g571(.A1(new_n348), .A2(new_n354), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n758), .A2(new_n751), .A3(new_n672), .A4(new_n241), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G134), .ZN(G36));
  NAND3_X1  g574(.A1(new_n405), .A2(new_n251), .A3(new_n407), .ZN(new_n761));
  INV_X1    g575(.A(new_n268), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n762), .B1(new_n384), .B2(KEYINPUT77), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n372), .B1(new_n763), .B2(new_n387), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n761), .B1(new_n764), .B2(KEYINPUT10), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(new_n412), .B2(new_n414), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n418), .B1(new_n766), .B2(new_n392), .ZN(new_n767));
  INV_X1    g581(.A(new_n419), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n426), .B(new_n428), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n397), .B1(new_n419), .B2(new_n417), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n769), .B(KEYINPUT45), .C1(new_n428), .C2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT105), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n433), .A2(new_n401), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(KEYINPUT105), .A3(KEYINPUT45), .A4(new_n769), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n769), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n430), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n432), .B1(new_n776), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n431), .B1(new_n780), .B2(KEYINPUT46), .ZN(new_n781));
  OAI21_X1  g595(.A(G469), .B1(new_n434), .B2(KEYINPUT45), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n782), .B1(new_n773), .B2(new_n775), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT46), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n783), .A2(new_n784), .A3(new_n432), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n357), .B1(new_n781), .B2(new_n785), .ZN(new_n786));
  OR3_X1    g600(.A1(new_n786), .A2(KEYINPUT106), .A3(new_n677), .ZN(new_n787));
  OAI21_X1  g601(.A(KEYINPUT106), .B1(new_n786), .B2(new_n677), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n499), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n790), .B1(new_n641), .B2(new_n642), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT43), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT43), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n702), .A2(new_n793), .A3(new_n790), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n618), .A2(new_n792), .A3(new_n664), .A4(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT44), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n644), .A2(new_n565), .ZN(new_n797));
  XOR2_X1   g611(.A(new_n797), .B(KEYINPUT107), .Z(new_n798));
  NAND3_X1  g612(.A1(new_n789), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G137), .ZN(G39));
  INV_X1    g614(.A(KEYINPUT47), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n786), .A2(new_n801), .ZN(new_n802));
  OAI211_X1 g616(.A(KEYINPUT47), .B(new_n357), .C1(new_n781), .C2(new_n785), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n797), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n758), .A2(new_n241), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n804), .A2(new_n735), .A3(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G140), .ZN(G42));
  OR4_X1    g622(.A1(new_n242), .A2(new_n791), .A3(new_n358), .A4(new_n565), .ZN(new_n809));
  XOR2_X1   g623(.A(new_n809), .B(KEYINPUT108), .Z(new_n810));
  INV_X1    g624(.A(new_n686), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n715), .A2(new_n716), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT49), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n810), .A2(new_n811), .A3(new_n690), .A4(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n758), .A2(new_n647), .A3(new_n241), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n815), .A2(new_n717), .B1(new_n659), .B2(new_n665), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n758), .A2(new_n655), .A3(new_n241), .ZN(new_n817));
  AOI211_X1 g631(.A(new_n605), .B(new_n663), .C1(new_n348), .C2(new_n354), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n717), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n614), .A2(new_n617), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n700), .A2(new_n499), .A3(new_n701), .ZN(new_n821));
  INV_X1    g635(.A(new_n646), .ZN(new_n822));
  INV_X1    g636(.A(new_n562), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n790), .A2(new_n823), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n820), .A2(new_n825), .A3(new_n241), .A4(new_n436), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n659), .A2(new_n355), .B1(new_n717), .B2(new_n730), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n816), .A2(new_n819), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n751), .A2(new_n697), .A3(new_n703), .A4(new_n739), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n759), .A2(new_n829), .ZN(new_n830));
  AND4_X1   g644(.A1(new_n823), .A2(new_n797), .A3(new_n653), .A4(new_n675), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n669), .A2(new_n436), .A3(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n830), .A2(new_n753), .A3(new_n755), .A4(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT109), .B1(new_n828), .B2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n666), .A2(new_n718), .A3(new_n607), .A4(new_n731), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n826), .A2(new_n721), .A3(new_n723), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT109), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n832), .A2(new_n759), .A3(new_n829), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n837), .A2(new_n756), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n834), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n604), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n691), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n843), .A2(new_n675), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n844), .A2(new_n436), .A3(new_n686), .A4(new_n663), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n735), .A2(new_n739), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n673), .B(new_n845), .C1(new_n846), .C2(new_n733), .ZN(new_n847));
  INV_X1    g661(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n848), .B1(new_n709), .B2(new_n712), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT52), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n708), .A2(new_n710), .A3(new_n705), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT103), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n847), .B1(new_n853), .B2(new_n711), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT52), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n841), .A2(new_n850), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(KEYINPUT53), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT110), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n855), .B1(new_n849), .B2(new_n860), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n854), .A2(KEYINPUT110), .A3(KEYINPUT52), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n859), .B(new_n841), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n858), .A2(new_n863), .A3(KEYINPUT54), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n857), .A2(new_n859), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n837), .A2(new_n756), .A3(new_n839), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n859), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(new_n861), .B2(new_n862), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n865), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n812), .A2(new_n358), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n802), .A2(new_n803), .A3(new_n872), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n242), .A2(new_n736), .A3(new_n738), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n792), .A3(new_n794), .A4(new_n504), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n876), .A2(new_n798), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n792), .A2(new_n794), .A3(new_n504), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n429), .A2(new_n231), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(G469), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n881), .A2(new_n357), .A3(new_n431), .A4(new_n797), .ZN(new_n882));
  INV_X1    g696(.A(new_n739), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n879), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n354), .A2(new_n685), .A3(new_n241), .A4(new_n504), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n702), .A2(new_n499), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n882), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT112), .B1(new_n884), .B2(new_n888), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n792), .A2(new_n794), .A3(new_n504), .ZN(new_n890));
  INV_X1    g704(.A(new_n882), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n890), .A2(new_n891), .A3(new_n739), .ZN(new_n892));
  INV_X1    g706(.A(new_n885), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n893), .A3(new_n886), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT112), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n889), .A2(new_n896), .A3(KEYINPUT51), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n690), .A2(new_n565), .ZN(new_n898));
  NOR4_X1   g712(.A1(new_n898), .A2(new_n715), .A3(new_n716), .A4(new_n358), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT50), .B1(new_n876), .B2(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n812), .A2(new_n357), .A3(new_n565), .A4(new_n690), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT50), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n901), .A2(new_n875), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n878), .A2(new_n897), .A3(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n879), .A2(new_n882), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n748), .A2(new_n241), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT48), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT48), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n907), .A2(new_n908), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  AOI211_X1 g727(.A(new_n500), .B(G953), .C1(new_n876), .C2(new_n734), .ZN(new_n914));
  OR3_X1    g728(.A1(new_n882), .A2(new_n885), .A3(new_n643), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n906), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g732(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n904), .B1(new_n873), .B2(new_n877), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n884), .A2(new_n888), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n918), .A2(new_n923), .A3(KEYINPUT113), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT113), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n878), .A2(new_n905), .A3(new_n922), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n919), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n916), .B1(new_n921), .B2(new_n897), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT114), .B1(new_n871), .B2(new_n930), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n930), .A2(KEYINPUT114), .A3(new_n864), .A4(new_n870), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n500), .A2(new_n223), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n814), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT115), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI211_X1 g751(.A(KEYINPUT115), .B(new_n814), .C1(new_n931), .C2(new_n934), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(G75));
  NOR2_X1   g753(.A1(new_n223), .A2(G952), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT56), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n857), .A2(new_n859), .ZN(new_n943));
  INV_X1    g757(.A(new_n868), .ZN(new_n944));
  OAI21_X1  g758(.A(G902), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(G210), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n942), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n576), .A2(new_n583), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT116), .Z(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT55), .Z(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT117), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(new_n581), .Z(new_n952));
  OAI21_X1  g766(.A(new_n941), .B1(new_n947), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n947), .A2(new_n952), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT118), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n947), .A2(KEYINPUT118), .A3(new_n952), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n953), .B1(new_n956), .B2(new_n957), .ZN(G51));
  OAI21_X1  g772(.A(KEYINPUT54), .B1(new_n943), .B2(new_n944), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n870), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n432), .B(KEYINPUT57), .Z(new_n962));
  OAI21_X1  g776(.A(new_n429), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n783), .B(KEYINPUT119), .Z(new_n964));
  OR2_X1    g778(.A1(new_n945), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n940), .B1(new_n963), .B2(new_n965), .ZN(G54));
  INV_X1    g780(.A(new_n945), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n967), .A2(KEYINPUT58), .A3(G475), .ZN(new_n968));
  INV_X1    g782(.A(new_n497), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n968), .A2(new_n969), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n970), .A2(new_n971), .A3(new_n940), .ZN(G60));
  NAND2_X1  g786(.A1(G478), .A2(G902), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT59), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n633), .A2(new_n621), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n940), .B1(new_n960), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n864), .A2(new_n870), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n974), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n633), .A2(new_n621), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n976), .A2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT120), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n976), .A2(new_n980), .A3(KEYINPUT120), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(G63));
  NAND2_X1  g799(.A1(G217), .A2(G902), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT60), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n987), .B1(new_n865), .B2(new_n868), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n940), .B1(new_n988), .B2(new_n662), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n662), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n990), .A2(KEYINPUT121), .ZN(new_n991));
  OAI221_X1 g805(.A(new_n989), .B1(new_n230), .B2(new_n988), .C1(new_n991), .C2(KEYINPUT61), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n991), .A2(KEYINPUT61), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n989), .B1(new_n230), .B2(new_n988), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n992), .A2(new_n995), .ZN(G66));
  INV_X1    g810(.A(G224), .ZN(new_n997));
  OAI21_X1  g811(.A(G953), .B1(new_n506), .B2(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n998), .B1(new_n837), .B2(G953), .ZN(new_n999));
  INV_X1    g813(.A(new_n949), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n1000), .B1(G898), .B2(new_n223), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n999), .B(new_n1001), .ZN(G69));
  INV_X1    g816(.A(KEYINPUT123), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n740), .A2(new_n673), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n713), .A2(new_n1004), .ZN(new_n1005));
  AND3_X1   g819(.A1(new_n1005), .A2(new_n756), .A3(new_n759), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n799), .A2(new_n807), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n789), .A2(new_n908), .A3(new_n843), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1006), .A2(new_n1007), .A3(new_n223), .A4(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n331), .A2(new_n333), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n479), .A2(new_n480), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1013), .B1(G900), .B2(G953), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1003), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n223), .B1(G227), .B2(G900), .ZN(new_n1016));
  NOR3_X1   g830(.A1(new_n1015), .A2(KEYINPUT124), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  OAI21_X1  g832(.A(KEYINPUT124), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT122), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1005), .A2(new_n693), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1020), .B1(new_n1021), .B2(KEYINPUT62), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT62), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n1005), .A2(KEYINPUT122), .A3(new_n1023), .A4(new_n693), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  AND2_X1   g839(.A1(new_n821), .A2(new_n824), .ZN(new_n1026));
  NAND4_X1  g840(.A1(new_n678), .A2(new_n355), .A3(new_n797), .A4(new_n1026), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n799), .A2(new_n807), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1028), .B1(KEYINPUT62), .B2(new_n1021), .ZN(new_n1029));
  AOI21_X1  g843(.A(G953), .B1(new_n1025), .B2(new_n1029), .ZN(new_n1030));
  OR2_X1    g844(.A1(new_n1030), .A2(new_n1012), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1009), .A2(new_n1014), .ZN(new_n1032));
  AOI22_X1  g846(.A1(new_n1018), .A2(new_n1019), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1019), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1032), .B1(new_n1030), .B2(new_n1012), .ZN(new_n1035));
  NOR3_X1   g849(.A1(new_n1034), .A2(new_n1035), .A3(new_n1017), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n1033), .A2(new_n1036), .ZN(G72));
  XNOR2_X1  g851(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1038));
  NOR2_X1   g852(.A1(new_n737), .A2(new_n231), .ZN(new_n1039));
  XOR2_X1   g853(.A(new_n1038), .B(new_n1039), .Z(new_n1040));
  INV_X1    g854(.A(new_n336), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1040), .B1(new_n1041), .B2(new_n339), .ZN(new_n1042));
  NAND3_X1  g856(.A1(new_n858), .A2(new_n863), .A3(new_n1042), .ZN(new_n1043));
  AND2_X1   g857(.A1(new_n1043), .A2(KEYINPUT126), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n1043), .A2(KEYINPUT126), .ZN(new_n1045));
  OR2_X1    g859(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AND3_X1   g860(.A1(new_n1025), .A2(new_n837), .A3(new_n1029), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n683), .B1(new_n1047), .B2(new_n1040), .ZN(new_n1048));
  INV_X1    g862(.A(new_n1040), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1049), .B1(new_n1050), .B2(new_n828), .ZN(new_n1051));
  AND3_X1   g865(.A1(new_n334), .A2(new_n295), .A3(new_n335), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n940), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n1046), .A2(new_n1048), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g868(.A(KEYINPUT127), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND4_X1  g870(.A1(new_n1046), .A2(KEYINPUT127), .A3(new_n1048), .A4(new_n1053), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1056), .A2(new_n1057), .ZN(G57));
endmodule


