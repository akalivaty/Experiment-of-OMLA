//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT11), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G197gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(new_n207), .B(KEYINPUT12), .Z(new_n208));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT16), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n209), .B1(new_n210), .B2(G1gat), .ZN(new_n211));
  INV_X1    g010(.A(G8gat), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n212), .A2(KEYINPUT92), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n211), .B(new_n213), .C1(G1gat), .C2(new_n209), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n212), .A2(KEYINPUT92), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT14), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G29gat), .B2(G36gat), .ZN(new_n218));
  OR3_X1    g017(.A1(new_n217), .A2(G29gat), .A3(G36gat), .ZN(new_n219));
  XOR2_X1   g018(.A(KEYINPUT91), .B(G29gat), .Z(new_n220));
  INV_X1    g019(.A(G36gat), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n218), .B(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G43gat), .B(G50gat), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n223), .A2(KEYINPUT15), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n223), .B(KEYINPUT15), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n227), .A2(new_n222), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n216), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT17), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(new_n226), .B2(new_n228), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n225), .B(KEYINPUT17), .C1(new_n222), .C2(new_n227), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n230), .B1(new_n234), .B2(KEYINPUT93), .ZN(new_n235));
  NAND2_X1  g034(.A1(G229gat), .A2(G233gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT93), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n216), .A2(new_n232), .A3(new_n237), .A4(new_n233), .ZN(new_n238));
  NAND4_X1  g037(.A1(new_n235), .A2(KEYINPUT18), .A3(new_n236), .A4(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n216), .B(new_n229), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n236), .B(KEYINPUT13), .Z(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n234), .A2(KEYINPUT93), .ZN(new_n245));
  INV_X1    g044(.A(new_n230), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n245), .A2(new_n236), .A3(new_n238), .A4(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT94), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT94), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n235), .A2(new_n249), .A3(new_n236), .A4(new_n238), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  XOR2_X1   g050(.A(KEYINPUT95), .B(KEYINPUT18), .Z(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n208), .B(new_n244), .C1(new_n251), .C2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n208), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n253), .B1(new_n248), .B2(new_n250), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n255), .B1(new_n256), .B2(new_n243), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT85), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n261), .A2(KEYINPUT28), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT27), .B(G183gat), .ZN(new_n263));
  INV_X1    g062(.A(G190gat), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G183gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT27), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT27), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G183gat), .ZN(new_n269));
  AND4_X1   g068(.A1(new_n264), .A2(new_n262), .A3(new_n267), .A4(new_n269), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n265), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT26), .ZN(new_n272));
  INV_X1    g071(.A(G176gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n272), .A2(new_n204), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G183gat), .A2(G190gat), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n204), .A2(new_n273), .A3(KEYINPUT23), .ZN(new_n280));
  AND2_X1   g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n204), .A2(new_n273), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT23), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT66), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT24), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n278), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n266), .A2(new_n264), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n290), .A2(new_n286), .ZN(new_n291));
  OAI211_X1 g090(.A(new_n280), .B(new_n284), .C1(new_n289), .C2(new_n291), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n271), .A2(new_n279), .B1(new_n292), .B2(KEYINPUT25), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT64), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n278), .B1(new_n294), .B2(KEYINPUT24), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n286), .A2(KEYINPUT64), .A3(G183gat), .A4(G190gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI22_X1  g096(.A1(new_n266), .A2(new_n264), .B1(new_n294), .B2(KEYINPUT24), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT65), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT65), .ZN(new_n301));
  NOR3_X1   g100(.A1(new_n278), .A2(new_n294), .A3(KEYINPUT24), .ZN(new_n302));
  AOI22_X1  g101(.A1(new_n286), .A2(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n301), .B(new_n298), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT25), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n283), .B1(G169gat), .B2(G176gat), .ZN(new_n306));
  AND4_X1   g105(.A1(new_n305), .A2(new_n280), .A3(new_n306), .A4(new_n275), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n300), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G226gat), .A2(G233gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G197gat), .B(G204gat), .ZN(new_n313));
  INV_X1    g112(.A(G211gat), .ZN(new_n314));
  INV_X1    g113(.A(G218gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n313), .B1(KEYINPUT22), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G211gat), .B(G218gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n312), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT29), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n292), .A2(KEYINPUT25), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n267), .A2(new_n269), .A3(new_n264), .ZN(new_n325));
  INV_X1    g124(.A(new_n262), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n262), .A2(new_n267), .A3(new_n269), .A4(new_n264), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n327), .A2(new_n277), .A3(new_n278), .A4(new_n328), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n308), .A2(KEYINPUT75), .A3(new_n324), .A4(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT75), .B1(new_n293), .B2(new_n308), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n323), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT76), .B1(new_n333), .B2(new_n310), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT75), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n280), .A2(new_n306), .A3(new_n275), .ZN(new_n336));
  INV_X1    g135(.A(new_n291), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n290), .A2(new_n286), .B1(new_n266), .B2(new_n264), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n329), .B1(new_n339), .B2(new_n305), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n304), .A2(new_n307), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n301), .B1(new_n297), .B2(new_n298), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n335), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT29), .B1(new_n344), .B2(new_n330), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT76), .ZN(new_n346));
  NOR3_X1   g145(.A1(new_n345), .A2(new_n346), .A3(new_n311), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n322), .B1(new_n334), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n344), .A2(new_n311), .A3(new_n330), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n309), .A2(new_n323), .A3(new_n310), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n349), .A2(new_n319), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G64gat), .B(G92gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(G8gat), .B(G36gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n355), .B(new_n356), .Z(new_n357));
  NAND4_X1  g156(.A1(new_n348), .A2(KEYINPUT30), .A3(new_n352), .A4(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n357), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n333), .A2(KEYINPUT76), .A3(new_n310), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n346), .B1(new_n345), .B2(new_n311), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n321), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n359), .B1(new_n362), .B2(new_n351), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n360), .A2(new_n361), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n351), .B1(new_n365), .B2(new_n322), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT30), .B1(new_n366), .B2(new_n357), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n260), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n348), .A2(new_n352), .A3(new_n357), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT30), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n371), .A2(KEYINPUT85), .A3(new_n358), .A4(new_n363), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n368), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G1gat), .B(G29gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n374), .B(KEYINPUT0), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(G57gat), .ZN(new_n376));
  INV_X1    g175(.A(G85gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT3), .ZN(new_n380));
  NAND2_X1  g179(.A1(G155gat), .A2(G162gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT2), .ZN(new_n382));
  INV_X1    g181(.A(G141gat), .ZN(new_n383));
  INV_X1    g182(.A(G148gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G141gat), .A2(G148gat), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n382), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT79), .ZN(new_n388));
  XNOR2_X1  g187(.A(G155gat), .B(G162gat), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n389), .B1(new_n387), .B2(new_n388), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n380), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n387), .A2(new_n388), .ZN(new_n393));
  INV_X1    g192(.A(new_n389), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(KEYINPUT3), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT1), .ZN(new_n398));
  INV_X1    g197(.A(G120gat), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n399), .A2(G113gat), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(G113gat), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n398), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G134gat), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n403), .A2(G127gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(G127gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  AND2_X1   g206(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(KEYINPUT68), .A2(G113gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n400), .B1(new_n410), .B2(G120gat), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n404), .A2(new_n398), .A3(new_n405), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n407), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n392), .A2(new_n397), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n396), .ZN(new_n415));
  INV_X1    g214(.A(new_n412), .ZN(new_n416));
  INV_X1    g215(.A(new_n400), .ZN(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT68), .B(G113gat), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n417), .B1(new_n418), .B2(new_n399), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n416), .A2(new_n419), .B1(new_n402), .B2(new_n406), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n415), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n390), .A2(new_n391), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT80), .B1(new_n423), .B2(new_n413), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT80), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n415), .A2(new_n420), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n421), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT82), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n422), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI211_X1 g228(.A(KEYINPUT82), .B(new_n421), .C1(new_n424), .C2(new_n426), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n414), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G225gat), .A2(G233gat), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT39), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n433), .B1(new_n424), .B2(new_n426), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT81), .B1(new_n415), .B2(new_n420), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT81), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n423), .A2(new_n438), .A3(new_n413), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n435), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n379), .B1(new_n434), .B2(new_n441), .ZN(new_n442));
  XOR2_X1   g241(.A(KEYINPUT86), .B(KEYINPUT39), .Z(new_n443));
  NAND3_X1  g242(.A1(new_n431), .A2(new_n433), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT87), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT40), .ZN(new_n446));
  OR2_X1    g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n433), .A2(KEYINPUT5), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n414), .B(new_n448), .C1(new_n429), .C2(new_n430), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n437), .A2(new_n439), .A3(new_n433), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n424), .A2(new_n426), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n432), .A2(KEYINPUT4), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n415), .A2(KEYINPUT4), .A3(new_n420), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n433), .B1(new_n414), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(KEYINPUT5), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n378), .B1(new_n449), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n457), .B1(new_n445), .B2(new_n446), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n373), .A2(new_n447), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n348), .A2(new_n352), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n357), .B1(new_n460), .B2(KEYINPUT37), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT37), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT88), .B1(new_n366), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT88), .ZN(new_n464));
  NOR4_X1   g263(.A1(new_n362), .A2(new_n464), .A3(KEYINPUT37), .A4(new_n351), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n461), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT38), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n449), .A2(new_n456), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n379), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT6), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n449), .A2(new_n456), .A3(new_n378), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n468), .A2(KEYINPUT6), .A3(new_n379), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT89), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT89), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n457), .A2(new_n475), .A3(KEYINPUT6), .ZN(new_n476));
  AND4_X1   g275(.A1(new_n472), .A2(new_n474), .A3(new_n369), .A4(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n365), .A2(new_n319), .A3(new_n312), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n349), .A2(new_n350), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n462), .B1(new_n479), .B2(new_n320), .ZN(new_n480));
  AOI211_X1 g279(.A(KEYINPUT38), .B(new_n357), .C1(new_n478), .C2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n481), .B1(new_n463), .B2(new_n465), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n467), .A2(new_n477), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(G22gat), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n380), .B1(new_n319), .B2(KEYINPUT29), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n485), .A2(new_n423), .ZN(new_n486));
  INV_X1    g285(.A(new_n392), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n319), .B1(new_n487), .B2(KEYINPUT29), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G228gat), .A2(G233gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n486), .A2(new_n488), .A3(G228gat), .A4(G233gat), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n484), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n491), .A2(new_n484), .A3(new_n492), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(KEYINPUT83), .A3(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G78gat), .B(G106gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(KEYINPUT31), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(G50gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT83), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n499), .B1(new_n493), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n494), .A2(new_n495), .A3(new_n499), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT84), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n494), .A2(KEYINPUT84), .A3(new_n495), .A4(new_n499), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n502), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n459), .A2(new_n483), .A3(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n420), .B1(new_n340), .B2(new_n343), .ZN(new_n509));
  NAND2_X1  g308(.A1(G227gat), .A2(G233gat), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n308), .A2(new_n413), .A3(new_n324), .A4(new_n329), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n509), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT32), .ZN(new_n514));
  INV_X1    g313(.A(G43gat), .ZN(new_n515));
  INV_X1    g314(.A(G99gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(G71gat), .ZN(new_n517));
  INV_X1    g316(.A(G71gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(G99gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT69), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n517), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n520), .B1(new_n517), .B2(new_n519), .ZN(new_n523));
  NOR3_X1   g322(.A1(new_n522), .A2(new_n523), .A3(G15gat), .ZN(new_n524));
  INV_X1    g323(.A(G15gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n517), .A2(new_n519), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT69), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n525), .B1(new_n527), .B2(new_n521), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n515), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(G15gat), .B1(new_n522), .B2(new_n523), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n527), .A2(new_n525), .A3(new_n521), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(new_n531), .A3(G43gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n514), .B1(new_n533), .B2(KEYINPUT33), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n513), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT70), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT70), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n513), .A2(new_n534), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n514), .A2(KEYINPUT33), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n513), .A2(new_n539), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n536), .A2(new_n538), .B1(new_n540), .B2(new_n533), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n509), .A2(new_n512), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n510), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT34), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n544), .B1(new_n510), .B2(KEYINPUT71), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n542), .B(new_n510), .C1(KEYINPUT71), .C2(new_n544), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n541), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT73), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT72), .B1(new_n541), .B2(new_n549), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n540), .A2(new_n533), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n513), .A2(new_n534), .A3(new_n537), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n537), .B1(new_n513), .B2(new_n534), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT72), .ZN(new_n557));
  NOR3_X1   g356(.A1(new_n556), .A2(new_n548), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n551), .B1(new_n552), .B2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n541), .A2(new_n549), .A3(KEYINPUT72), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n557), .B1(new_n556), .B2(new_n548), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(new_n561), .A3(KEYINPUT73), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n550), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(KEYINPUT74), .B1(new_n563), .B2(KEYINPUT36), .ZN(new_n564));
  INV_X1    g363(.A(new_n550), .ZN(new_n565));
  AND3_X1   g364(.A1(new_n560), .A2(new_n561), .A3(KEYINPUT73), .ZN(new_n566));
  AOI21_X1  g365(.A(KEYINPUT73), .B1(new_n560), .B2(new_n561), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT74), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT36), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n550), .B1(new_n561), .B2(new_n560), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT36), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n564), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n502), .A2(new_n505), .A3(new_n506), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n472), .A2(new_n473), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n371), .A2(new_n358), .A3(new_n363), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n508), .A2(new_n574), .A3(new_n579), .ZN(new_n580));
  XOR2_X1   g379(.A(KEYINPUT90), .B(KEYINPUT35), .Z(new_n581));
  NOR2_X1   g380(.A1(new_n575), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n472), .A2(new_n474), .A3(new_n476), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n582), .A2(new_n583), .A3(new_n368), .A4(new_n372), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n507), .A2(new_n572), .ZN(new_n585));
  NOR3_X1   g384(.A1(new_n585), .A2(new_n577), .A3(new_n578), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT35), .ZN(new_n587));
  OAI22_X1  g386(.A1(new_n584), .A2(new_n568), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n259), .B1(new_n580), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT21), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT9), .ZN(new_n591));
  XNOR2_X1  g390(.A(G57gat), .B(G64gat), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n591), .B1(new_n592), .B2(KEYINPUT97), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n593), .B1(KEYINPUT97), .B2(new_n592), .ZN(new_n594));
  NAND2_X1  g393(.A1(G71gat), .A2(G78gat), .ZN(new_n595));
  NOR2_X1   g394(.A1(G71gat), .A2(G78gat), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT96), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n598), .B1(new_n597), .B2(new_n596), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n596), .A2(KEYINPUT9), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n601), .A2(new_n595), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n602), .A2(new_n592), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n216), .B1(new_n590), .B2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(G183gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n590), .ZN(new_n607));
  XNOR2_X1  g406(.A(G127gat), .B(G155gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n606), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT98), .ZN(new_n612));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(KEYINPUT99), .B(G211gat), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n610), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G190gat), .B(G218gat), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT101), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(KEYINPUT100), .A2(G85gat), .A3(G92gat), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT7), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g426(.A1(G99gat), .A2(G106gat), .ZN(new_n628));
  INV_X1    g427(.A(G92gat), .ZN(new_n629));
  AOI22_X1  g428(.A1(KEYINPUT8), .A2(new_n628), .B1(new_n377), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n626), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G99gat), .B(G106gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT41), .ZN(new_n635));
  AND2_X1   g434(.A1(G232gat), .A2(G233gat), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  OAI22_X1  g436(.A1(new_n229), .A2(new_n634), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n232), .A2(new_n233), .A3(new_n634), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n623), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G134gat), .B(G162gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n621), .A2(new_n622), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n637), .A2(new_n635), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n643), .A2(new_n646), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(G230gat), .ZN(new_n651));
  INV_X1    g450(.A(G233gat), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n600), .A2(new_n603), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n633), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT10), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n634), .A2(new_n604), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n654), .A2(KEYINPUT10), .A3(new_n633), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n653), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n655), .A2(new_n657), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n660), .B1(new_n661), .B2(new_n653), .ZN(new_n662));
  XNOR2_X1  g461(.A(G120gat), .B(G148gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT103), .B(G204gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT102), .B(G176gat), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n665), .B(new_n666), .Z(new_n667));
  OR2_X1    g466(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n660), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n661), .A2(new_n653), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(new_n670), .A3(new_n667), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n620), .A2(new_n650), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n589), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n576), .B(KEYINPUT104), .Z(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(G1gat), .Z(G1324gat));
  INV_X1    g477(.A(new_n373), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n674), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT16), .B(G8gat), .Z(new_n681));
  AND2_X1   g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(KEYINPUT42), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(KEYINPUT42), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n683), .B(new_n684), .C1(new_n212), .C2(new_n680), .ZN(G1325gat));
  OAI21_X1  g484(.A(G15gat), .B1(new_n674), .B2(new_n574), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n563), .A2(new_n525), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n686), .B1(new_n674), .B2(new_n687), .ZN(G1326gat));
  NOR2_X1   g487(.A1(new_n674), .A2(new_n507), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT43), .B(G22gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT105), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n689), .B(new_n691), .ZN(G1327gat));
  NOR3_X1   g491(.A1(new_n619), .A2(new_n649), .A3(new_n672), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n589), .A2(new_n220), .A3(new_n675), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT45), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n580), .A2(new_n588), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n696), .B1(new_n697), .B2(new_n650), .ZN(new_n698));
  AOI211_X1 g497(.A(KEYINPUT44), .B(new_n649), .C1(new_n580), .C2(new_n588), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n619), .B(KEYINPUT106), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n701), .A2(new_n259), .A3(new_n672), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(new_n676), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n695), .B1(new_n704), .B2(new_n220), .ZN(G1328gat));
  NAND4_X1  g504(.A1(new_n589), .A2(new_n221), .A3(new_n373), .A4(new_n693), .ZN(new_n706));
  AND2_X1   g505(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n707));
  NOR2_X1   g506(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n710), .B1(new_n703), .B2(new_n679), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(G36gat), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n703), .A2(new_n710), .A3(new_n679), .ZN(new_n713));
  OAI221_X1 g512(.A(new_n709), .B1(new_n707), .B2(new_n706), .C1(new_n712), .C2(new_n713), .ZN(G1329gat));
  INV_X1    g513(.A(KEYINPUT47), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(KEYINPUT109), .ZN(new_n716));
  OAI21_X1  g515(.A(G43gat), .B1(new_n703), .B2(new_n574), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n589), .A2(new_n515), .A3(new_n563), .A4(new_n693), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n715), .A2(KEYINPUT109), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n719), .B(new_n720), .ZN(G1330gat));
  OAI21_X1  g520(.A(G50gat), .B1(new_n703), .B2(new_n507), .ZN(new_n722));
  INV_X1    g521(.A(G50gat), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n589), .A2(new_n723), .A3(new_n575), .A4(new_n693), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(KEYINPUT48), .Z(G1331gat));
  NAND3_X1  g525(.A1(new_n259), .A2(new_n619), .A3(new_n649), .ZN(new_n727));
  INV_X1    g526(.A(new_n672), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT110), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n730), .B1(new_n580), .B2(new_n588), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n675), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g532(.A1(new_n731), .A2(new_n373), .ZN(new_n734));
  NOR2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  AND2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n734), .B2(new_n735), .ZN(G1333gat));
  INV_X1    g537(.A(new_n574), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n518), .B1(new_n731), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n568), .A2(G71gat), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n740), .B1(new_n731), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g542(.A1(new_n731), .A2(new_n575), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G78gat), .ZN(G1335gat));
  AOI21_X1  g544(.A(new_n649), .B1(new_n580), .B2(new_n588), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n619), .A2(new_n258), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n746), .A2(KEYINPUT51), .A3(new_n747), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n728), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n752), .A2(new_n377), .A3(new_n675), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n619), .A2(new_n258), .A3(new_n728), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n698), .B2(new_n699), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT111), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI211_X1 g556(.A(KEYINPUT111), .B(new_n754), .C1(new_n698), .C2(new_n699), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n757), .A2(new_n675), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n753), .B1(new_n759), .B2(new_n377), .ZN(G1336gat));
  AND3_X1   g559(.A1(new_n752), .A2(new_n629), .A3(new_n373), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(KEYINPUT52), .ZN(new_n762));
  OAI21_X1  g561(.A(G92gat), .B1(new_n755), .B2(new_n679), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n757), .A2(new_n373), .A3(new_n758), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n765), .A2(new_n766), .A3(G92gat), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n766), .B1(new_n765), .B2(G92gat), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n767), .A2(new_n768), .A3(new_n761), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n764), .B1(new_n769), .B2(new_n770), .ZN(G1337gat));
  NAND2_X1  g570(.A1(new_n750), .A2(new_n751), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n568), .A2(G99gat), .A3(new_n728), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT113), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n757), .A2(new_n739), .A3(new_n758), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n775), .B1(new_n776), .B2(new_n516), .ZN(G1338gat));
  NOR2_X1   g576(.A1(new_n507), .A2(G106gat), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT53), .B1(new_n752), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n780));
  XOR2_X1   g579(.A(KEYINPUT114), .B(G106gat), .Z(new_n781));
  OAI21_X1  g580(.A(new_n781), .B1(new_n755), .B2(new_n507), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n779), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n780), .B1(new_n779), .B2(new_n782), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n757), .A2(new_n575), .A3(new_n758), .ZN(new_n785));
  AOI22_X1  g584(.A1(new_n785), .A2(new_n781), .B1(new_n752), .B2(new_n778), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787));
  OAI22_X1  g586(.A1(new_n783), .A2(new_n784), .B1(new_n786), .B2(new_n787), .ZN(G1339gat));
  NOR2_X1   g587(.A1(new_n727), .A2(new_n672), .ZN(new_n789));
  INV_X1    g588(.A(new_n207), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n236), .B1(new_n235), .B2(new_n238), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n240), .A2(new_n241), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n254), .A2(new_n672), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n658), .A2(new_n659), .A3(new_n653), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n669), .A2(KEYINPUT54), .A3(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n667), .B1(new_n660), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(KEYINPUT55), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n671), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT55), .B1(new_n798), .B2(new_n800), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n258), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n254), .A2(new_n672), .A3(KEYINPUT116), .A4(new_n793), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n796), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n649), .ZN(new_n808));
  INV_X1    g607(.A(new_n804), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(new_n649), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n254), .A2(new_n793), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n701), .B1(new_n813), .B2(KEYINPUT117), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n808), .A2(new_n815), .A3(new_n812), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n789), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n676), .A2(new_n373), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n817), .A2(new_n575), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n563), .ZN(new_n821));
  OAI21_X1  g620(.A(G113gat), .B1(new_n821), .B2(new_n259), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n820), .A2(new_n572), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n258), .A2(new_n410), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(KEYINPUT118), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n822), .B1(new_n823), .B2(new_n825), .ZN(G1340gat));
  OAI21_X1  g625(.A(G120gat), .B1(new_n821), .B2(new_n728), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n672), .A2(new_n399), .ZN(new_n828));
  XOR2_X1   g627(.A(new_n828), .B(KEYINPUT119), .Z(new_n829));
  OAI21_X1  g628(.A(new_n827), .B1(new_n823), .B2(new_n829), .ZN(G1341gat));
  INV_X1    g629(.A(new_n701), .ZN(new_n831));
  OAI21_X1  g630(.A(G127gat), .B1(new_n821), .B2(new_n831), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n620), .A2(G127gat), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n823), .B2(new_n833), .ZN(G1342gat));
  NAND2_X1  g633(.A1(new_n650), .A2(new_n403), .ZN(new_n835));
  OR3_X1    g634(.A1(new_n823), .A2(KEYINPUT56), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(G134gat), .B1(new_n821), .B2(new_n649), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT56), .B1(new_n823), .B2(new_n835), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(G1343gat));
  NOR3_X1   g638(.A1(new_n817), .A2(KEYINPUT57), .A3(new_n507), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n805), .A2(new_n794), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n649), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n812), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n789), .B1(new_n843), .B2(new_n620), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT57), .B1(new_n844), .B2(new_n507), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n819), .A2(new_n739), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n840), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(G141gat), .B1(new_n849), .B2(new_n259), .ZN(new_n850));
  AOI22_X1  g649(.A1(new_n795), .A2(new_n794), .B1(new_n258), .B2(new_n804), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n650), .B1(new_n851), .B2(new_n806), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n810), .A2(new_n811), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT117), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n831), .A3(new_n816), .ZN(new_n855));
  INV_X1    g654(.A(new_n789), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n507), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n846), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n383), .A3(new_n258), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n850), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT58), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT58), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n850), .A2(new_n863), .A3(new_n860), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(G1344gat));
  NAND3_X1  g664(.A1(new_n859), .A2(new_n384), .A3(new_n672), .ZN(new_n866));
  AOI211_X1 g665(.A(KEYINPUT59), .B(new_n384), .C1(new_n848), .C2(new_n672), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868));
  OAI21_X1  g667(.A(KEYINPUT57), .B1(new_n817), .B2(new_n507), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT57), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n810), .A2(KEYINPUT120), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n810), .A2(KEYINPUT120), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n811), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n619), .B1(new_n873), .B2(new_n842), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n870), .B(new_n575), .C1(new_n874), .C2(new_n789), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n869), .A2(new_n672), .A3(new_n846), .A4(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n868), .B1(new_n876), .B2(G148gat), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n866), .B1(new_n867), .B2(new_n877), .ZN(G1345gat));
  OAI21_X1  g677(.A(G155gat), .B1(new_n849), .B2(new_n831), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n620), .A2(G155gat), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n879), .B1(new_n858), .B2(new_n880), .ZN(G1346gat));
  OAI21_X1  g680(.A(G162gat), .B1(new_n849), .B2(new_n649), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n649), .A2(G162gat), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n858), .B2(new_n883), .ZN(G1347gat));
  NOR2_X1   g683(.A1(new_n675), .A2(new_n679), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n817), .A2(new_n585), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(G169gat), .B1(new_n887), .B2(new_n258), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n817), .A2(new_n575), .ZN(new_n889));
  XNOR2_X1  g688(.A(new_n886), .B(KEYINPUT121), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(new_n568), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n259), .A2(new_n204), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n888), .B1(new_n893), .B2(new_n894), .ZN(G1348gat));
  OAI21_X1  g694(.A(G176gat), .B1(new_n892), .B2(new_n728), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n887), .A2(new_n273), .A3(new_n672), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1349gat));
  OAI21_X1  g697(.A(G183gat), .B1(new_n892), .B2(new_n831), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT123), .B1(KEYINPUT122), .B2(KEYINPUT60), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n887), .A2(new_n263), .A3(new_n619), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n899), .A2(new_n901), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n903), .B1(KEYINPUT123), .B2(KEYINPUT60), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n902), .B1(new_n904), .B2(new_n900), .ZN(G1350gat));
  AOI21_X1  g704(.A(new_n264), .B1(new_n893), .B2(new_n650), .ZN(new_n906));
  OR2_X1    g705(.A1(new_n906), .A2(KEYINPUT61), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n887), .A2(new_n264), .A3(new_n650), .ZN(new_n908));
  XOR2_X1   g707(.A(new_n908), .B(KEYINPUT124), .Z(new_n909));
  NAND2_X1  g708(.A1(new_n906), .A2(KEYINPUT61), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n907), .A2(new_n909), .A3(new_n910), .ZN(G1351gat));
  NOR2_X1   g710(.A1(new_n886), .A2(new_n739), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n857), .A2(new_n912), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n913), .A2(G197gat), .A3(new_n259), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT125), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n890), .A2(new_n739), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n916), .B(new_n875), .C1(new_n870), .C2(new_n857), .ZN(new_n917));
  OAI21_X1  g716(.A(G197gat), .B1(new_n917), .B2(new_n259), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n915), .A2(new_n918), .ZN(G1352gat));
  NOR2_X1   g718(.A1(new_n728), .A2(G204gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n857), .A2(new_n912), .A3(new_n920), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT126), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n869), .A2(new_n672), .A3(new_n875), .ZN(new_n926));
  INV_X1    g725(.A(new_n916), .ZN(new_n927));
  OAI21_X1  g726(.A(G204gat), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n924), .A2(new_n925), .A3(new_n928), .ZN(G1353gat));
  NAND4_X1  g728(.A1(new_n857), .A2(new_n314), .A3(new_n619), .A4(new_n912), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n869), .A2(new_n619), .A3(new_n875), .A4(new_n916), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT63), .B1(new_n931), .B2(G211gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT127), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT127), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n937), .B(new_n930), .C1(new_n933), .C2(new_n934), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1354gat));
  OAI21_X1  g738(.A(new_n315), .B1(new_n913), .B2(new_n649), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n650), .A2(G218gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n917), .B2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(G1355gat));
endmodule


