//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1185, new_n1186, new_n1187, new_n1188, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1241, new_n1242, new_n1243;
  OR3_X1    g0000(.A1(KEYINPUT64), .A2(G58), .A3(G68), .ZN(new_n201));
  OAI21_X1  g0001(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(G50), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G77), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT65), .Z(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NOR2_X1   g0008(.A1(new_n203), .A2(new_n204), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n213), .B1(new_n214), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n219), .B(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT66), .Z(new_n225));
  AOI211_X1 g0025(.A(new_n223), .B(new_n225), .C1(G77), .C2(G244), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(G1), .B2(G20), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT1), .Z(new_n228));
  AOI211_X1 g0028(.A(new_n218), .B(new_n228), .C1(new_n214), .C2(new_n217), .ZN(G361));
  XOR2_X1   g0029(.A(G226), .B(G232), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  INV_X1    g0045(.A(KEYINPUT10), .ZN(new_n246));
  OR2_X1    g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G1698), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G222), .ZN(new_n251));
  INV_X1    g0051(.A(G223), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n249), .B(new_n251), .C1(new_n252), .C2(new_n250), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  OAI211_X1 g0055(.A(G1), .B(G13), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n253), .B(new_n257), .C1(G77), .C2(new_n249), .ZN(new_n258));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G226), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  OR2_X1    g0064(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n258), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  OR2_X1    g0066(.A1(new_n266), .A2(KEYINPUT68), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(KEYINPUT68), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G200), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT73), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n267), .A2(new_n268), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n271), .B1(new_n272), .B2(G190), .ZN(new_n273));
  INV_X1    g0073(.A(G190), .ZN(new_n274));
  AOI211_X1 g0074(.A(KEYINPUT73), .B(new_n274), .C1(new_n267), .C2(new_n268), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n270), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n205), .A2(G20), .ZN(new_n277));
  INV_X1    g0077(.A(G150), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G20), .A2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT8), .B(G58), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT70), .ZN(new_n282));
  XNOR2_X1  g0082(.A(new_n281), .B(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n211), .A2(G33), .ZN(new_n284));
  OAI221_X1 g0084(.A(new_n277), .B1(new_n278), .B2(new_n280), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n210), .B1(new_n215), .B2(new_n254), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT69), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(KEYINPUT69), .B(new_n210), .C1(new_n215), .C2(new_n254), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n285), .A2(new_n290), .B1(new_n204), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n290), .B1(new_n259), .B2(G20), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G50), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT9), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT9), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n293), .A2(new_n298), .A3(new_n295), .ZN(new_n299));
  AND2_X1   g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n246), .B1(new_n276), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT73), .B1(new_n269), .B2(new_n274), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n272), .A2(new_n271), .A3(G190), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n297), .A2(new_n299), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n304), .A2(KEYINPUT10), .A3(new_n270), .A4(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n269), .A2(G179), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n296), .B1(new_n272), .B2(G169), .ZN(new_n308));
  OR2_X1    g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT72), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n294), .A2(G77), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT71), .ZN(new_n312));
  INV_X1    g0112(.A(G77), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n292), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT71), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n294), .A2(new_n315), .A3(G77), .ZN(new_n316));
  XOR2_X1   g0116(.A(KEYINPUT15), .B(G87), .Z(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n280), .A2(new_n281), .B1(new_n318), .B2(new_n284), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n211), .A2(new_n313), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n290), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n312), .A2(new_n314), .A3(new_n316), .A4(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n250), .A2(G232), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n249), .B(new_n323), .C1(new_n222), .C2(new_n250), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n324), .B(new_n257), .C1(G107), .C2(new_n249), .ZN(new_n325));
  INV_X1    g0125(.A(G244), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n325), .B(new_n265), .C1(new_n326), .C2(new_n261), .ZN(new_n327));
  AND2_X1   g0127(.A1(new_n327), .A2(G200), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n327), .A2(new_n274), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  OR2_X1    g0131(.A1(new_n327), .A2(G179), .ZN(new_n332));
  INV_X1    g0132(.A(G169), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n322), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n310), .B1(new_n331), .B2(new_n336), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n301), .A2(new_n306), .A3(new_n309), .A4(new_n337), .ZN(new_n338));
  AND2_X1   g0138(.A1(KEYINPUT3), .A2(G33), .ZN(new_n339));
  NOR2_X1   g0139(.A1(KEYINPUT3), .A2(G33), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT7), .B1(new_n341), .B2(new_n211), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT7), .ZN(new_n343));
  NOR4_X1   g0143(.A1(new_n339), .A2(new_n340), .A3(new_n343), .A4(G20), .ZN(new_n344));
  OAI21_X1  g0144(.A(G68), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n279), .A2(G159), .ZN(new_n346));
  INV_X1    g0146(.A(G58), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n347), .A2(new_n221), .ZN(new_n348));
  OAI21_X1  g0148(.A(G20), .B1(new_n203), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n345), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT16), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n345), .A2(KEYINPUT16), .A3(new_n346), .A4(new_n349), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(new_n290), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n283), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n355), .A2(new_n291), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n356), .B1(new_n355), .B2(new_n294), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n256), .A2(G232), .A3(new_n260), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n265), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(G190), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n252), .A2(new_n250), .ZN(new_n361));
  INV_X1    g0161(.A(G226), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G1698), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n361), .B(new_n363), .C1(new_n339), .C2(new_n340), .ZN(new_n364));
  NAND2_X1  g0164(.A1(G33), .A2(G87), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n256), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT74), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI211_X1 g0168(.A(KEYINPUT74), .B(new_n256), .C1(new_n364), .C2(new_n365), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n360), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G200), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n366), .B2(new_n359), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n354), .A2(new_n357), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT17), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n354), .A2(new_n357), .A3(KEYINPUT17), .A4(new_n373), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT18), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n354), .A2(new_n357), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n359), .A2(G179), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n381), .B1(new_n368), .B2(new_n369), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n333), .B1(new_n366), .B2(new_n359), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n379), .B1(new_n380), .B2(new_n385), .ZN(new_n386));
  AOI211_X1 g0186(.A(KEYINPUT18), .B(new_n384), .C1(new_n354), .C2(new_n357), .ZN(new_n387));
  NOR3_X1   g0187(.A1(new_n378), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n362), .A2(new_n250), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n249), .B(new_n389), .C1(G232), .C2(new_n250), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G33), .A2(G97), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n256), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n265), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n261), .A2(new_n222), .ZN(new_n394));
  NOR3_X1   g0194(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT13), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NOR4_X1   g0197(.A1(new_n392), .A2(KEYINPUT13), .A3(new_n393), .A4(new_n394), .ZN(new_n398));
  OAI21_X1  g0198(.A(G169), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT14), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n397), .A2(new_n398), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G179), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT14), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n403), .B(G169), .C1(new_n397), .C2(new_n398), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n400), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n284), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n406), .A2(G77), .B1(new_n279), .B2(G50), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n211), .B2(G68), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n290), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT11), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n294), .A2(G68), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n408), .A2(KEYINPUT11), .A3(new_n290), .ZN(new_n413));
  INV_X1    g0213(.A(G13), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n414), .A2(G1), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n415), .A2(G20), .A3(new_n221), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT12), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n411), .A2(new_n412), .A3(new_n413), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n405), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n418), .B1(new_n401), .B2(G190), .ZN(new_n420));
  OAI21_X1  g0220(.A(G200), .B1(new_n397), .B2(new_n398), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(KEYINPUT72), .B(new_n335), .C1(new_n329), .C2(new_n330), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n388), .A2(new_n419), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n338), .A2(new_n424), .ZN(new_n425));
  AOI22_X1  g0225(.A1(new_n415), .A2(G20), .B1(new_n259), .B2(G33), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n288), .A2(new_n426), .A3(new_n289), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT76), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n288), .A2(new_n426), .A3(KEYINPUT76), .A4(new_n289), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(G107), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(G107), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n415), .A2(G20), .A3(new_n432), .ZN(new_n433));
  OR2_X1    g0233(.A1(new_n433), .A2(KEYINPUT25), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n432), .A2(G20), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT23), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n211), .B(G87), .C1(new_n339), .C2(new_n340), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT22), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT22), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n249), .A2(new_n440), .A3(new_n211), .A4(G87), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n437), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n406), .A2(G116), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n442), .A2(KEYINPUT24), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT24), .B1(new_n442), .B2(new_n443), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n435), .B1(new_n446), .B2(new_n290), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n433), .A2(KEYINPUT25), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT77), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT5), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n449), .B1(new_n450), .B2(G41), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n255), .A2(KEYINPUT77), .A3(KEYINPUT5), .ZN(new_n452));
  INV_X1    g0252(.A(G45), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(G1), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n450), .A2(G41), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n451), .A2(new_n452), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n456), .A2(G264), .A3(new_n256), .ZN(new_n457));
  INV_X1    g0257(.A(G257), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(G1698), .ZN(new_n459));
  OAI221_X1 g0259(.A(new_n459), .B1(G250), .B2(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G294), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n256), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  OR2_X1    g0263(.A1(new_n456), .A2(new_n264), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G190), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(G200), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n447), .A2(new_n448), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n442), .A2(new_n443), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT24), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n442), .A2(KEYINPUT24), .A3(new_n443), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(new_n290), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n435), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n474), .A2(new_n448), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n465), .A2(new_n333), .ZN(new_n477));
  INV_X1    g0277(.A(G179), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n466), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n476), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n291), .A2(G116), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT80), .ZN(new_n482));
  XNOR2_X1  g0282(.A(new_n481), .B(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n288), .A2(new_n426), .A3(G116), .A4(new_n289), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G283), .ZN(new_n485));
  INV_X1    g0285(.A(G97), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n485), .B(new_n211), .C1(G33), .C2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(G116), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G20), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n286), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT20), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n490), .A2(new_n491), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n483), .B(new_n484), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G264), .A2(G1698), .ZN(new_n495));
  OAI221_X1 g0295(.A(new_n495), .B1(new_n458), .B2(G1698), .C1(new_n339), .C2(new_n340), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n496), .B(new_n257), .C1(G303), .C2(new_n249), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n456), .A2(G270), .A3(new_n256), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n497), .A2(new_n464), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n494), .A2(G169), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT21), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n499), .A2(new_n478), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n494), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n494), .A2(KEYINPUT21), .A3(G169), .A4(new_n499), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n502), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n469), .A2(new_n480), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n290), .ZN(new_n508));
  OR2_X1    g0308(.A1(KEYINPUT6), .A2(G97), .ZN(new_n509));
  OAI21_X1  g0309(.A(KEYINPUT6), .B1(G97), .B2(G107), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT75), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n511), .B1(new_n509), .B2(new_n510), .ZN(new_n514));
  NOR3_X1   g0314(.A1(new_n513), .A2(new_n514), .A3(new_n432), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n509), .A2(new_n510), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT75), .ZN(new_n517));
  AOI21_X1  g0317(.A(G107), .B1(new_n517), .B2(new_n512), .ZN(new_n518));
  OAI21_X1  g0318(.A(G20), .B1(new_n515), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n343), .B1(new_n249), .B2(G20), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n341), .A2(KEYINPUT7), .A3(new_n211), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n522), .A2(G107), .B1(G77), .B2(new_n279), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n508), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n429), .A2(G97), .A3(new_n430), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n292), .A2(new_n486), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(KEYINPUT78), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  AND2_X1   g0328(.A1(new_n525), .A2(new_n526), .ZN(new_n529));
  OAI21_X1  g0329(.A(G107), .B1(new_n342), .B2(new_n344), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n313), .B2(new_n280), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n432), .B1(new_n513), .B2(new_n514), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n517), .A2(G107), .A3(new_n512), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n211), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n290), .B1(new_n531), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT78), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n529), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n528), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT4), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(G1698), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n540), .B(G244), .C1(new_n340), .C2(new_n339), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n326), .B1(new_n247), .B2(new_n248), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n541), .B(new_n485), .C1(new_n542), .C2(KEYINPUT4), .ZN(new_n543));
  OAI21_X1  g0343(.A(G250), .B1(new_n339), .B2(new_n340), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n250), .B1(new_n544), .B2(KEYINPUT4), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n257), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n456), .A2(G257), .A3(new_n256), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n546), .A2(new_n464), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G179), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n546), .A2(new_n464), .A3(new_n547), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(G169), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n538), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n550), .A2(G200), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n546), .A2(G190), .A3(new_n464), .A4(new_n547), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n529), .A2(new_n535), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT19), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n284), .B2(new_n486), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT79), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n249), .A2(new_n211), .A3(G68), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n211), .B1(new_n391), .B2(new_n560), .ZN(new_n564));
  INV_X1    g0364(.A(G87), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n565), .A2(new_n486), .A3(new_n432), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT79), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n568), .B(new_n560), .C1(new_n284), .C2(new_n486), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n562), .A2(new_n563), .A3(new_n567), .A4(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n570), .A2(new_n290), .B1(new_n292), .B2(new_n318), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n429), .A2(G87), .A3(new_n430), .ZN(new_n572));
  AND2_X1   g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n222), .A2(new_n250), .ZN(new_n574));
  OAI221_X1 g0374(.A(new_n574), .B1(G244), .B2(new_n250), .C1(new_n339), .C2(new_n340), .ZN(new_n575));
  NAND2_X1  g0375(.A1(G33), .A2(G116), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n256), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n454), .A2(new_n264), .ZN(new_n578));
  INV_X1    g0378(.A(G250), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n453), .B2(G1), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n256), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n577), .A2(new_n274), .A3(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n247), .A2(new_n248), .B1(new_n326), .B2(G1698), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n584), .A2(new_n574), .B1(G33), .B2(G116), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n581), .B1(new_n585), .B2(new_n256), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n583), .B1(G200), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n429), .A2(new_n317), .A3(new_n430), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n571), .A2(new_n588), .B1(new_n333), .B2(new_n586), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n577), .A2(new_n582), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n478), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n573), .A2(new_n587), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  AND3_X1   g0392(.A1(new_n553), .A2(new_n559), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n494), .B1(G200), .B2(new_n499), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n274), .B2(new_n499), .ZN(new_n595));
  AND4_X1   g0395(.A1(new_n425), .A2(new_n507), .A3(new_n593), .A4(new_n595), .ZN(G372));
  NAND2_X1  g0396(.A1(new_n480), .A2(new_n506), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n538), .A2(new_n552), .B1(new_n558), .B2(new_n556), .ZN(new_n598));
  AND4_X1   g0398(.A1(new_n597), .A2(new_n598), .A3(new_n469), .A4(new_n592), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n538), .A2(new_n592), .A3(new_n552), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT26), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n571), .A2(new_n588), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n586), .A2(new_n333), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n602), .A2(new_n603), .A3(new_n591), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT26), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n592), .A2(new_n552), .A3(new_n605), .A4(new_n557), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n601), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n425), .B1(new_n599), .B2(new_n607), .ZN(new_n608));
  XOR2_X1   g0408(.A(new_n608), .B(KEYINPUT81), .Z(new_n609));
  INV_X1    g0409(.A(new_n309), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n301), .A2(new_n306), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n386), .A2(new_n387), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n418), .A2(new_n405), .B1(new_n422), .B2(new_n336), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n612), .B1(new_n613), .B2(new_n378), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n610), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n609), .A2(new_n615), .ZN(G369));
  NAND2_X1  g0416(.A1(new_n506), .A2(new_n595), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n414), .A2(G20), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n259), .ZN(new_n619));
  OR2_X1    g0419(.A1(new_n619), .A2(KEYINPUT27), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(KEYINPUT27), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(G213), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT82), .ZN(new_n623));
  XNOR2_X1  g0423(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(G343), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n494), .ZN(new_n627));
  MUX2_X1   g0427(.A(new_n506), .B(new_n617), .S(new_n627), .Z(new_n628));
  INV_X1    g0428(.A(G330), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n480), .A2(new_n626), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n476), .A2(new_n626), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n469), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n631), .B1(new_n480), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(new_n480), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n506), .A2(new_n626), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n631), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n635), .A2(new_n638), .ZN(G399));
  NOR2_X1   g0439(.A1(new_n566), .A2(G116), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n640), .B(KEYINPUT83), .ZN(new_n641));
  INV_X1    g0441(.A(new_n216), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n642), .A2(G41), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n641), .A2(new_n259), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n644), .B1(new_n209), .B2(new_n643), .ZN(new_n645));
  XOR2_X1   g0445(.A(new_n645), .B(KEYINPUT28), .Z(new_n646));
  AOI22_X1  g0446(.A1(new_n528), .A2(new_n537), .B1(new_n551), .B2(new_n549), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n605), .B1(new_n647), .B2(new_n592), .ZN(new_n648));
  INV_X1    g0448(.A(new_n604), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n550), .A2(G169), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n550), .A2(new_n478), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n557), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n583), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n586), .A2(G200), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n653), .A2(new_n654), .A3(new_n571), .A4(new_n572), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n604), .A2(new_n655), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n652), .A2(new_n656), .A3(KEYINPUT26), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n648), .A2(new_n649), .A3(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n598), .A2(new_n597), .A3(new_n469), .A4(new_n592), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n626), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XOR2_X1   g0460(.A(KEYINPUT85), .B(KEYINPUT29), .Z(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT86), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n626), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n599), .B2(new_n607), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT86), .ZN(new_n665));
  INV_X1    g0465(.A(new_n661), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n647), .A2(new_n605), .A3(new_n592), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n592), .A2(new_n552), .A3(new_n557), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n649), .B1(new_n669), .B2(KEYINPUT26), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n659), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n671), .A2(KEYINPUT29), .A3(new_n663), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n662), .A2(new_n667), .A3(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n593), .A2(new_n507), .A3(new_n595), .A4(new_n663), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n590), .B1(new_n463), .B2(new_n464), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n499), .A2(new_n478), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n675), .A2(new_n676), .A3(new_n550), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT84), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n550), .A2(new_n586), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n680), .A2(KEYINPUT30), .A3(new_n503), .A4(new_n463), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT30), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n503), .A2(new_n463), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n546), .A2(new_n590), .A3(new_n464), .A4(new_n547), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n675), .A2(new_n676), .A3(KEYINPUT84), .A4(new_n550), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n679), .A2(new_n681), .A3(new_n685), .A4(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n626), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT31), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n681), .A2(new_n685), .A3(new_n677), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n691), .A2(KEYINPUT31), .A3(new_n626), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n674), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n673), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n646), .B1(new_n695), .B2(G1), .ZN(G364));
  NOR2_X1   g0496(.A1(G179), .A2(G200), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(G20), .A3(new_n274), .ZN(new_n698));
  INV_X1    g0498(.A(G329), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n371), .A2(G179), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n700), .A2(G20), .A3(G190), .ZN(new_n701));
  INV_X1    g0501(.A(G303), .ZN(new_n702));
  OAI221_X1 g0502(.A(new_n341), .B1(new_n698), .B2(new_n699), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n211), .A2(new_n478), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT89), .Z(new_n705));
  NAND3_X1  g0505(.A1(new_n705), .A2(new_n274), .A3(new_n371), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n703), .B1(new_n707), .B2(G311), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n700), .A2(G20), .A3(new_n274), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G283), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n704), .A2(G190), .A3(G200), .ZN(new_n712));
  INV_X1    g0512(.A(G326), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n211), .B1(new_n697), .B2(G190), .ZN(new_n714));
  INV_X1    g0514(.A(G294), .ZN(new_n715));
  OAI22_X1  g0515(.A1(new_n712), .A2(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n704), .A2(new_n274), .A3(G200), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  XNOR2_X1  g0518(.A(KEYINPUT33), .B(G317), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n716), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n705), .A2(G190), .A3(new_n371), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G322), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n708), .A2(new_n711), .A3(new_n720), .A4(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n714), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G97), .ZN(new_n726));
  OAI221_X1 g0526(.A(new_n726), .B1(new_n204), .B2(new_n712), .C1(new_n221), .C2(new_n717), .ZN(new_n727));
  INV_X1    g0527(.A(new_n701), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n727), .B1(G87), .B2(new_n728), .ZN(new_n729));
  OAI221_X1 g0529(.A(new_n249), .B1(new_n432), .B2(new_n709), .C1(new_n706), .C2(new_n313), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  XOR2_X1   g0531(.A(new_n721), .B(KEYINPUT90), .Z(new_n732));
  OAI211_X1 g0532(.A(new_n729), .B(new_n731), .C1(new_n732), .C2(new_n347), .ZN(new_n733));
  INV_X1    g0533(.A(G159), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n698), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT91), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT32), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n724), .B1(new_n733), .B2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n210), .B1(G20), .B2(new_n333), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n259), .B1(new_n618), .B2(G45), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n643), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n642), .A2(new_n249), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n209), .A2(new_n453), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n745), .B(new_n746), .C1(new_n241), .C2(new_n453), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n249), .A2(G355), .A3(new_n216), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n747), .B(new_n748), .C1(G116), .C2(new_n216), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT87), .ZN(new_n750));
  NOR2_X1   g0550(.A1(G13), .A2(G33), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT88), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n739), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n744), .B1(new_n750), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n740), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT92), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n628), .A2(new_n754), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n628), .A2(new_n629), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n744), .B1(new_n628), .B2(new_n629), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(new_n761), .ZN(G396));
  NOR2_X1   g0562(.A1(new_n335), .A2(new_n626), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n322), .A2(new_n626), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n764), .B1(new_n329), .B2(new_n330), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n763), .B1(new_n765), .B2(new_n335), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n664), .A2(new_n767), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n663), .B(new_n766), .C1(new_n599), .C2(new_n607), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(new_n694), .Z(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n744), .ZN(new_n772));
  INV_X1    g0572(.A(G132), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n698), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n709), .A2(new_n221), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n249), .B1(new_n701), .B2(new_n204), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n775), .B(new_n776), .C1(G58), .C2(new_n725), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n707), .A2(G159), .B1(G150), .B2(new_n718), .ZN(new_n778));
  INV_X1    g0578(.A(G137), .ZN(new_n779));
  INV_X1    g0579(.A(G143), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n778), .B1(new_n779), .B2(new_n712), .C1(new_n732), .C2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT94), .ZN(new_n782));
  INV_X1    g0582(.A(KEYINPUT34), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n777), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n774), .B(new_n784), .C1(new_n783), .C2(new_n782), .ZN(new_n785));
  XOR2_X1   g0585(.A(KEYINPUT93), .B(G283), .Z(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n726), .B1(new_n702), .B2(new_n712), .C1(new_n717), .C2(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n341), .B1(new_n701), .B2(new_n432), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(G87), .B2(new_n710), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n790), .B1(new_n721), .B2(new_n715), .C1(new_n488), .C2(new_n706), .ZN(new_n791));
  INV_X1    g0591(.A(new_n698), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n788), .B(new_n791), .C1(G311), .C2(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n739), .B1(new_n785), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n744), .B1(new_n767), .B2(new_n752), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n739), .A2(new_n751), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n794), .B(new_n795), .C1(G77), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n772), .A2(new_n798), .ZN(G384));
  INV_X1    g0599(.A(KEYINPUT38), .ZN(new_n800));
  INV_X1    g0600(.A(new_n624), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n380), .A2(new_n801), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n376), .A2(new_n377), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n802), .B1(new_n803), .B2(new_n612), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n380), .B1(new_n385), .B2(new_n801), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT37), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n805), .A2(new_n806), .A3(new_n374), .ZN(new_n807));
  AND3_X1   g0607(.A1(new_n354), .A2(new_n357), .A3(new_n373), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n354), .A2(new_n357), .B1(new_n384), .B2(new_n624), .ZN(new_n809));
  OAI21_X1  g0609(.A(KEYINPUT37), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n800), .B1(new_n804), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n807), .A2(new_n810), .ZN(new_n813));
  OAI211_X1 g0613(.A(KEYINPUT38), .B(new_n813), .C1(new_n388), .C2(new_n802), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n812), .A2(KEYINPUT96), .A3(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT96), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n816), .B(new_n800), .C1(new_n804), .C2(new_n811), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT100), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n818), .B1(new_n688), .B2(new_n689), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(new_n690), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n688), .A2(new_n818), .A3(new_n689), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n820), .A2(new_n674), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n626), .A2(new_n418), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n419), .A2(new_n422), .A3(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n422), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n418), .B(new_n626), .C1(new_n825), .C2(new_n405), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n767), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n815), .A2(new_n817), .A3(new_n822), .A4(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT40), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT97), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n810), .B(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT98), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n808), .A2(new_n809), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n833), .B1(new_n834), .B2(new_n806), .ZN(new_n835));
  NOR4_X1   g0635(.A1(new_n808), .A2(new_n809), .A3(KEYINPUT98), .A4(KEYINPUT37), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n804), .B1(new_n832), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n814), .B1(new_n838), .B2(KEYINPUT38), .ZN(new_n839));
  NAND4_X1  g0639(.A1(new_n839), .A2(KEYINPUT40), .A3(new_n822), .A4(new_n827), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n830), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n425), .A2(new_n822), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n841), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(G330), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n662), .A2(new_n667), .A3(new_n425), .A4(new_n672), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n615), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT99), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n844), .B(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n815), .A2(KEYINPUT39), .A3(new_n817), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT39), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n850), .B(new_n814), .C1(new_n838), .C2(KEYINPUT38), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n419), .A2(new_n626), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n612), .A2(new_n801), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n815), .A2(new_n817), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n826), .A2(new_n824), .ZN(new_n857));
  INV_X1    g0657(.A(new_n763), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n857), .B1(new_n769), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n855), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n848), .B(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n259), .B2(new_n618), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n532), .A2(new_n533), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n488), .B1(new_n864), .B2(KEYINPUT35), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n865), .B(new_n212), .C1(KEYINPUT35), .C2(new_n864), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT36), .ZN(new_n867));
  NOR4_X1   g0667(.A1(new_n203), .A2(new_n204), .A3(new_n313), .A4(new_n348), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n204), .A2(G68), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n869), .B(KEYINPUT95), .ZN(new_n870));
  OAI211_X1 g0670(.A(G1), .B(new_n414), .C1(new_n868), .C2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n863), .A2(new_n867), .A3(new_n871), .ZN(G367));
  INV_X1    g0672(.A(KEYINPUT45), .ZN(new_n873));
  INV_X1    g0673(.A(new_n638), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n652), .A2(new_n663), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n557), .A2(new_n626), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n553), .A2(new_n559), .A3(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT102), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n598), .A2(KEYINPUT102), .A3(new_n876), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n875), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n873), .B1(new_n874), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n879), .A2(new_n880), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n552), .A2(new_n557), .A3(new_n626), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n885), .A2(KEYINPUT45), .A3(new_n638), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT106), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT44), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n874), .A2(new_n881), .A3(new_n888), .A4(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  NAND2_X1  g0691(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n891), .B(new_n892), .C1(new_n885), .C2(new_n638), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n887), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n635), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n887), .A2(new_n635), .A3(new_n890), .A4(new_n893), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n634), .B(new_n637), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(new_n630), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n695), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n643), .B(KEYINPUT41), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n742), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OR3_X1    g0704(.A1(new_n663), .A2(new_n604), .A3(new_n573), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n592), .B1(new_n573), .B2(new_n663), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  MUX2_X1   g0707(.A(new_n905), .B(new_n907), .S(KEYINPUT101), .Z(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(KEYINPUT43), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT104), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n553), .B1(new_n881), .B2(new_n480), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n663), .ZN(new_n912));
  INV_X1    g0712(.A(new_n631), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n636), .A2(new_n913), .A3(new_n637), .ZN(new_n914));
  OAI21_X1  g0714(.A(KEYINPUT42), .B1(new_n881), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT103), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n912), .A2(KEYINPUT103), .A3(new_n915), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n881), .A2(new_n914), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n921), .A2(KEYINPUT42), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n910), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  AOI211_X1 g0724(.A(KEYINPUT104), .B(new_n922), .C1(new_n918), .C2(new_n919), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n909), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n919), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT103), .B1(new_n912), .B2(new_n915), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n923), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(KEYINPUT104), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n908), .B(KEYINPUT43), .Z(new_n931));
  NAND3_X1  g0731(.A1(new_n920), .A2(new_n910), .A3(new_n923), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n926), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n635), .A2(new_n881), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n904), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n926), .A2(new_n933), .A3(new_n935), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT105), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT105), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n926), .A2(new_n933), .A3(new_n940), .A4(new_n935), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n937), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  OAI221_X1 g0742(.A(new_n249), .B1(new_n709), .B2(new_n313), .C1(new_n347), .C2(new_n701), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(new_n722), .B2(G150), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n717), .A2(new_n734), .B1(new_n712), .B2(new_n780), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(G68), .B2(new_n725), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n944), .B(new_n946), .C1(new_n204), .C2(new_n706), .ZN(new_n947));
  XOR2_X1   g0747(.A(KEYINPUT108), .B(G137), .Z(new_n948));
  AOI21_X1  g0748(.A(new_n947), .B1(new_n792), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n707), .A2(new_n786), .ZN(new_n950));
  INV_X1    g0750(.A(G311), .ZN(new_n951));
  OAI22_X1  g0751(.A1(new_n717), .A2(new_n715), .B1(new_n712), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n952), .B1(G107), .B2(new_n725), .ZN(new_n953));
  OAI21_X1  g0753(.A(KEYINPUT107), .B1(new_n701), .B2(new_n488), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n954), .A2(KEYINPUT46), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n249), .B1(new_n792), .B2(G317), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n954), .A2(KEYINPUT46), .B1(G97), .B2(new_n710), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n953), .A2(new_n955), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n732), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n958), .B1(new_n959), .B2(G303), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n949), .B1(new_n950), .B2(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT47), .Z(new_n962));
  AOI21_X1  g0762(.A(new_n744), .B1(new_n962), .B2(new_n739), .ZN(new_n963));
  INV_X1    g0763(.A(new_n745), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n755), .B1(new_n216), .B2(new_n318), .C1(new_n237), .C2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n754), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n963), .B(new_n965), .C1(new_n908), .C2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n942), .A2(new_n967), .ZN(G387));
  OR2_X1    g0768(.A1(new_n695), .A2(new_n900), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n695), .A2(new_n900), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n969), .A2(new_n643), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n725), .A2(new_n317), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n721), .B2(new_n204), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT110), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n706), .A2(new_n221), .B1(new_n283), .B2(new_n717), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n341), .B1(new_n710), .B2(G97), .ZN(new_n976));
  XNOR2_X1  g0776(.A(KEYINPUT109), .B(G150), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n792), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n976), .B(new_n978), .C1(new_n734), .C2(new_n712), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n975), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n728), .A2(G77), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n974), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT111), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n707), .A2(G303), .B1(G311), .B2(new_n718), .ZN(new_n984));
  INV_X1    g0784(.A(G322), .ZN(new_n985));
  INV_X1    g0785(.A(G317), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n984), .B1(new_n985), .B2(new_n712), .C1(new_n732), .C2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT48), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n715), .B2(new_n701), .C1(new_n714), .C2(new_n787), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT49), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n249), .B1(new_n792), .B2(G326), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n709), .A2(new_n488), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n983), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AND2_X1   g0796(.A1(new_n996), .A2(new_n739), .ZN(new_n997));
  INV_X1    g0797(.A(new_n281), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n204), .ZN(new_n999));
  AOI21_X1  g0799(.A(G45), .B1(new_n999), .B2(KEYINPUT50), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(KEYINPUT50), .B2(new_n999), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n641), .B(new_n1001), .C1(G68), .C2(G77), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n745), .B1(new_n234), .B2(new_n453), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n641), .A2(new_n216), .A3(new_n249), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1002), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n216), .A2(G107), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n755), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n743), .B(new_n1007), .C1(new_n634), .C2(new_n966), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n971), .B1(new_n741), .B2(new_n901), .C1(new_n997), .C2(new_n1008), .ZN(G393));
  AOI211_X1 g0809(.A(G41), .B(new_n642), .C1(new_n898), .C2(new_n970), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n898), .B2(new_n970), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n896), .A2(new_n742), .A3(new_n897), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n755), .B1(new_n486), .B2(new_n216), .C1(new_n244), .C2(new_n964), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n721), .A2(new_n734), .B1(new_n278), .B2(new_n712), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT51), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n717), .A2(new_n204), .B1(new_n714), .B2(new_n313), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n249), .B1(new_n698), .B2(new_n780), .C1(new_n709), .C2(new_n565), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1016), .B(new_n1017), .C1(new_n707), .C2(new_n998), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1015), .B(new_n1018), .C1(new_n221), .C2(new_n701), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n249), .B1(new_n710), .B2(G107), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1020), .B1(new_n985), .B2(new_n698), .C1(new_n701), .C2(new_n787), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT112), .Z(new_n1022));
  OAI22_X1  g0822(.A1(new_n721), .A2(new_n951), .B1(new_n986), .B2(new_n712), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT52), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n707), .A2(G294), .B1(G303), .B2(new_n718), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1022), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n714), .A2(new_n488), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1019), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n744), .B1(new_n1028), .B2(new_n739), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1013), .B(new_n1029), .C1(new_n885), .C2(new_n966), .ZN(new_n1030));
  AND2_X1   g0830(.A1(new_n1012), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1011), .A2(new_n1031), .ZN(G390));
  NAND2_X1  g0832(.A1(new_n826), .A2(new_n824), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n767), .A2(new_n629), .ZN(new_n1034));
  AND3_X1   g0834(.A1(new_n822), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n849), .B(new_n851), .C1(new_n859), .C2(new_n853), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n853), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n765), .A2(new_n335), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n671), .A2(new_n663), .A3(new_n1038), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1039), .A2(new_n858), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1037), .B(new_n839), .C1(new_n1040), .C2(new_n857), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1035), .B1(new_n1036), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n693), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1044));
  AND2_X1   g0844(.A1(new_n822), .A2(new_n1034), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1040), .B(new_n1044), .C1(new_n1045), .C2(new_n1033), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n769), .A2(new_n858), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1033), .B1(new_n693), .B2(new_n1034), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1047), .B1(new_n1035), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n425), .A2(G330), .A3(new_n822), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n845), .A2(new_n615), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1050), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1044), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1036), .A2(new_n1041), .A3(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1043), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1052), .B1(new_n1049), .B2(new_n1046), .ZN(new_n1058));
  AND3_X1   g0858(.A1(new_n1036), .A2(new_n1041), .A3(new_n1055), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1058), .B1(new_n1059), .B2(new_n1042), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1057), .A2(new_n1060), .A3(new_n643), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n706), .A2(new_n486), .B1(new_n432), .B2(new_n717), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT115), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1065));
  INV_X1    g0865(.A(G283), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1064), .B(new_n1065), .C1(new_n1066), .C2(new_n712), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1067), .A2(KEYINPUT116), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n775), .B1(G77), .B2(new_n725), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(KEYINPUT116), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n341), .B1(new_n698), .B2(new_n715), .C1(new_n701), .C2(new_n565), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n722), .B2(G116), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n718), .A2(new_n948), .ZN(new_n1074));
  XOR2_X1   g0874(.A(KEYINPUT54), .B(G143), .Z(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1074), .B1(new_n734), .B2(new_n714), .C1(new_n706), .C2(new_n1076), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT113), .Z(new_n1078));
  NAND2_X1  g0878(.A1(new_n728), .A2(new_n977), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1079), .A2(KEYINPUT53), .B1(G125), .B2(new_n792), .ZN(new_n1080));
  INV_X1    g0880(.A(G128), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1080), .B1(KEYINPUT53), .B2(new_n1079), .C1(new_n1081), .C2(new_n712), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(G132), .B2(new_n722), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n249), .B1(new_n709), .B2(new_n204), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT114), .Z(new_n1085));
  NAND3_X1  g0885(.A1(new_n1078), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1073), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n744), .B1(new_n1087), .B2(new_n739), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n852), .B2(new_n753), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n283), .B2(new_n796), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1043), .A2(new_n1056), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1090), .B1(new_n1091), .B2(new_n742), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1061), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(G378));
  NAND2_X1  g0894(.A1(new_n1060), .A2(new_n1053), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n830), .A2(G330), .A3(new_n840), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n861), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n611), .A2(new_n309), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT55), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n296), .A2(new_n801), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT56), .Z(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1098), .A2(KEYINPUT55), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1098), .A2(KEYINPUT55), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1104), .A2(new_n1105), .A3(new_n1101), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n830), .A2(G330), .A3(new_n840), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1108), .A2(new_n854), .A3(new_n860), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n1097), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1107), .B1(new_n1097), .B2(new_n1109), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1095), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT57), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1095), .B(KEYINPUT57), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1114), .A2(new_n643), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1103), .A2(new_n752), .A3(new_n1106), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n725), .A2(G150), .ZN(new_n1118));
  INV_X1    g0918(.A(G125), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n1118), .B1(new_n1119), .B2(new_n712), .C1(new_n701), .C2(new_n1076), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n1081), .A2(new_n721), .B1(new_n706), .B2(new_n779), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1120), .B(new_n1121), .C1(G132), .C2(new_n718), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT119), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT59), .ZN(new_n1124));
  OR2_X1    g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1126));
  AOI21_X1  g0926(.A(G33), .B1(new_n792), .B2(G124), .ZN(new_n1127));
  AOI21_X1  g0927(.A(G41), .B1(new_n710), .B2(G159), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n981), .B1(new_n347), .B2(new_n709), .C1(new_n1066), .C2(new_n698), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n707), .B2(new_n317), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n722), .A2(G107), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n712), .A2(new_n488), .B1(new_n714), .B2(new_n221), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n249), .B(new_n1133), .C1(G97), .C2(new_n718), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1131), .A2(new_n255), .A3(new_n1132), .A4(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT117), .ZN(new_n1140));
  AOI21_X1  g0940(.A(G50), .B1(new_n248), .B2(new_n255), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1138), .B(new_n1139), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1129), .B(new_n1142), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n744), .B1(new_n1143), .B2(new_n739), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1117), .B(new_n1144), .C1(G50), .C2(new_n797), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT120), .ZN(new_n1146));
  OR2_X1    g0946(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1146), .B1(new_n742), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1116), .A2(new_n1148), .ZN(G375));
  OAI221_X1 g0949(.A(new_n341), .B1(new_n698), .B2(new_n702), .C1(new_n709), .C2(new_n313), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n707), .B2(G107), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n728), .A2(G97), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n972), .B1(new_n488), .B2(new_n717), .C1(new_n715), .C2(new_n712), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n722), .A2(G283), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n959), .A2(new_n948), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n712), .A2(new_n773), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n718), .A2(new_n1075), .B1(new_n725), .B2(G50), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n249), .B1(new_n698), .B2(new_n1081), .C1(new_n709), .C2(new_n347), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n707), .B2(G150), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .A4(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n701), .A2(new_n734), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1156), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n744), .B1(new_n1164), .B2(new_n739), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n751), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n1033), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n221), .B2(new_n796), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n1050), .B2(new_n742), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n903), .B(KEYINPUT121), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1054), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1050), .A2(new_n1053), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1169), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  XOR2_X1   g0973(.A(new_n1173), .B(KEYINPUT122), .Z(G381));
  NAND3_X1  g0974(.A1(new_n1116), .A2(new_n1093), .A3(new_n1148), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NOR3_X1   g0976(.A1(G381), .A2(G384), .A3(G390), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  OR3_X1    g0978(.A1(G387), .A2(G396), .A3(G393), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT123), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1178), .A2(new_n1179), .A3(KEYINPUT123), .ZN(new_n1183));
  OR2_X1    g0983(.A1(new_n1182), .A2(new_n1183), .ZN(G407));
  INV_X1    g0984(.A(G213), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1185), .A2(G343), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1176), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1185), .B1(new_n1187), .B2(KEYINPUT124), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(KEYINPUT124), .B2(new_n1187), .C1(new_n1182), .C2(new_n1183), .ZN(G409));
  NOR2_X1   g0989(.A1(new_n1172), .A2(KEYINPUT60), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1052), .A2(new_n1046), .A3(new_n1049), .A4(KEYINPUT60), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1054), .A2(new_n1191), .A3(new_n643), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1169), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1193), .A2(new_n772), .A3(new_n798), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT125), .ZN(new_n1195));
  OAI211_X1 g0995(.A(G384), .B(new_n1169), .C1(new_n1190), .C2(new_n1192), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1195), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1186), .A2(G2897), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1197), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1093), .B1(new_n1116), .B2(new_n1148), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n742), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1095), .B(new_n1170), .C1(new_n1110), .C2(new_n1111), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1093), .A2(new_n1203), .A3(new_n1204), .A4(new_n1145), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1186), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1200), .B(new_n1201), .C1(new_n1202), .C2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT61), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT62), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1202), .A2(new_n1212), .A3(new_n1207), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT127), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1211), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(G375), .A2(G378), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1212), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1207), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1219), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1210), .A2(new_n1215), .A3(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(G393), .B(G396), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n942), .A2(G390), .A3(new_n967), .ZN(new_n1223));
  AOI21_X1  g1023(.A(G390), .B1(new_n942), .B2(new_n967), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1222), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(G390), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(G387), .A2(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n942), .A2(G390), .A3(new_n967), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1222), .A2(KEYINPUT126), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1224), .A2(KEYINPUT126), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1225), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1221), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT63), .ZN(new_n1234));
  NOR4_X1   g1034(.A1(new_n1202), .A2(new_n1207), .A3(new_n1234), .A4(new_n1212), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1232), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1208), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1219), .B1(new_n1237), .B2(new_n1234), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1238), .A3(new_n1209), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1233), .A2(new_n1239), .ZN(G405));
  NOR3_X1   g1040(.A1(new_n1176), .A2(new_n1217), .A3(new_n1202), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1212), .B1(new_n1216), .B2(new_n1175), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(new_n1232), .ZN(G402));
endmodule


