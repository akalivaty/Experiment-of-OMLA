//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1280, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(new_n207), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(G50), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n212), .B1(new_n215), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G226), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT65), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n232), .B(new_n233), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XOR2_X1   g0039(.A(G50), .B(G58), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  XNOR2_X1  g0045(.A(KEYINPUT66), .B(KEYINPUT8), .ZN(new_n246));
  INV_X1    g0046(.A(G58), .ZN(new_n247));
  OR3_X1    g0047(.A1(new_n246), .A2(KEYINPUT67), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(KEYINPUT8), .ZN(new_n249));
  OAI211_X1 g0049(.A(KEYINPUT67), .B(new_n249), .C1(new_n246), .C2(new_n247), .ZN(new_n250));
  AND2_X1   g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G20), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n218), .A2(new_n247), .A3(new_n220), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  AOI22_X1  g0056(.A1(new_n255), .A2(G20), .B1(G150), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n254), .A2(new_n257), .B1(new_n213), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(new_n213), .A3(new_n258), .ZN(new_n261));
  OR2_X1    g0061(.A1(new_n261), .A2(KEYINPUT68), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n206), .A2(G20), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(KEYINPUT68), .ZN(new_n264));
  AND3_X1   g0064(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G50), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G50), .B2(new_n260), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n259), .A2(new_n267), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n268), .A2(KEYINPUT9), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(KEYINPUT9), .ZN(new_n270));
  INV_X1    g0070(.A(G41), .ZN(new_n271));
  INV_X1    g0071(.A(G45), .ZN(new_n272));
  AOI21_X1  g0072(.A(G1), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G1), .A3(G13), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(new_n275), .A3(G274), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n276), .B1(new_n219), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT3), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n252), .ZN(new_n282));
  NAND2_X1  g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n280), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AND2_X1   g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NOR2_X1   g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n284), .A2(G223), .B1(new_n287), .B2(G77), .ZN(new_n288));
  AOI21_X1  g0088(.A(G1698), .B1(new_n282), .B2(new_n283), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G222), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n279), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G200), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n295), .B1(G190), .B2(new_n293), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n269), .A2(new_n270), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT10), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT10), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n269), .A2(new_n299), .A3(new_n270), .A4(new_n296), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G179), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n293), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(G169), .B2(new_n293), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n268), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  XOR2_X1   g0107(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n308));
  NAND2_X1  g0108(.A1(new_n219), .A2(new_n280), .ZN(new_n309));
  INV_X1    g0109(.A(G232), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G1698), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n309), .B(new_n311), .C1(new_n285), .C2(new_n286), .ZN(new_n312));
  NAND2_X1  g0112(.A1(G33), .A2(G97), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n275), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n275), .A2(G238), .A3(new_n277), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n276), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n308), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT70), .ZN(new_n318));
  OR3_X1    g0118(.A1(new_n314), .A2(new_n316), .A3(new_n308), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT70), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n320), .B(new_n308), .C1(new_n314), .C2(new_n316), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n318), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G169), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT14), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT13), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n314), .A2(new_n316), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n319), .B(G179), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT14), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n322), .A2(new_n328), .A3(G169), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n324), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n260), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n220), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n332), .B(KEYINPUT12), .ZN(new_n333));
  AOI22_X1  g0133(.A1(new_n253), .A2(G77), .B1(G20), .B2(new_n220), .ZN(new_n334));
  INV_X1    g0134(.A(new_n256), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n334), .B1(new_n218), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n258), .A2(new_n213), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(KEYINPUT11), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n261), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n339), .A2(G68), .A3(new_n263), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n333), .A2(new_n338), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT11), .B1(new_n336), .B2(new_n337), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n330), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n322), .A2(G200), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT71), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n322), .A2(KEYINPUT71), .A3(G200), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n319), .B(G190), .C1(new_n325), .C2(new_n326), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n351), .A2(new_n343), .ZN(new_n352));
  AOI21_X1  g0152(.A(KEYINPUT72), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  AND3_X1   g0153(.A1(new_n322), .A2(KEYINPUT71), .A3(G200), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT71), .B1(new_n322), .B2(G200), .ZN(new_n355));
  OAI211_X1 g0155(.A(KEYINPUT72), .B(new_n352), .C1(new_n354), .C2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n345), .B1(new_n353), .B2(new_n357), .ZN(new_n358));
  XOR2_X1   g0158(.A(KEYINPUT8), .B(G58), .Z(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n360), .A2(new_n335), .ZN(new_n361));
  XNOR2_X1  g0161(.A(KEYINPUT15), .B(G87), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n207), .A2(G33), .ZN(new_n363));
  INV_X1    g0163(.A(G77), .ZN(new_n364));
  OAI22_X1  g0164(.A1(new_n362), .A2(new_n363), .B1(new_n207), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n337), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n364), .B1(new_n206), .B2(G20), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n339), .A2(new_n367), .B1(new_n364), .B2(new_n331), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n282), .A2(new_n283), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n310), .A2(new_n280), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n221), .A2(G1698), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n375), .B(new_n292), .C1(G107), .C2(new_n371), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n275), .A2(G244), .A3(new_n277), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(new_n276), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G200), .ZN(new_n379));
  INV_X1    g0179(.A(G190), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n370), .B(new_n379), .C1(new_n380), .C2(new_n378), .ZN(new_n381));
  INV_X1    g0181(.A(G169), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n376), .A2(new_n302), .A3(new_n276), .A4(new_n377), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n369), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n381), .A2(new_n385), .ZN(new_n386));
  OR3_X1    g0186(.A1(new_n307), .A2(new_n358), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT7), .B1(new_n287), .B2(new_n207), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n282), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n283), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(G68), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  AND2_X1   g0191(.A1(G58), .A2(G68), .ZN(new_n392));
  NOR2_X1   g0192(.A1(G58), .A2(G68), .ZN(new_n393));
  OAI21_X1  g0193(.A(G20), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G159), .ZN(new_n395));
  NOR4_X1   g0195(.A1(new_n395), .A2(KEYINPUT73), .A3(G20), .A4(G33), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT73), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(new_n256), .B2(G159), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n394), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT74), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT74), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n401), .B(new_n394), .C1(new_n396), .C2(new_n398), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n391), .A2(new_n400), .A3(KEYINPUT16), .A4(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT16), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n282), .A2(new_n207), .A3(new_n283), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT7), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n220), .B1(new_n407), .B2(new_n389), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n404), .B1(new_n408), .B2(new_n399), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n403), .A2(new_n409), .A3(new_n337), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT75), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n260), .B1(new_n248), .B2(new_n250), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n265), .B2(new_n251), .ZN(new_n413));
  AND3_X1   g0213(.A1(new_n410), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n411), .B1(new_n410), .B2(new_n413), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT18), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n219), .A2(G1698), .ZN(new_n418));
  OAI221_X1 g0218(.A(new_n418), .B1(G223), .B2(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G33), .A2(G87), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n292), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n276), .B1(new_n310), .B2(new_n278), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(G169), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n302), .B2(new_n425), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n416), .A2(new_n417), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n410), .A2(new_n413), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT75), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n410), .A2(new_n411), .A3(new_n413), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n430), .A2(new_n431), .A3(new_n427), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT18), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n422), .A2(new_n424), .A3(new_n380), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n275), .B1(new_n419), .B2(new_n420), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n294), .B1(new_n435), .B2(new_n423), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n410), .A2(new_n413), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n410), .A2(new_n413), .A3(new_n437), .A4(KEYINPUT17), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n428), .A2(new_n433), .A3(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n387), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT77), .ZN(new_n446));
  OAI211_X1 g0246(.A(G250), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT76), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT76), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n371), .A2(new_n449), .A3(G250), .A4(G1698), .ZN(new_n450));
  AND2_X1   g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(G244), .B(new_n280), .C1(new_n285), .C2(new_n286), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT4), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(G33), .A2(G283), .ZN(new_n455));
  INV_X1    g0255(.A(G244), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n371), .A2(new_n280), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n454), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n446), .B1(new_n451), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n448), .A2(new_n450), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n289), .A2(new_n457), .B1(G33), .B2(G283), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n461), .A2(KEYINPUT77), .A3(new_n454), .A4(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n460), .A2(new_n292), .A3(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n271), .A2(KEYINPUT5), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n206), .A2(G45), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n271), .A2(KEYINPUT5), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n292), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G257), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n468), .B(KEYINPUT78), .ZN(new_n471));
  INV_X1    g0271(.A(G274), .ZN(new_n472));
  INV_X1    g0272(.A(new_n213), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n472), .B1(new_n473), .B2(new_n274), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n471), .A2(new_n474), .A3(new_n467), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n464), .A2(new_n302), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT6), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n479), .A2(new_n202), .A3(G107), .ZN(new_n480));
  XNOR2_X1  g0280(.A(G97), .B(G107), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n480), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  OAI22_X1  g0282(.A1(new_n482), .A2(new_n207), .B1(new_n364), .B2(new_n335), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n203), .B1(new_n407), .B2(new_n389), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n337), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n331), .A2(new_n202), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n206), .A2(G33), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n260), .A2(new_n487), .A3(new_n213), .A4(new_n258), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G97), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n485), .A2(new_n486), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n449), .B1(new_n284), .B2(G250), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n447), .A2(KEYINPUT76), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n462), .B(new_n454), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n275), .B1(new_n494), .B2(new_n446), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n476), .B1(new_n495), .B2(new_n463), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n478), .B(new_n491), .C1(G169), .C2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n464), .A2(G190), .A3(new_n477), .ZN(new_n498));
  INV_X1    g0298(.A(new_n491), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n498), .B(new_n499), .C1(new_n294), .C2(new_n496), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n272), .A2(G1), .ZN(new_n501));
  OR2_X1    g0301(.A1(new_n501), .A2(G250), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n472), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n502), .A2(new_n275), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n221), .A2(new_n280), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n456), .A2(G1698), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n506), .B(new_n507), .C1(new_n285), .C2(new_n286), .ZN(new_n508));
  INV_X1    g0308(.A(G116), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n252), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT79), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n275), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(G238), .A2(G1698), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n515), .B1(new_n456), .B2(G1698), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n510), .B1(new_n516), .B2(new_n371), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT79), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n505), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n302), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n292), .B1(new_n517), .B2(KEYINPUT79), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n508), .A2(KEYINPUT79), .A3(new_n511), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n504), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n488), .A2(new_n362), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT80), .ZN(new_n525));
  XNOR2_X1  g0325(.A(new_n524), .B(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT19), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n207), .B1(new_n313), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(G87), .B2(new_n204), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n527), .B1(new_n363), .B2(new_n202), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n207), .B(G68), .C1(new_n285), .C2(new_n286), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n532), .A2(new_n337), .B1(new_n331), .B2(new_n362), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n523), .A2(new_n382), .B1(new_n526), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n337), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n489), .A2(G87), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n362), .A2(new_n331), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(G190), .B2(new_n519), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n523), .A2(G200), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n520), .A2(new_n534), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n497), .A2(new_n500), .A3(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(G257), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n543));
  OAI211_X1 g0343(.A(G250), .B(new_n280), .C1(new_n285), .C2(new_n286), .ZN(new_n544));
  NAND2_X1  g0344(.A1(G33), .A2(G294), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n292), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n469), .A2(G264), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT83), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n549), .A2(new_n550), .A3(G179), .A4(new_n475), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(new_n548), .A3(new_n475), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT83), .B1(new_n552), .B2(G169), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n552), .A2(new_n302), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n551), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n207), .B(G87), .C1(new_n285), .C2(new_n286), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT22), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT22), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n371), .A2(new_n558), .A3(new_n207), .A4(G87), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT24), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT23), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n207), .B2(G107), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n203), .A2(KEYINPUT23), .A3(G20), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n563), .A2(new_n564), .B1(new_n510), .B2(new_n207), .ZN(new_n565));
  AND3_X1   g0365(.A1(new_n560), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n561), .B1(new_n560), .B2(new_n565), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n337), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT25), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n260), .B2(G107), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n260), .A2(new_n569), .A3(G107), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n570), .A2(new_n572), .B1(new_n489), .B2(G107), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n555), .A2(new_n574), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n552), .A2(new_n294), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n552), .A2(G190), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n568), .B(new_n573), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(G264), .B(G1698), .C1(new_n285), .C2(new_n286), .ZN(new_n580));
  OAI211_X1 g0380(.A(G257), .B(new_n280), .C1(new_n285), .C2(new_n286), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n282), .A2(G303), .A3(new_n283), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT81), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n580), .A2(new_n581), .A3(KEYINPUT81), .A4(new_n582), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n292), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n469), .A2(G270), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n475), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n588), .A2(G190), .A3(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n455), .B(new_n207), .C1(G33), .C2(new_n202), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n509), .A2(G20), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n337), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT20), .ZN(new_n596));
  XNOR2_X1  g0396(.A(new_n595), .B(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n260), .A2(G116), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n489), .B2(G116), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n275), .B1(new_n585), .B2(new_n586), .ZN(new_n602));
  OAI21_X1  g0402(.A(G200), .B1(new_n602), .B2(new_n590), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n592), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  XOR2_X1   g0404(.A(KEYINPUT82), .B(KEYINPUT21), .Z(new_n605));
  NAND2_X1  g0405(.A1(new_n600), .A2(G169), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n602), .A2(new_n590), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n589), .A2(new_n475), .A3(G179), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n600), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n382), .B1(new_n597), .B2(new_n599), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n612), .B(KEYINPUT21), .C1(new_n590), .C2(new_n602), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n604), .A2(new_n608), .A3(new_n611), .A4(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n579), .A2(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n445), .A2(new_n542), .A3(new_n615), .ZN(G372));
  OAI21_X1  g0416(.A(new_n352), .B1(new_n354), .B2(new_n355), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT72), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n356), .ZN(new_n620));
  INV_X1    g0420(.A(new_n385), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n442), .B1(new_n622), .B2(new_n345), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n429), .A2(new_n427), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT18), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n429), .A2(new_n417), .A3(new_n427), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n301), .B1(new_n623), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n628), .A2(new_n306), .ZN(new_n629));
  INV_X1    g0429(.A(new_n445), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT26), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n534), .A2(new_n520), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n539), .A2(new_n540), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n631), .B1(new_n497), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n464), .A2(new_n477), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n499), .B1(new_n636), .B2(new_n382), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n637), .A2(new_n541), .A3(KEYINPUT26), .A4(new_n478), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n632), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n578), .A2(new_n632), .A3(new_n633), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n641), .A2(KEYINPUT84), .A3(new_n497), .A4(new_n500), .ZN(new_n642));
  INV_X1    g0442(.A(new_n575), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n608), .A2(new_n611), .A3(new_n613), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n641), .A2(new_n497), .A3(new_n500), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT84), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n640), .B1(new_n642), .B2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n629), .B1(new_n630), .B2(new_n649), .ZN(G369));
  NAND3_X1  g0450(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n651), .A2(KEYINPUT27), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(G213), .A3(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(G343), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n601), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n644), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n614), .B2(new_n658), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n660), .A2(G330), .ZN(new_n661));
  INV_X1    g0461(.A(new_n579), .ZN(new_n662));
  INV_X1    g0462(.A(new_n574), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n662), .B1(new_n663), .B2(new_n657), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n643), .A2(new_n656), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n644), .A2(new_n657), .ZN(new_n668));
  XOR2_X1   g0468(.A(new_n656), .B(KEYINPUT85), .Z(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OAI22_X1  g0470(.A1(new_n668), .A2(new_n579), .B1(new_n575), .B2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT86), .ZN(G399));
  INV_X1    g0474(.A(new_n210), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G41), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n204), .A2(G87), .A3(G116), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G1), .A3(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n216), .B2(new_n677), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT28), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT29), .ZN(new_n682));
  OAI211_X1 g0482(.A(KEYINPUT89), .B(new_n682), .C1(new_n649), .C2(new_n670), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT89), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n497), .A2(new_n500), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n541), .A2(new_n578), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n647), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n645), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(new_n642), .A3(new_n688), .ZN(new_n689));
  AOI22_X1  g0489(.A1(new_n635), .A2(new_n638), .B1(new_n520), .B2(new_n534), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n670), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n684), .B1(new_n691), .B2(KEYINPUT29), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n690), .B1(new_n646), .B2(new_n645), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n693), .A2(KEYINPUT29), .A3(new_n657), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n683), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n464), .A2(new_n610), .A3(new_n477), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT87), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n519), .B2(new_n549), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n519), .A2(new_n549), .A3(new_n697), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n696), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n588), .A2(new_n591), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n514), .A2(new_n518), .ZN(new_n703));
  AOI21_X1  g0503(.A(G179), .B1(new_n703), .B2(new_n504), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n702), .A2(new_n552), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT30), .B1(new_n705), .B2(new_n496), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n701), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  AOI21_X1  g0508(.A(KEYINPUT79), .B1(new_n508), .B2(new_n511), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n522), .A2(new_n709), .A3(new_n275), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n552), .B(new_n302), .C1(new_n710), .C2(new_n505), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(new_n607), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n708), .B1(new_n712), .B2(new_n636), .ZN(new_n713));
  INV_X1    g0513(.A(new_n700), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n496), .B(new_n610), .C1(new_n714), .C2(new_n698), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n707), .A2(new_n656), .A3(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT31), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n542), .A2(new_n615), .A3(new_n669), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n707), .A2(new_n716), .A3(KEYINPUT31), .A4(new_n670), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n722), .A2(KEYINPUT88), .A3(G330), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT88), .B1(new_n722), .B2(G330), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n695), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n681), .B1(new_n726), .B2(G1), .ZN(G364));
  NOR2_X1   g0527(.A1(G13), .A2(G33), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n660), .A2(G20), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n213), .B1(G20), .B2(new_n382), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n207), .A2(new_n380), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n294), .A2(G179), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT94), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G303), .ZN(new_n738));
  INV_X1    g0538(.A(G283), .ZN(new_n739));
  OR3_X1    g0539(.A1(new_n207), .A2(KEYINPUT91), .A3(G190), .ZN(new_n740));
  OAI21_X1  g0540(.A(KEYINPUT91), .B1(new_n207), .B2(G190), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n740), .A2(new_n741), .A3(new_n734), .ZN(new_n742));
  OAI22_X1  g0542(.A1(new_n737), .A2(new_n738), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G179), .A2(G200), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n740), .A2(new_n744), .A3(new_n741), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n743), .B1(G329), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G190), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  XOR2_X1   g0550(.A(KEYINPUT33), .B(G317), .Z(new_n751));
  NOR2_X1   g0551(.A1(new_n302), .A2(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n733), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G322), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n750), .A2(new_n751), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT95), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n207), .B1(new_n744), .B2(G190), .ZN(new_n757));
  INV_X1    g0557(.A(G294), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n207), .A2(G190), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n752), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(G311), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n287), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n748), .A2(new_n380), .ZN(new_n764));
  XOR2_X1   g0564(.A(KEYINPUT93), .B(G326), .Z(new_n765));
  AOI211_X1 g0565(.A(new_n759), .B(new_n763), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n747), .A2(new_n756), .A3(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n753), .ZN(new_n768));
  INV_X1    g0568(.A(new_n735), .ZN(new_n769));
  AOI22_X1  g0569(.A1(G58), .A2(new_n768), .B1(new_n769), .B2(G87), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n770), .B(new_n371), .C1(new_n364), .C2(new_n761), .ZN(new_n771));
  INV_X1    g0571(.A(new_n742), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n771), .B1(G107), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n757), .A2(new_n202), .ZN(new_n774));
  INV_X1    g0574(.A(new_n764), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n218), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n774), .B(new_n776), .C1(G68), .C2(new_n749), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n745), .A2(new_n395), .ZN(new_n778));
  XOR2_X1   g0578(.A(KEYINPUT92), .B(KEYINPUT32), .Z(new_n779));
  XNOR2_X1  g0579(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n773), .A2(new_n777), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n732), .B1(new_n767), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n207), .A2(G13), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n206), .B1(new_n783), .B2(G45), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n676), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n210), .A2(new_n371), .ZN(new_n787));
  INV_X1    g0587(.A(G355), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n787), .A2(new_n788), .B1(G116), .B2(new_n210), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n210), .A2(new_n287), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT90), .Z(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n216), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n792), .B1(new_n272), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n241), .A2(G45), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n789), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n729), .A2(G20), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n731), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n786), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n730), .A2(new_n782), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n660), .A2(G330), .ZN(new_n802));
  NOR3_X1   g0602(.A1(new_n661), .A2(new_n802), .A3(new_n786), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(G396));
  NAND2_X1  g0605(.A1(new_n369), .A2(new_n656), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n381), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT97), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT96), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n385), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n383), .A2(new_n369), .A3(KEYINPUT96), .A4(new_n384), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n807), .A2(new_n808), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n621), .A2(new_n656), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n381), .A2(new_n806), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n810), .A2(new_n811), .ZN(new_n815));
  OAI21_X1  g0615(.A(KEYINPUT97), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AND3_X1   g0616(.A1(new_n812), .A2(new_n813), .A3(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n691), .B(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n786), .B1(new_n819), .B2(new_n725), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n725), .B2(new_n819), .ZN(new_n821));
  INV_X1    g0621(.A(new_n786), .ZN(new_n822));
  INV_X1    g0622(.A(new_n761), .ZN(new_n823));
  AOI22_X1  g0623(.A1(G143), .A2(new_n768), .B1(new_n823), .B2(G159), .ZN(new_n824));
  INV_X1    g0624(.A(G150), .ZN(new_n825));
  INV_X1    g0625(.A(G137), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n824), .B1(new_n750), .B2(new_n825), .C1(new_n826), .C2(new_n775), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT34), .ZN(new_n828));
  OR2_X1    g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n742), .A2(new_n220), .ZN(new_n831));
  INV_X1    g0631(.A(new_n757), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n287), .B(new_n831), .C1(G58), .C2(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n736), .A2(G50), .B1(G132), .B2(new_n746), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n829), .A2(new_n830), .A3(new_n833), .A4(new_n834), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n287), .B1(new_n761), .B2(new_n509), .C1(new_n758), .C2(new_n753), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G87), .B2(new_n772), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n775), .A2(new_n738), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n774), .B(new_n838), .C1(G283), .C2(new_n749), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n736), .A2(G107), .B1(G311), .B2(new_n746), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n837), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n732), .B1(new_n835), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n731), .A2(new_n728), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n822), .B(new_n842), .C1(new_n364), .C2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n818), .B2(new_n729), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n821), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(G384));
  INV_X1    g0647(.A(KEYINPUT35), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n482), .A2(new_n848), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n509), .B(new_n215), .C1(new_n482), .C2(new_n848), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n849), .B1(new_n851), .B2(KEYINPUT98), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(KEYINPUT98), .B2(new_n851), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT36), .Z(new_n854));
  OAI211_X1 g0654(.A(new_n793), .B(G77), .C1(new_n247), .C2(new_n220), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n218), .A2(G68), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n206), .B(G13), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(G330), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n707), .A2(new_n716), .A3(KEYINPUT31), .A4(new_n656), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n719), .A2(new_n720), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n445), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n862), .B(KEYINPUT101), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n861), .A2(new_n818), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n343), .A2(new_n657), .ZN(new_n865));
  AOI221_X4 g0665(.A(new_n865), .B1(new_n344), .B2(new_n330), .C1(new_n619), .C2(new_n356), .ZN(new_n866));
  INV_X1    g0666(.A(new_n865), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(new_n620), .B2(new_n345), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n864), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT99), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n435), .A2(new_n423), .A3(new_n302), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(G169), .B2(new_n425), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n391), .A2(new_n400), .A3(new_n402), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n404), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n875), .A2(new_n337), .A3(new_n403), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n873), .B1(new_n876), .B2(new_n413), .ZN(new_n877));
  INV_X1    g0677(.A(new_n438), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n871), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n265), .A2(new_n251), .ZN(new_n880));
  INV_X1    g0680(.A(new_n412), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n403), .A2(new_n337), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n882), .B1(new_n883), .B2(new_n875), .ZN(new_n884));
  OAI211_X1 g0684(.A(KEYINPUT99), .B(new_n438), .C1(new_n884), .C2(new_n873), .ZN(new_n885));
  OR2_X1    g0685(.A1(new_n884), .A2(new_n654), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n879), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  INV_X1    g0688(.A(new_n654), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n430), .A2(new_n431), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT37), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n432), .A2(new_n890), .A3(new_n891), .A4(new_n438), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n884), .A2(new_n654), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n444), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n893), .A2(KEYINPUT38), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n438), .A2(new_n891), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n416), .B2(new_n427), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n887), .A2(KEYINPUT37), .B1(new_n899), .B2(new_n890), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n442), .B1(KEYINPUT18), .B2(new_n432), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n886), .B1(new_n901), .B2(new_n428), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n897), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n896), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT40), .B1(new_n870), .B2(new_n904), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n893), .A2(KEYINPUT100), .A3(KEYINPUT38), .A4(new_n895), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n900), .A2(new_n902), .A3(new_n897), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT100), .ZN(new_n908));
  NOR3_X1   g0708(.A1(new_n414), .A2(new_n415), .A3(new_n654), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n624), .A2(new_n438), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT37), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n625), .A2(new_n440), .A3(new_n441), .A4(new_n626), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n911), .A2(new_n892), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n908), .B1(new_n913), .B2(KEYINPUT38), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n906), .B1(new_n907), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n358), .A2(new_n865), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n620), .A2(new_n345), .A3(new_n867), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n918), .A2(KEYINPUT40), .A3(new_n818), .A4(new_n861), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n915), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n905), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n859), .B1(new_n863), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n921), .B2(new_n863), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n630), .A2(new_n695), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(new_n629), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n815), .A2(new_n657), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n691), .B2(new_n818), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(new_n904), .A3(new_n918), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT39), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n906), .B(new_n931), .C1(new_n907), .C2(new_n914), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n330), .A2(new_n344), .A3(new_n657), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n896), .A2(new_n903), .A3(KEYINPUT39), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n932), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n627), .A2(new_n654), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n930), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n925), .B(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n923), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n206), .B2(new_n783), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n923), .A2(new_n939), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n858), .B1(new_n941), .B2(new_n942), .ZN(G367));
  OAI21_X1  g0743(.A(new_n798), .B1(new_n210), .B2(new_n362), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n791), .B2(new_n237), .ZN(new_n945));
  OAI22_X1  g0745(.A1(new_n735), .A2(new_n247), .B1(new_n761), .B2(new_n218), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n287), .B(new_n946), .C1(G150), .C2(new_n768), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n772), .A2(G77), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n947), .B(new_n948), .C1(new_n826), .C2(new_n745), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n764), .A2(G143), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n950), .B1(new_n757), .B2(new_n220), .C1(new_n750), .C2(new_n395), .ZN(new_n951));
  OR2_X1    g0751(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n952));
  NAND2_X1  g0752(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n952), .B(new_n953), .C1(new_n735), .C2(new_n509), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n749), .A2(G294), .B1(new_n764), .B2(G311), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n954), .B(new_n955), .C1(new_n203), .C2(new_n757), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n736), .A2(KEYINPUT46), .A3(G116), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n746), .A2(G317), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n287), .B1(new_n753), .B2(new_n738), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n959), .B1(G283), .B2(new_n823), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n772), .A2(G97), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n957), .A2(new_n958), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n949), .A2(new_n951), .B1(new_n956), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT47), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n822), .B(new_n945), .C1(new_n964), .C2(new_n731), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n538), .A2(new_n656), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n632), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(new_n541), .B2(new_n966), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n797), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n668), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n662), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n666), .B2(new_n971), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(new_n661), .ZN(new_n974));
  NAND3_X1  g0774(.A1(new_n695), .A2(new_n974), .A3(new_n725), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(KEYINPUT105), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT105), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n695), .A2(new_n974), .A3(new_n977), .A4(new_n725), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT45), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n497), .B(new_n500), .C1(new_n499), .C2(new_n669), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n637), .A2(new_n478), .A3(new_n670), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n979), .B1(new_n983), .B2(new_n671), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n672), .A2(new_n982), .A3(KEYINPUT45), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT44), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n672), .B2(new_n982), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n983), .A2(KEYINPUT44), .A3(new_n671), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n986), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n667), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n991), .A2(new_n992), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n993), .B1(new_n994), .B2(KEYINPUT104), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT104), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n991), .A2(new_n996), .A3(new_n992), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n976), .A2(new_n978), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n726), .ZN(new_n999));
  XOR2_X1   g0799(.A(KEYINPUT103), .B(KEYINPUT41), .Z(new_n1000));
  XNOR2_X1  g0800(.A(new_n676), .B(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n785), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n982), .A2(new_n662), .A3(new_n971), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT42), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n497), .B1(new_n980), .B2(new_n575), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n1005), .A2(new_n669), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n968), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1008), .A2(KEYINPUT43), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1008), .A2(KEYINPUT43), .ZN(new_n1010));
  OR3_X1    g0810(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  AND3_X1   g0811(.A1(new_n1007), .A2(KEYINPUT102), .A3(new_n1010), .ZN(new_n1012));
  AOI21_X1  g0812(.A(KEYINPUT102), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1014), .B1(new_n667), .B2(new_n983), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n667), .A2(new_n983), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1011), .B(new_n1016), .C1(new_n1013), .C2(new_n1012), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n970), .B1(new_n1002), .B2(new_n1018), .ZN(G387));
  NAND2_X1  g0819(.A1(new_n976), .A2(new_n978), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1020), .B(new_n676), .C1(new_n726), .C2(new_n974), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n974), .A2(new_n785), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n287), .B1(new_n769), .B2(G77), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n961), .B(new_n1023), .C1(new_n825), .C2(new_n745), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT107), .Z(new_n1025));
  AOI22_X1  g0825(.A1(G50), .A2(new_n768), .B1(new_n823), .B2(G68), .ZN(new_n1026));
  OR2_X1    g0826(.A1(new_n757), .A2(new_n362), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1026), .B(new_n1027), .C1(new_n395), .C2(new_n775), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n251), .B2(new_n749), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n371), .B1(new_n746), .B2(new_n765), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n735), .A2(new_n758), .B1(new_n757), .B2(new_n739), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT108), .Z(new_n1033));
  AOI22_X1  g0833(.A1(G317), .A2(new_n768), .B1(new_n823), .B2(G303), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n750), .B2(new_n762), .C1(new_n754), .C2(new_n775), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT48), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1033), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n1036), .B2(new_n1035), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT49), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1031), .B1(new_n509), .B2(new_n742), .C1(new_n1038), .C2(new_n1039), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1030), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n732), .B1(new_n1042), .B2(KEYINPUT109), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(KEYINPUT109), .B2(new_n1042), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n234), .A2(G45), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n359), .A2(new_n218), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT50), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n678), .B(new_n272), .C1(new_n220), .C2(new_n364), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1045), .B(new_n791), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(G107), .B2(new_n210), .C1(new_n678), .C2(new_n787), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n822), .B1(new_n1050), .B2(new_n798), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n797), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1044), .B(new_n1051), .C1(new_n666), .C2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1021), .A2(new_n1022), .A3(new_n1053), .ZN(G393));
  INV_X1    g0854(.A(new_n993), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1055), .A2(new_n994), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1056), .B1(new_n976), .B2(new_n978), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n1057), .A2(KEYINPUT111), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n998), .A2(new_n676), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1057), .A2(KEYINPUT111), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1058), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n983), .A2(new_n797), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n798), .B1(new_n202), .B2(new_n210), .C1(new_n792), .C2(new_n244), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n786), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n757), .A2(new_n364), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n371), .B1(new_n220), .B2(new_n735), .C1(new_n360), .C2(new_n761), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(G50), .C2(new_n749), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n775), .A2(new_n825), .B1(new_n753), .B2(new_n395), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT51), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G87), .A2(new_n772), .B1(new_n746), .B2(G143), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1067), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT110), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n768), .A2(G311), .B1(G317), .B2(new_n764), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT52), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n287), .B1(new_n761), .B2(new_n758), .C1(new_n739), .C2(new_n735), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n750), .A2(new_n738), .B1(new_n757), .B2(new_n509), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n203), .A2(new_n742), .B1(new_n745), .B2(new_n754), .ZN(new_n1078));
  OR4_X1    g0878(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1073), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1064), .B1(new_n1081), .B2(new_n731), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1056), .A2(new_n785), .B1(new_n1062), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(KEYINPUT112), .B1(new_n1061), .B2(new_n1083), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n676), .B(new_n998), .C1(new_n1057), .C2(KEYINPUT111), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT111), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1086), .B(new_n1056), .C1(new_n976), .C2(new_n978), .ZN(new_n1087));
  OAI211_X1 g0887(.A(KEYINPUT112), .B(new_n1083), .C1(new_n1085), .C2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1084), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(G390));
  NOR3_X1   g0891(.A1(new_n864), .A2(new_n869), .A3(new_n859), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n670), .B(new_n817), .C1(new_n689), .C2(new_n690), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n918), .B1(new_n1093), .B2(new_n927), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n1094), .A2(new_n933), .B1(new_n932), .B2(new_n935), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n812), .A2(new_n816), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n693), .A2(new_n657), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n869), .B1(new_n1097), .B2(new_n926), .ZN(new_n1098));
  NOR3_X1   g0898(.A1(new_n1098), .A2(new_n915), .A3(new_n934), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1092), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1100));
  OR3_X1    g0900(.A1(new_n1098), .A2(new_n915), .A3(new_n934), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n933), .B1(new_n928), .B2(new_n869), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n932), .A2(new_n935), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n818), .B(new_n918), .C1(new_n723), .C2(new_n724), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1101), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1100), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n785), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n843), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n786), .B1(new_n251), .B2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT54), .B(G143), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT115), .Z(new_n1112));
  AOI22_X1  g0912(.A1(new_n1112), .A2(new_n823), .B1(new_n772), .B2(G50), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n746), .A2(G125), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n749), .A2(G137), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n287), .B1(new_n768), .B2(G132), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n735), .A2(new_n825), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT53), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1118), .A2(new_n1119), .B1(G159), .B2(new_n832), .ZN(new_n1120));
  INV_X1    g0920(.A(G128), .ZN(new_n1121));
  OAI221_X1 g0921(.A(new_n1120), .B1(new_n1119), .B2(new_n1118), .C1(new_n1121), .C2(new_n775), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n287), .B1(new_n761), .B2(new_n202), .C1(new_n509), .C2(new_n753), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1123), .A2(new_n831), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n736), .A2(G87), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1124), .B(new_n1125), .C1(new_n758), .C2(new_n745), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1065), .B1(new_n764), .B2(G283), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1127), .B1(new_n203), .B2(new_n750), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n1117), .A2(new_n1122), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1110), .B1(new_n1129), .B2(new_n731), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1103), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n729), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1108), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1105), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n869), .B1(new_n864), .B2(new_n859), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1136), .A2(new_n926), .A3(new_n1097), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n818), .B1(new_n723), .B2(new_n724), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1092), .B1(new_n1140), .B2(new_n869), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT113), .ZN(new_n1142));
  NOR3_X1   g0942(.A1(new_n1141), .A2(new_n1142), .A3(new_n928), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1092), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n722), .A2(G330), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT88), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n722), .A2(KEYINPUT88), .A3(G330), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n817), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1144), .B1(new_n1149), .B2(new_n918), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT113), .B1(new_n1150), .B2(new_n929), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1139), .B1(new_n1143), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n445), .A2(G330), .A3(new_n861), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n924), .A2(new_n629), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1100), .A2(new_n1106), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n677), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1152), .A2(new_n1154), .A3(new_n1107), .ZN(new_n1158));
  AOI21_X1  g0958(.A(KEYINPUT114), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1142), .B1(new_n1141), .B2(new_n928), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n918), .B1(new_n1161), .B2(new_n818), .ZN(new_n1162));
  OAI211_X1 g0962(.A(KEYINPUT113), .B(new_n929), .C1(new_n1162), .C2(new_n1092), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1138), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n924), .A2(new_n629), .A3(new_n1153), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1156), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1158), .A2(new_n1166), .A3(KEYINPUT114), .A4(new_n676), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1134), .B1(new_n1159), .B2(new_n1168), .ZN(G378));
  INV_X1    g0969(.A(KEYINPUT57), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1165), .B1(new_n1152), .B2(new_n1107), .ZN(new_n1171));
  XOR2_X1   g0971(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n301), .B2(new_n306), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n889), .B1(new_n259), .B2(new_n267), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1176), .B(KEYINPUT118), .Z(new_n1177));
  NAND3_X1  g0977(.A1(new_n301), .A2(new_n306), .A3(new_n1173), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1175), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1177), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n305), .B(new_n1172), .C1(new_n298), .C2(new_n300), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1180), .B1(new_n1174), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(new_n921), .B2(G330), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT40), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n896), .A2(new_n903), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n918), .A2(new_n818), .A3(new_n861), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1185), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n911), .A2(new_n892), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n912), .A2(new_n909), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(KEYINPUT100), .B1(new_n1191), .B2(new_n897), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n896), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n870), .A2(new_n1193), .A3(KEYINPUT40), .A4(new_n906), .ZN(new_n1194));
  AND4_X1   g0994(.A1(G330), .A2(new_n1188), .A3(new_n1183), .A4(new_n1194), .ZN(new_n1195));
  NOR3_X1   g0995(.A1(new_n1184), .A2(new_n1195), .A3(new_n938), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n938), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1183), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1188), .A2(new_n1194), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1198), .B1(new_n1199), .B2(new_n859), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n921), .A2(G330), .A3(new_n1183), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1197), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1196), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1170), .B1(new_n1171), .B2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1154), .B1(new_n1164), .B2(new_n1156), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n938), .B1(new_n1184), .B2(new_n1195), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1200), .A2(new_n1197), .A3(new_n1201), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1206), .A2(KEYINPUT120), .A3(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT120), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1197), .A2(new_n1200), .A3(new_n1201), .A4(new_n1209), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1205), .A2(new_n1208), .A3(KEYINPUT57), .A4(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1204), .A2(new_n676), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n785), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n822), .B1(new_n218), .B2(new_n843), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n768), .A2(G107), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n1216), .A2(KEYINPUT116), .B1(new_n220), .B2(new_n757), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n371), .A2(G41), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n364), .B2(new_n735), .C1(new_n362), .C2(new_n761), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n247), .A2(new_n742), .B1(new_n745), .B2(new_n739), .ZN(new_n1220));
  NOR3_X1   g1020(.A1(new_n1217), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1216), .A2(KEYINPUT116), .B1(new_n749), .B2(G97), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1221), .B(new_n1222), .C1(new_n509), .C2(new_n775), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT58), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n753), .A2(new_n1121), .B1(new_n761), .B2(new_n826), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G150), .B2(new_n832), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n749), .A2(G132), .B1(new_n764), .B2(G125), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1112), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1226), .B(new_n1227), .C1(new_n1228), .C2(new_n735), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1229), .A2(KEYINPUT59), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(KEYINPUT59), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n772), .A2(G159), .ZN(new_n1232));
  AOI211_X1 g1032(.A(G33), .B(G41), .C1(new_n746), .C2(G124), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1218), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1235), .B(new_n218), .C1(G33), .C2(G41), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1224), .A2(new_n1234), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1238), .A2(KEYINPUT117), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n731), .B1(new_n1238), .B2(KEYINPUT117), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n1215), .B1(new_n1239), .B2(new_n1240), .C1(new_n1183), .C2(new_n729), .ZN(new_n1241));
  XOR2_X1   g1041(.A(new_n1241), .B(KEYINPUT119), .Z(new_n1242));
  NAND2_X1  g1042(.A1(new_n1214), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1212), .A2(new_n1244), .ZN(G375));
  OAI22_X1  g1045(.A1(new_n1228), .A2(new_n750), .B1(new_n1121), .B2(new_n745), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n737), .A2(new_n395), .B1(new_n247), .B2(new_n742), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n287), .B1(new_n768), .B2(G137), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n832), .A2(G50), .B1(G132), .B2(new_n764), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1248), .B(new_n1249), .C1(new_n825), .C2(new_n761), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1246), .A2(new_n1247), .A3(new_n1250), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n737), .A2(new_n202), .B1(new_n738), .B2(new_n745), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n371), .B1(new_n823), .B2(G107), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n948), .B(new_n1253), .C1(new_n739), .C2(new_n753), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n1027), .B1(new_n750), .B2(new_n509), .C1(new_n758), .C2(new_n775), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1252), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n731), .B1(new_n1251), .B2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n822), .B1(new_n220), .B2(new_n843), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1257), .B(new_n1258), .C1(new_n918), .C2(new_n729), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1259), .B1(new_n1164), .B2(new_n784), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT121), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT121), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1262), .B(new_n1259), .C1(new_n1164), .C2(new_n784), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1155), .A2(new_n1001), .A3(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(G381));
  NAND3_X1  g1067(.A1(new_n1158), .A2(new_n1166), .A3(new_n676), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1134), .ZN(new_n1269));
  OR2_X1    g1069(.A1(G393), .A2(G396), .ZN(new_n1270));
  NOR4_X1   g1070(.A1(G381), .A2(new_n1269), .A3(new_n1270), .A4(G384), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n999), .A2(new_n1001), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n784), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1018), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(new_n1273), .A2(new_n1274), .B1(new_n969), .B2(new_n965), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1205), .A2(new_n1213), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n677), .B1(new_n1276), .B2(new_n1170), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1243), .B1(new_n1277), .B2(new_n1211), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1271), .A2(new_n1275), .A3(new_n1090), .A4(new_n1278), .ZN(G407));
  INV_X1    g1079(.A(new_n1269), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1278), .A2(new_n655), .A3(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(G407), .A2(G213), .A3(new_n1281), .ZN(G409));
  NAND2_X1  g1082(.A1(new_n655), .A2(G213), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT114), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1268), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1133), .B1(new_n1285), .B2(new_n1167), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(G375), .A2(new_n1286), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1205), .A2(new_n1001), .A3(new_n1213), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1208), .A2(new_n785), .A3(new_n1210), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1241), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1288), .B1(new_n1290), .B2(KEYINPUT122), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT122), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1289), .A2(new_n1292), .A3(new_n1241), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1269), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1283), .B1(new_n1287), .B2(new_n1294), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n677), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT60), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1164), .A2(new_n1297), .A3(new_n1165), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1297), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1296), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  AND3_X1   g1100(.A1(new_n1264), .A2(new_n1300), .A3(G384), .ZN(new_n1301));
  AOI21_X1  g1101(.A(G384), .B1(new_n1264), .B2(new_n1300), .ZN(new_n1302));
  INV_X1    g1102(.A(G2897), .ZN(new_n1303));
  OAI22_X1  g1103(.A1(new_n1301), .A2(new_n1302), .B1(new_n1303), .B2(new_n1283), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1264), .A2(new_n1300), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n846), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1264), .A2(new_n1300), .A3(G384), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1283), .A2(new_n1303), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1304), .A2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT61), .B1(new_n1295), .B2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(G378), .A2(new_n1278), .ZN(new_n1312));
  AND2_X1   g1112(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1312), .B1(new_n1313), .B2(new_n1269), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT62), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1314), .A2(new_n1315), .A3(new_n1316), .A4(new_n1283), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1316), .B(new_n1283), .C1(new_n1287), .C2(new_n1294), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(KEYINPUT62), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1311), .A2(new_n1317), .A3(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1275), .B1(new_n1084), .B2(new_n1089), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1083), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT112), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1324), .A2(G387), .A3(new_n1088), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1321), .A2(new_n1325), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(G393), .A2(G396), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1326), .A2(new_n1270), .A3(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT125), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1321), .A2(new_n1329), .ZN(new_n1330));
  OAI211_X1 g1130(.A(new_n1275), .B(KEYINPUT125), .C1(new_n1084), .C2(new_n1089), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT124), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1325), .A2(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1330), .A2(new_n1331), .A3(new_n1333), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1324), .A2(G387), .A3(KEYINPUT124), .A4(new_n1088), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1270), .A2(new_n1327), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1328), .B1(new_n1334), .B2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT123), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1314), .A2(new_n1339), .A3(new_n1283), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1295), .A2(KEYINPUT123), .ZN(new_n1341));
  AOI22_X1  g1141(.A1(new_n1340), .A2(new_n1341), .B1(new_n1309), .B2(new_n1304), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT63), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1318), .A2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT61), .ZN(new_n1345));
  NOR3_X1   g1145(.A1(new_n1301), .A2(new_n1302), .A3(new_n1343), .ZN(new_n1346));
  OAI211_X1 g1146(.A(new_n1346), .B(new_n1283), .C1(new_n1287), .C2(new_n1294), .ZN(new_n1347));
  NAND4_X1  g1147(.A1(new_n1344), .A2(new_n1345), .A3(new_n1338), .A4(new_n1347), .ZN(new_n1348));
  OAI22_X1  g1148(.A1(new_n1320), .A2(new_n1338), .B1(new_n1342), .B2(new_n1348), .ZN(G405));
  INV_X1    g1149(.A(KEYINPUT127), .ZN(new_n1350));
  AND2_X1   g1150(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1351), .A2(new_n1331), .A3(new_n1330), .A4(new_n1333), .ZN(new_n1352));
  AND2_X1   g1152(.A1(new_n1352), .A2(new_n1328), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1269), .B1(new_n1212), .B2(new_n1244), .ZN(new_n1354));
  NOR3_X1   g1154(.A1(new_n1287), .A2(new_n1316), .A3(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(G375), .A2(new_n1280), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1356), .B1(new_n1312), .B2(new_n1357), .ZN(new_n1358));
  NOR2_X1   g1158(.A1(new_n1355), .A2(new_n1358), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1350), .B1(new_n1353), .B2(new_n1359), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1316), .B1(new_n1287), .B2(new_n1354), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1312), .A2(new_n1356), .A3(new_n1357), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1363), .A2(new_n1338), .A3(KEYINPUT127), .ZN(new_n1364));
  INV_X1    g1164(.A(KEYINPUT126), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1353), .A2(new_n1359), .A3(new_n1365), .ZN(new_n1366));
  OAI21_X1  g1166(.A(KEYINPUT126), .B1(new_n1363), .B2(new_n1338), .ZN(new_n1367));
  AOI22_X1  g1167(.A1(new_n1360), .A2(new_n1364), .B1(new_n1366), .B2(new_n1367), .ZN(G402));
endmodule


