//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  INV_X1    g0013(.A(G107), .ZN(new_n214));
  INV_X1    g0014(.A(G264), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G58), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR4_X1   g0025(.A1(new_n216), .A2(new_n219), .A3(new_n222), .A4(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(KEYINPUT64), .B(G68), .Z(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G238), .ZN(new_n228));
  AOI22_X1  g0028(.A1(new_n226), .A2(new_n228), .B1(G1), .B2(G20), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT1), .Z(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n231), .A2(new_n207), .ZN(new_n232));
  INV_X1    g0032(.A(new_n201), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(G50), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  AOI211_X1 g0035(.A(new_n210), .B(new_n230), .C1(new_n232), .C2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  INV_X1    g0045(.A(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(KEYINPUT65), .B(G107), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G68), .B(G77), .Z(new_n250));
  XOR2_X1   g0050(.A(G50), .B(G58), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G41), .ZN(new_n255));
  OAI211_X1 g0055(.A(G1), .B(G13), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n257));
  AND3_X1   g0057(.A1(new_n256), .A2(G238), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n261));
  NAND4_X1  g0061(.A1(new_n260), .A2(new_n261), .A3(G232), .A4(G1698), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT70), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT3), .B(G33), .ZN(new_n265));
  NAND4_X1  g0065(.A1(new_n265), .A2(KEYINPUT70), .A3(G232), .A4(G1698), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(G226), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G97), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n264), .A2(new_n266), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n256), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n258), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT13), .ZN(new_n273));
  INV_X1    g0073(.A(G274), .ZN(new_n274));
  OR2_X1    g0074(.A1(new_n257), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT66), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n275), .B(new_n276), .ZN(new_n277));
  AND3_X1   g0077(.A1(new_n272), .A2(new_n273), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n273), .B1(new_n272), .B2(new_n277), .ZN(new_n279));
  OAI21_X1  g0079(.A(G169), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT14), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n272), .A2(new_n277), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT13), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n272), .A2(new_n273), .A3(new_n277), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n283), .A2(G179), .A3(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT14), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n286), .B(G169), .C1(new_n278), .C2(new_n279), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n281), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n231), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(G1), .B2(new_n207), .ZN(new_n292));
  INV_X1    g0092(.A(G68), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT72), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n296));
  OR3_X1    g0096(.A1(new_n296), .A2(KEYINPUT12), .A3(G68), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n297), .A2(KEYINPUT73), .ZN(new_n298));
  OAI21_X1  g0098(.A(KEYINPUT12), .B1(new_n227), .B2(new_n296), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(KEYINPUT73), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(G20), .A2(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G50), .ZN(new_n303));
  XOR2_X1   g0103(.A(new_n303), .B(KEYINPUT71), .Z(new_n304));
  NAND2_X1  g0104(.A1(new_n207), .A2(G33), .ZN(new_n305));
  OAI221_X1 g0105(.A(new_n304), .B1(new_n207), .B2(new_n227), .C1(new_n220), .C2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT11), .ZN(new_n307));
  AND3_X1   g0107(.A1(new_n306), .A2(new_n307), .A3(new_n290), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n307), .B1(new_n306), .B2(new_n290), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n295), .B(new_n301), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n288), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n265), .A2(G238), .A3(G1698), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(new_n214), .B2(new_n265), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n260), .A2(new_n261), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n314), .A2(new_n224), .A3(G1698), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n271), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n256), .A2(new_n257), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n316), .B(new_n277), .C1(new_n221), .C2(new_n317), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n318), .A2(G179), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G20), .A2(G77), .ZN(new_n320));
  XOR2_X1   g0120(.A(KEYINPUT15), .B(G87), .Z(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n302), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT8), .B(G58), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n320), .B1(new_n322), .B2(new_n305), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n296), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n325), .A2(new_n290), .B1(new_n220), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n327), .B1(new_n220), .B2(new_n292), .ZN(new_n328));
  INV_X1    g0128(.A(G169), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n318), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n319), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n311), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n328), .B1(G200), .B2(new_n318), .ZN(new_n333));
  INV_X1    g0133(.A(G190), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n333), .B1(new_n334), .B2(new_n318), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT16), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT64), .B(G68), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT74), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n254), .ZN(new_n339));
  NAND2_X1  g0139(.A1(KEYINPUT74), .A2(G33), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT3), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n261), .ZN(new_n342));
  OAI211_X1 g0142(.A(KEYINPUT7), .B(new_n207), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT7), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n344), .B1(new_n265), .B2(G20), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n337), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n302), .A2(G159), .ZN(new_n347));
  XOR2_X1   g0147(.A(KEYINPUT67), .B(G58), .Z(new_n348));
  AOI21_X1  g0148(.A(new_n201), .B1(new_n227), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n347), .B1(new_n349), .B2(new_n207), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n336), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT67), .B(G58), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n233), .B1(new_n337), .B2(new_n352), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(G20), .B1(G159), .B2(new_n302), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n339), .A2(KEYINPUT3), .A3(new_n340), .ZN(new_n355));
  AOI21_X1  g0155(.A(G20), .B1(new_n355), .B2(new_n260), .ZN(new_n356));
  OAI21_X1  g0156(.A(G68), .B1(new_n356), .B2(new_n344), .ZN(new_n357));
  AOI211_X1 g0157(.A(KEYINPUT7), .B(G20), .C1(new_n355), .C2(new_n260), .ZN(new_n358));
  OAI211_X1 g0158(.A(KEYINPUT16), .B(new_n354), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n351), .A2(new_n290), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT8), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n223), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n362), .B1(new_n352), .B2(new_n361), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n326), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n363), .B2(new_n292), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G200), .ZN(new_n368));
  XNOR2_X1  g0168(.A(new_n275), .B(KEYINPUT66), .ZN(new_n369));
  INV_X1    g0169(.A(new_n260), .ZN(new_n370));
  AND2_X1   g0170(.A1(KEYINPUT74), .A2(G33), .ZN(new_n371));
  NOR2_X1   g0171(.A1(KEYINPUT74), .A2(G33), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n370), .B1(new_n373), .B2(KEYINPUT3), .ZN(new_n374));
  AND2_X1   g0174(.A1(G226), .A2(G1698), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n374), .A2(new_n375), .B1(G33), .B2(G87), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT75), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n374), .A2(new_n377), .A3(G223), .A4(new_n267), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n355), .A2(G223), .A3(new_n267), .A4(new_n260), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT75), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n376), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n369), .B1(new_n381), .B2(new_n271), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n317), .A2(new_n224), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n368), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n367), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT17), .ZN(new_n387));
  OR2_X1    g0187(.A1(new_n387), .A2(KEYINPUT76), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n382), .A2(G190), .A3(new_n384), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(KEYINPUT76), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n386), .A2(new_n388), .A3(new_n389), .A4(new_n390), .ZN(new_n391));
  AOI211_X1 g0191(.A(new_n369), .B(new_n383), .C1(new_n381), .C2(new_n271), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n366), .B(new_n360), .C1(new_n392), .C2(new_n368), .ZN(new_n393));
  INV_X1    g0193(.A(new_n389), .ZN(new_n394));
  OAI211_X1 g0194(.A(KEYINPUT76), .B(new_n387), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n381), .A2(new_n271), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n396), .A2(G179), .A3(new_n277), .A4(new_n384), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n392), .B2(new_n329), .ZN(new_n398));
  AND3_X1   g0198(.A1(new_n398), .A2(KEYINPUT18), .A3(new_n367), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT18), .B1(new_n398), .B2(new_n367), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n391), .B(new_n395), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n335), .B1(new_n402), .B2(KEYINPUT77), .ZN(new_n403));
  AOI211_X1 g0203(.A(new_n332), .B(new_n403), .C1(KEYINPUT77), .C2(new_n402), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n326), .A2(G50), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n405), .B1(new_n292), .B2(G50), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT68), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n203), .A2(G20), .ZN(new_n408));
  INV_X1    g0208(.A(G150), .ZN(new_n409));
  OAI221_X1 g0209(.A(new_n408), .B1(new_n409), .B2(new_n323), .C1(new_n363), .C2(new_n305), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n290), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT9), .ZN(new_n413));
  INV_X1    g0213(.A(new_n317), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G226), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n314), .A2(new_n220), .ZN(new_n416));
  MUX2_X1   g0216(.A(G222), .B(G223), .S(G1698), .Z(new_n417));
  OAI211_X1 g0217(.A(new_n416), .B(new_n271), .C1(new_n314), .C2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n277), .A2(new_n415), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G200), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n407), .A2(new_n411), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT9), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n419), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G190), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n413), .A2(new_n420), .A3(new_n423), .A4(new_n425), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT10), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n424), .A2(G169), .ZN(new_n428));
  OR3_X1    g0228(.A1(new_n412), .A2(new_n428), .A3(KEYINPUT69), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT69), .B1(new_n412), .B2(new_n428), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n429), .B(new_n430), .C1(G179), .C2(new_n419), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n283), .A2(G190), .A3(new_n284), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n283), .A2(new_n284), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n310), .B1(G200), .B2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n432), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n404), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT22), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(new_n212), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n355), .A2(new_n207), .A3(new_n260), .A4(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n260), .A2(new_n261), .A3(new_n207), .A4(G87), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n439), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n214), .A2(G20), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT23), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n444), .B(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n339), .A2(new_n340), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(new_n207), .A3(G116), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n441), .A2(new_n443), .A3(new_n446), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT81), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n246), .B1(new_n339), .B2(new_n340), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n439), .A2(new_n442), .B1(new_n451), .B2(new_n207), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT81), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n452), .A2(new_n453), .A3(new_n441), .A4(new_n446), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT24), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n450), .A2(new_n454), .A3(KEYINPUT24), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(new_n290), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n206), .A2(G33), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n291), .A2(new_n296), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G107), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n326), .B(new_n214), .C1(KEYINPUT82), .C2(KEYINPUT25), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT82), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT25), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n464), .B(new_n465), .C1(new_n296), .C2(G107), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n463), .B(new_n466), .C1(new_n464), .C2(new_n465), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n459), .A2(new_n462), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n213), .A2(new_n267), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n218), .A2(G1698), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n355), .A2(new_n260), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n447), .A2(G294), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n256), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G45), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(G1), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n255), .A2(KEYINPUT5), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT5), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G41), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n475), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(new_n274), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n256), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(new_n215), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n473), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(G169), .ZN(new_n484));
  INV_X1    g0284(.A(G179), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n484), .B1(new_n485), .B2(new_n483), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n468), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n483), .A2(new_n334), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(G200), .B2(new_n483), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n459), .A2(new_n489), .A3(new_n462), .A4(new_n467), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  XNOR2_X1  g0291(.A(G97), .B(G107), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT6), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NOR3_X1   g0294(.A1(new_n493), .A2(new_n217), .A3(G107), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n497), .A2(G20), .B1(G77), .B2(new_n302), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT7), .B1(new_n314), .B2(new_n207), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n259), .B1(new_n371), .B2(new_n372), .ZN(new_n500));
  AOI21_X1  g0300(.A(G20), .B1(new_n500), .B2(new_n261), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n499), .B1(new_n501), .B2(KEYINPUT7), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n498), .B1(new_n502), .B2(new_n214), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n503), .A2(new_n290), .B1(new_n217), .B2(new_n326), .ZN(new_n504));
  INV_X1    g0304(.A(new_n480), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n481), .A2(new_n218), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n260), .A2(new_n261), .A3(G250), .A4(G1698), .ZN(new_n508));
  AND2_X1   g0308(.A1(KEYINPUT4), .A2(G244), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n260), .A2(new_n261), .A3(new_n509), .A4(new_n267), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G283), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n508), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT4), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n355), .A2(G244), .A3(new_n267), .A4(new_n260), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n505), .B(new_n507), .C1(new_n515), .C2(new_n256), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G200), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n461), .A2(G97), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n514), .A2(new_n513), .ZN(new_n519));
  AND3_X1   g0319(.A1(new_n508), .A2(new_n510), .A3(new_n511), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n271), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n522), .A2(G190), .A3(new_n505), .A4(new_n507), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n504), .A2(new_n517), .A3(new_n518), .A4(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n326), .A2(new_n217), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n495), .B1(new_n493), .B2(new_n492), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n526), .A2(new_n207), .B1(new_n220), .B2(new_n323), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n343), .A2(new_n345), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n527), .B1(G107), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n525), .B(new_n518), .C1(new_n529), .C2(new_n291), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n256), .B1(new_n519), .B2(new_n520), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n531), .A2(new_n506), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n532), .A2(new_n485), .A3(new_n505), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n516), .A2(new_n329), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n530), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n524), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(G238), .A2(G1698), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n537), .B1(new_n221), .B2(G1698), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(new_n355), .A3(new_n260), .ZN(new_n539));
  INV_X1    g0339(.A(new_n451), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n271), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n475), .A2(G274), .ZN(new_n543));
  INV_X1    g0343(.A(new_n475), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n256), .A2(new_n544), .A3(G250), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT78), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT78), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n256), .A2(new_n544), .A3(new_n547), .A4(G250), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n542), .A2(new_n543), .A3(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n355), .A2(new_n207), .A3(G68), .A4(new_n260), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT19), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n207), .B1(new_n269), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n212), .A2(new_n217), .A3(new_n214), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n553), .A2(new_n554), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n551), .A2(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n557), .A2(new_n290), .B1(new_n326), .B2(new_n322), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n461), .A2(new_n321), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n550), .A2(new_n329), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n541), .A2(new_n271), .B1(G274), .B2(new_n475), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n561), .A2(new_n485), .A3(new_n549), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n550), .A2(G200), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n561), .A2(G190), .A3(new_n549), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n461), .A2(G87), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n564), .A2(new_n558), .A3(new_n565), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(KEYINPUT79), .B1(new_n536), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n557), .A2(new_n290), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n322), .A2(new_n326), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n570), .A2(new_n571), .A3(new_n566), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(G200), .B2(new_n550), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n565), .A2(new_n573), .B1(new_n560), .B2(new_n562), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT79), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n574), .A2(new_n575), .A3(new_n524), .A4(new_n535), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n296), .A2(G116), .ZN(new_n577));
  AND4_X1   g0377(.A1(G116), .A2(new_n291), .A3(new_n296), .A4(new_n460), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n511), .B(new_n207), .C1(G33), .C2(new_n217), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT80), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n289), .A2(new_n231), .B1(G20), .B2(new_n246), .ZN(new_n582));
  AOI21_X1  g0382(.A(G20), .B1(new_n254), .B2(G97), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(KEYINPUT80), .A3(new_n511), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT20), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n581), .A2(new_n584), .A3(KEYINPUT20), .A4(new_n582), .ZN(new_n588));
  AOI211_X1 g0388(.A(new_n577), .B(new_n578), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n218), .A2(new_n267), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n215), .A2(G1698), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n355), .A2(new_n260), .A3(new_n590), .A4(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n314), .A2(G303), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n271), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n479), .A2(G270), .A3(new_n256), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n595), .A2(G179), .A3(new_n505), .A4(new_n596), .ZN(new_n597));
  OR2_X1    g0397(.A1(new_n589), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n595), .A2(new_n505), .A3(new_n596), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G200), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n600), .B(new_n589), .C1(new_n334), .C2(new_n599), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n577), .B1(new_n587), .B2(new_n588), .ZN(new_n602));
  INV_X1    g0402(.A(new_n578), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n604), .A2(KEYINPUT21), .A3(G169), .A4(new_n599), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT21), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n599), .A2(G169), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n606), .B1(new_n607), .B2(new_n589), .ZN(new_n608));
  AND4_X1   g0408(.A1(new_n598), .A2(new_n601), .A3(new_n605), .A4(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n576), .A2(new_n609), .ZN(new_n610));
  AND4_X1   g0410(.A1(new_n438), .A2(new_n491), .A3(new_n569), .A4(new_n610), .ZN(G372));
  AND4_X1   g0411(.A1(new_n490), .A2(new_n567), .A3(new_n535), .A4(new_n524), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n608), .A2(new_n605), .A3(new_n598), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n487), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT26), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n568), .B2(new_n535), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n530), .A2(new_n533), .A3(new_n534), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n619), .A2(new_n574), .A3(KEYINPUT26), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n618), .A2(new_n620), .B1(new_n562), .B2(new_n560), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n438), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g0423(.A(new_n623), .B(KEYINPUT83), .Z(new_n624));
  INV_X1    g0424(.A(new_n431), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n311), .A2(new_n433), .A3(new_n435), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n391), .A2(new_n395), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(new_n627), .A3(new_n332), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(new_n400), .B2(new_n399), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n625), .B1(new_n629), .B2(new_n427), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n624), .A2(new_n630), .ZN(G369));
  INV_X1    g0431(.A(G343), .ZN(new_n632));
  XOR2_X1   g0432(.A(KEYINPUT84), .B(KEYINPUT27), .Z(new_n633));
  INV_X1    g0433(.A(G13), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n634), .A2(G1), .A3(G20), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n633), .A2(new_n635), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n636), .A2(G213), .A3(new_n637), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n589), .A2(new_n632), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n613), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n614), .A2(new_n601), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n640), .B1(new_n641), .B2(new_n639), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(KEYINPUT85), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT85), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n644), .B(new_n640), .C1(new_n641), .C2(new_n639), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(G330), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n638), .A2(new_n632), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n468), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n487), .A2(new_n649), .A3(new_n490), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n468), .A2(new_n486), .A3(new_n648), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT86), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n647), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n614), .A2(new_n648), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n653), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g0458(.A(new_n648), .B(KEYINPUT87), .Z(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n468), .A2(new_n660), .A3(new_n486), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n656), .A2(new_n662), .ZN(G399));
  INV_X1    g0463(.A(new_n208), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(G41), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n554), .A2(G116), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G1), .A3(new_n667), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n668), .A2(KEYINPUT88), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(KEYINPUT88), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n669), .B(new_n670), .C1(new_n234), .C2(new_n666), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT28), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n610), .A2(new_n491), .A3(new_n569), .A4(new_n660), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n483), .B1(new_n532), .B2(new_n505), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n674), .A2(new_n485), .A3(new_n550), .A4(new_n599), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT30), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n550), .A2(new_n531), .A3(new_n506), .ZN(new_n677));
  INV_X1    g0477(.A(new_n482), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n471), .A2(new_n472), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n505), .B(new_n678), .C1(new_n679), .C2(new_n256), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n597), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n676), .B1(new_n677), .B2(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n522), .A2(new_n561), .A3(new_n549), .A4(new_n507), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n473), .A2(new_n482), .ZN(new_n684));
  INV_X1    g0484(.A(new_n596), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n685), .B1(new_n594), .B2(new_n271), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n684), .A2(new_n686), .A3(G179), .A4(new_n505), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n683), .A2(new_n687), .A3(KEYINPUT30), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n675), .B1(new_n682), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT89), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT89), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n675), .B(new_n691), .C1(new_n682), .C2(new_n688), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n690), .A2(new_n648), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT31), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n689), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n673), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT90), .B1(new_n697), .B2(G330), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n697), .A2(KEYINPUT90), .A3(G330), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT92), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n618), .A2(new_n620), .A3(new_n702), .ZN(new_n703));
  OAI211_X1 g0503(.A(KEYINPUT92), .B(new_n617), .C1(new_n568), .C2(new_n535), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n703), .A2(new_n563), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT93), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n615), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n487), .A2(KEYINPUT93), .A3(new_n614), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(new_n708), .A3(new_n612), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n648), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n659), .B1(new_n616), .B2(new_n621), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  XOR2_X1   g0512(.A(KEYINPUT91), .B(KEYINPUT29), .Z(new_n713));
  AOI22_X1  g0513(.A1(new_n710), .A2(KEYINPUT29), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n701), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n672), .B1(new_n715), .B2(G1), .ZN(G364));
  NOR3_X1   g0516(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n640), .B(new_n717), .C1(new_n641), .C2(new_n639), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n634), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n206), .B1(new_n719), .B2(G45), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n665), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n374), .A2(new_n664), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n724), .B1(new_n252), .B2(G45), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(G45), .B2(new_n234), .ZN(new_n726));
  INV_X1    g0526(.A(G355), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n265), .A2(new_n208), .ZN(new_n728));
  OAI221_X1 g0528(.A(new_n726), .B1(G116), .B2(new_n208), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n231), .B1(G20), .B2(new_n329), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n717), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n733), .A2(KEYINPUT95), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(KEYINPUT95), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n734), .A2(new_n334), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g0536(.A(KEYINPUT33), .B(G317), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n207), .A2(G190), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n485), .A2(G200), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n736), .A2(new_n737), .B1(G311), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G179), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n738), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G329), .ZN(new_n746));
  INV_X1    g0546(.A(G283), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n368), .A2(G179), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(new_n738), .ZN(new_n749));
  OAI211_X1 g0549(.A(new_n742), .B(new_n746), .C1(new_n747), .C2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n207), .A2(new_n334), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(new_n748), .ZN(new_n752));
  INV_X1    g0552(.A(G303), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n734), .A2(G190), .A3(new_n735), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AND2_X1   g0556(.A1(new_n756), .A2(G326), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n207), .B1(new_n743), .B2(G190), .ZN(new_n758));
  INV_X1    g0558(.A(G294), .ZN(new_n759));
  INV_X1    g0559(.A(G322), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n751), .A2(new_n739), .ZN(new_n761));
  OAI221_X1 g0561(.A(new_n314), .B1(new_n758), .B2(new_n759), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  NOR4_X1   g0562(.A1(new_n750), .A2(new_n754), .A3(new_n757), .A4(new_n762), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n740), .A2(KEYINPUT94), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n740), .A2(KEYINPUT94), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n265), .B1(new_n766), .B2(new_n220), .ZN(new_n767));
  INV_X1    g0567(.A(new_n736), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n293), .ZN(new_n769));
  INV_X1    g0569(.A(G159), .ZN(new_n770));
  OR3_X1    g0570(.A1(new_n744), .A2(KEYINPUT32), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(KEYINPUT32), .B1(new_n744), .B2(new_n770), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n771), .B(new_n772), .C1(new_n202), .C2(new_n755), .ZN(new_n773));
  INV_X1    g0573(.A(new_n752), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G87), .ZN(new_n775));
  INV_X1    g0575(.A(new_n761), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n348), .ZN(new_n777));
  INV_X1    g0577(.A(new_n749), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G107), .ZN(new_n779));
  INV_X1    g0579(.A(new_n758), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G97), .ZN(new_n781));
  NAND4_X1  g0581(.A1(new_n775), .A2(new_n777), .A3(new_n779), .A4(new_n781), .ZN(new_n782));
  NOR4_X1   g0582(.A1(new_n767), .A2(new_n769), .A3(new_n773), .A4(new_n782), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n730), .B1(new_n763), .B2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n718), .A2(new_n722), .A3(new_n732), .A4(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n722), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n647), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n646), .A2(G330), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n785), .B1(new_n787), .B2(new_n788), .ZN(G396));
  INV_X1    g0589(.A(new_n331), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n328), .A2(new_n648), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n790), .B1(new_n335), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n331), .A2(new_n648), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AND4_X1   g0594(.A1(KEYINPUT98), .A2(new_n622), .A3(new_n660), .A4(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(KEYINPUT98), .B1(new_n711), .B2(new_n794), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n794), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n797), .B1(new_n712), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n799), .A2(new_n701), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(new_n786), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n801), .A2(KEYINPUT99), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(KEYINPUT99), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n802), .B(new_n803), .C1(new_n701), .C2(new_n799), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G13), .A2(G33), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n730), .A2(new_n805), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT96), .Z(new_n807));
  AOI21_X1  g0607(.A(new_n786), .B1(new_n807), .B2(new_n220), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n798), .A2(new_n805), .B1(KEYINPUT97), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G132), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n374), .B1(new_n811), .B2(new_n744), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G137), .A2(new_n756), .B1(new_n736), .B2(G150), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n770), .B2(new_n766), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G143), .B2(new_n776), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT34), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n812), .B(new_n816), .C1(G68), .C2(new_n778), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n817), .B1(new_n202), .B2(new_n752), .C1(new_n352), .C2(new_n758), .ZN(new_n818));
  INV_X1    g0618(.A(G311), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n761), .A2(new_n759), .B1(new_n744), .B2(new_n819), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n781), .B(new_n314), .C1(new_n214), .C2(new_n752), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n820), .B(new_n821), .C1(G87), .C2(new_n778), .ZN(new_n822));
  INV_X1    g0622(.A(new_n766), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n823), .A2(G116), .B1(G303), .B2(new_n756), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n822), .B(new_n824), .C1(new_n747), .C2(new_n768), .ZN(new_n825));
  AND2_X1   g0625(.A1(new_n818), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n730), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n810), .B1(KEYINPUT97), .B2(new_n809), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n804), .A2(new_n828), .ZN(G384));
  NAND4_X1  g0629(.A1(new_n690), .A2(KEYINPUT31), .A3(new_n648), .A4(new_n692), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n673), .A2(new_n695), .A3(new_n830), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n435), .A2(new_n433), .B1(new_n310), .B2(new_n648), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT101), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n287), .A2(new_n285), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n286), .B1(new_n434), .B2(G169), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n833), .B(new_n310), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n833), .B1(new_n288), .B2(new_n310), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n832), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n310), .B(new_n648), .C1(new_n834), .C2(new_n835), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT102), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n288), .A2(KEYINPUT102), .A3(new_n310), .A4(new_n648), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  AND3_X1   g0645(.A1(new_n831), .A2(new_n845), .A3(new_n794), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT38), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n354), .B1(new_n357), .B2(new_n358), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n291), .B1(new_n848), .B2(new_n336), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n359), .B1(new_n849), .B2(KEYINPUT103), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT7), .B1(new_n374), .B2(G20), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n356), .A2(new_n344), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n851), .A2(G68), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT16), .B1(new_n853), .B2(new_n354), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT103), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n854), .A2(new_n855), .A3(new_n291), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n366), .B1(new_n850), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n638), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n397), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n329), .B1(new_n382), .B2(new_n384), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n367), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT18), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n862), .B(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n859), .B1(new_n627), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT37), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n354), .B1(new_n502), .B2(new_n337), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n291), .B1(new_n867), .B2(new_n336), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n365), .B1(new_n868), .B2(new_n359), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n396), .A2(new_n277), .A3(new_n384), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(G200), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n869), .A2(new_n871), .A3(new_n389), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n367), .A2(new_n858), .ZN(new_n873));
  AND4_X1   g0673(.A1(new_n866), .A2(new_n862), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n857), .B1(new_n398), .B2(new_n858), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n872), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n874), .B1(new_n876), .B2(KEYINPUT37), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n847), .B1(new_n865), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n398), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n855), .B1(new_n854), .B2(new_n291), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n848), .A2(new_n336), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n881), .A2(KEYINPUT103), .A3(new_n290), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n880), .A2(new_n882), .A3(new_n359), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n879), .A2(new_n638), .B1(new_n883), .B2(new_n366), .ZN(new_n884));
  INV_X1    g0684(.A(new_n872), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT37), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n862), .A2(new_n872), .A3(new_n866), .A4(new_n873), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n859), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n401), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n888), .A2(new_n890), .A3(KEYINPUT38), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n878), .A2(KEYINPUT104), .A3(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT40), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT104), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n888), .A2(new_n890), .A3(new_n894), .A4(KEYINPUT38), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n846), .A2(new_n892), .A3(new_n893), .A4(new_n895), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n888), .A2(new_n890), .A3(KEYINPUT38), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n401), .A2(new_n367), .A3(new_n858), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n862), .A2(new_n872), .A3(new_n873), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT37), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(new_n887), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n897), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n831), .A2(new_n845), .A3(new_n794), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT40), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n896), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(G330), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n404), .A2(G330), .A3(new_n436), .A4(new_n831), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n438), .A2(new_n906), .A3(new_n831), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n793), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n795), .B2(new_n796), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n913), .A2(new_n845), .A3(new_n895), .A4(new_n892), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n864), .A2(new_n858), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n837), .A2(new_n838), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n917), .A2(new_n648), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n892), .A2(KEYINPUT39), .A3(new_n895), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n903), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n919), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n916), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n911), .B(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n404), .A2(new_n436), .A3(new_n714), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(new_n630), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n925), .B(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n206), .B2(new_n719), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n526), .B(KEYINPUT100), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n246), .B1(new_n930), .B2(KEYINPUT35), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n931), .B(new_n232), .C1(KEYINPUT35), .C2(new_n930), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT36), .ZN(new_n933));
  NAND2_X1  g0733(.A1(G50), .A2(G58), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n206), .B1(new_n934), .B2(new_n293), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n220), .B1(new_n227), .B2(new_n348), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n634), .B(new_n935), .C1(new_n936), .C2(new_n202), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n929), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT105), .ZN(G367));
  INV_X1    g0739(.A(KEYINPUT42), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n659), .A2(new_n530), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(new_n535), .A3(new_n524), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n619), .A2(new_n659), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n653), .A2(new_n654), .A3(new_n657), .A4(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(KEYINPUT107), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n945), .A2(KEYINPUT107), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n940), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n948), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n950), .A2(KEYINPUT42), .A3(new_n946), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n535), .B1(new_n942), .B2(new_n487), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n660), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n949), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n572), .A2(new_n648), .ZN(new_n955));
  MUX2_X1   g0755(.A(new_n563), .B(new_n568), .S(new_n955), .Z(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT106), .Z(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n954), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n960), .B1(new_n954), .B2(new_n961), .ZN(new_n964));
  INV_X1    g0764(.A(new_n656), .ZN(new_n965));
  INV_X1    g0765(.A(new_n944), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n963), .A2(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n964), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n965), .A2(new_n966), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n968), .A2(new_n969), .A3(new_n962), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n665), .B(KEYINPUT41), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT108), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n647), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n658), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n657), .B1(new_n653), .B2(new_n654), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n647), .B(new_n973), .C1(new_n975), .C2(new_n976), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR3_X1   g0780(.A1(new_n980), .A2(new_n701), .A3(new_n714), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n658), .A2(new_n661), .A3(new_n944), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT45), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n982), .A2(new_n983), .ZN(new_n985));
  AND3_X1   g0785(.A1(new_n662), .A2(KEYINPUT44), .A3(new_n966), .ZN(new_n986));
  AOI21_X1  g0786(.A(KEYINPUT44), .B1(new_n662), .B2(new_n966), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n984), .A2(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n656), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n965), .B1(new_n986), .B2(new_n987), .C1(new_n984), .C2(new_n985), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n981), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n972), .B1(new_n991), .B2(new_n715), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n967), .B(new_n970), .C1(new_n992), .C2(new_n721), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n314), .B1(new_n774), .B2(new_n348), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n776), .A2(G150), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n745), .A2(G137), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n780), .A2(G68), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n994), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n823), .A2(G50), .B1(G143), .B2(new_n756), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n770), .B2(new_n768), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n998), .B(new_n1000), .C1(G77), .C2(new_n778), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n778), .A2(G97), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n756), .A2(G311), .B1(G303), .B2(new_n776), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n1004), .A2(KEYINPUT109), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1004), .A2(KEYINPUT109), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1002), .B1(new_n759), .B2(new_n768), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n752), .A2(new_n246), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT46), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n374), .ZN(new_n1010));
  INV_X1    g0810(.A(G317), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1010), .B1(new_n1011), .B2(new_n744), .C1(new_n766), .C2(new_n747), .ZN(new_n1012));
  NOR3_X1   g0812(.A1(new_n1007), .A2(new_n1009), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n780), .A2(G107), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1001), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT110), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT47), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n730), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n957), .A2(new_n717), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n731), .B1(new_n208), .B2(new_n322), .C1(new_n724), .C2(new_n243), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1018), .A2(new_n722), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n993), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(KEYINPUT111), .ZN(new_n1023));
  INV_X1    g0823(.A(KEYINPUT111), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n993), .A2(new_n1024), .A3(new_n1021), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(G387));
  AOI22_X1  g0827(.A1(G322), .A2(new_n756), .B1(new_n736), .B2(G311), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n753), .B2(new_n766), .C1(new_n1011), .C2(new_n761), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT48), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n747), .B2(new_n758), .C1(new_n759), .C2(new_n752), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT49), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n374), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n778), .A2(G116), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n745), .A2(G326), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n756), .A2(G159), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n780), .A2(new_n321), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n774), .A2(G77), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1038), .A2(new_n1002), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G150), .B2(new_n745), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n374), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G68), .B2(new_n741), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n202), .B2(new_n761), .C1(new_n363), .C2(new_n768), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n827), .B1(new_n1037), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n723), .B1(new_n240), .B2(new_n474), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n667), .B2(new_n728), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n324), .A2(G50), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT50), .ZN(new_n1050));
  AOI21_X1  g0850(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1050), .A2(new_n667), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1048), .A2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(G107), .B2(new_n208), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n786), .B(new_n1046), .C1(new_n731), .C2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n655), .A2(new_n717), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n980), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n1055), .A2(new_n1056), .B1(new_n1057), .B2(new_n721), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n665), .B1(new_n715), .B2(new_n1057), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1058), .B1(new_n1059), .B2(new_n981), .ZN(G393));
  INV_X1    g0860(.A(new_n981), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n989), .A2(new_n990), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n666), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1063), .A2(new_n991), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n758), .A2(new_n220), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G87), .B2(new_n778), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1066), .B(new_n374), .C1(new_n766), .C2(new_n324), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n755), .A2(new_n409), .B1(new_n770), .B2(new_n761), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT51), .Z(new_n1069));
  AOI211_X1 g0869(.A(new_n1067), .B(new_n1069), .C1(G143), .C2(new_n745), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n1070), .B1(new_n202), .B2(new_n768), .C1(new_n337), .C2(new_n752), .ZN(new_n1071));
  XOR2_X1   g0871(.A(new_n1071), .B(KEYINPUT112), .Z(new_n1072));
  OAI22_X1  g0872(.A1(new_n755), .A2(new_n1011), .B1(new_n819), .B2(new_n761), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT52), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n752), .A2(new_n747), .B1(new_n744), .B2(new_n760), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n736), .B2(G303), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1074), .B(new_n1076), .C1(new_n759), .C2(new_n740), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G116), .B2(new_n780), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n1078), .A2(new_n314), .A3(new_n779), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n730), .B1(new_n1072), .B2(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n249), .A2(new_n723), .B1(G97), .B2(new_n664), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1081), .A2(new_n731), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n966), .A2(new_n717), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1080), .A2(new_n722), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n1062), .B2(new_n720), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1064), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(G390));
  INV_X1    g0887(.A(new_n792), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n793), .B1(new_n710), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n845), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n919), .B1(new_n897), .B2(new_n902), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n920), .A2(new_n922), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n918), .B1(new_n913), .B2(new_n845), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1091), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(G330), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n904), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n697), .A2(KEYINPUT90), .A3(G330), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n794), .B(new_n845), .C1(new_n1098), .C2(new_n698), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n831), .A2(G330), .A3(new_n794), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n1090), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(KEYINPUT113), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT113), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1100), .A2(new_n1103), .A3(new_n1090), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1099), .A2(new_n1089), .A3(new_n1102), .A4(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n794), .B1(new_n1098), .B2(new_n698), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1096), .B1(new_n1106), .B2(new_n1090), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n913), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1105), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1099), .B(new_n1091), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1110));
  AND3_X1   g0910(.A1(new_n908), .A2(new_n630), .A3(new_n926), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1097), .A2(new_n1109), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n665), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT114), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1097), .A2(new_n1110), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1112), .A2(KEYINPUT114), .A3(new_n665), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1115), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1097), .A2(new_n721), .A3(new_n1110), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n920), .A2(new_n805), .A3(new_n922), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n807), .A2(new_n363), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n758), .A2(new_n770), .ZN(new_n1124));
  INV_X1    g0924(.A(G137), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n768), .A2(new_n1125), .B1(new_n811), .B2(new_n761), .ZN(new_n1126));
  XOR2_X1   g0926(.A(KEYINPUT54), .B(G143), .Z(new_n1127));
  AOI211_X1 g0927(.A(new_n1124), .B(new_n1126), .C1(new_n823), .C2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n756), .A2(G128), .ZN(new_n1129));
  INV_X1    g0929(.A(G125), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n752), .A2(new_n409), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT53), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n265), .B1(new_n1130), .B2(new_n744), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(new_n1132), .B2(new_n1131), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n778), .A2(G50), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1128), .A2(new_n1129), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n823), .A2(G97), .B1(G283), .B2(new_n756), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n214), .B2(new_n768), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT115), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(G68), .B2(new_n778), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n776), .A2(G116), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n265), .B1(new_n745), .B2(G294), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1140), .A2(new_n775), .A3(new_n1141), .A4(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1136), .B1(new_n1143), .B2(new_n1065), .ZN(new_n1144));
  XOR2_X1   g0944(.A(new_n1144), .B(KEYINPUT116), .Z(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n730), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1122), .A2(new_n722), .A3(new_n1123), .A4(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1120), .A2(new_n1121), .A3(new_n1147), .ZN(G378));
  XNOR2_X1  g0948(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n412), .A2(new_n638), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n427), .B2(new_n431), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n427), .A2(new_n431), .A3(new_n1151), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1149), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1154), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1149), .ZN(new_n1157));
  NOR3_X1   g0957(.A1(new_n1156), .A2(new_n1152), .A3(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1155), .A2(new_n1158), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1095), .B(new_n1159), .C1(new_n896), .C2(new_n905), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1159), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n906), .B2(G330), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n1160), .A2(new_n1162), .B1(new_n923), .B2(new_n916), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT118), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT119), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1166), .B1(new_n1167), .B2(new_n924), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n907), .A2(new_n1159), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n906), .A2(new_n1161), .A3(G330), .ZN(new_n1170));
  AND4_X1   g0970(.A1(new_n1166), .A2(new_n1169), .A3(new_n924), .A4(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1165), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1169), .A2(new_n924), .A3(new_n1170), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(KEYINPUT119), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1169), .A2(new_n1166), .A3(new_n924), .A4(new_n1170), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1174), .A2(new_n1164), .A3(new_n1163), .A4(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1172), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1112), .A2(new_n1111), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT120), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1112), .A2(KEYINPUT120), .A3(new_n1111), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT57), .B1(new_n1177), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT57), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n1163), .B2(new_n1173), .ZN(new_n1185));
  AND3_X1   g0985(.A1(new_n1112), .A2(KEYINPUT120), .A3(new_n1111), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT120), .B1(new_n1112), .B2(new_n1111), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1185), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n665), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1183), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1159), .A2(new_n805), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n749), .A2(new_n352), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n756), .A2(G116), .B1(G283), .B2(new_n745), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1193), .B1(new_n214), .B2(new_n761), .C1(new_n322), .C2(new_n740), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1192), .B(new_n1194), .C1(G97), .C2(new_n736), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n374), .A2(G41), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1195), .A2(new_n997), .A3(new_n1040), .A4(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(KEYINPUT117), .B(KEYINPUT58), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1197), .B(new_n1198), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n755), .A2(new_n1130), .B1(new_n1125), .B2(new_n740), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n774), .A2(new_n1127), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n776), .A2(G128), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(new_n409), .C2(new_n758), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1200), .B(new_n1203), .C1(G132), .C2(new_n736), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT59), .ZN(new_n1205));
  AOI21_X1  g1005(.A(G33), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(G41), .B1(new_n745), .B2(G124), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n770), .C2(new_n749), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1209));
  AOI21_X1  g1009(.A(G41), .B1(new_n371), .B2(KEYINPUT3), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n1208), .A2(new_n1209), .B1(G50), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n730), .B1(new_n1199), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n806), .A2(new_n202), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1191), .A2(new_n722), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(new_n1177), .B2(new_n721), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1190), .A2(new_n1216), .ZN(G375));
  NAND2_X1  g1017(.A1(new_n1090), .A2(new_n805), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G77), .A2(new_n778), .B1(new_n745), .B2(G303), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n776), .A2(G283), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1219), .A2(new_n314), .A3(new_n1039), .A4(new_n1220), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n823), .A2(G107), .B1(G294), .B2(new_n756), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n246), .B2(new_n768), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1221), .B(new_n1223), .C1(G97), .C2(new_n774), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n736), .A2(new_n1127), .B1(G128), .B2(new_n745), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n811), .B2(new_n755), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1010), .B1(G150), .B2(new_n741), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1192), .B1(G50), .B2(new_n780), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1227), .B(new_n1228), .C1(new_n770), .C2(new_n752), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1226), .B(new_n1229), .C1(G137), .C2(new_n776), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n730), .B1(new_n1224), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n807), .A2(new_n293), .ZN(new_n1232));
  AND4_X1   g1032(.A1(new_n722), .A2(new_n1218), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n1109), .B2(new_n721), .ZN(new_n1234));
  OR2_X1    g1034(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n971), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1117), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1234), .B1(new_n1236), .B2(new_n1237), .ZN(G381));
  NAND2_X1  g1038(.A1(G375), .A2(KEYINPUT122), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT122), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1190), .A2(new_n1240), .A3(new_n1216), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(G378), .ZN(new_n1243));
  INV_X1    g1043(.A(G381), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1245), .B(KEYINPUT121), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1246), .A2(new_n1026), .A3(new_n1086), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .A4(new_n1248), .ZN(G407));
  NAND3_X1  g1049(.A1(new_n1242), .A2(new_n632), .A3(new_n1243), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(G407), .A2(G213), .A3(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT123), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(G407), .A2(new_n1250), .A3(KEYINPUT123), .A4(G213), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(G409));
  INV_X1    g1055(.A(KEYINPUT126), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT60), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1235), .A2(new_n1257), .ZN(new_n1258));
  OR3_X1    g1058(.A1(new_n1109), .A2(new_n1111), .A3(new_n1257), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1258), .A2(new_n665), .A3(new_n1117), .A4(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1234), .ZN(new_n1261));
  INV_X1    g1061(.A(G384), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1260), .A2(G384), .A3(new_n1234), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(G213), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1266), .A2(G343), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(G2897), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1265), .A2(new_n1270), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1263), .B(new_n1264), .C1(new_n1269), .C2(new_n1268), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1177), .A2(new_n971), .A3(new_n1182), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1163), .A2(new_n1173), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n721), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1274), .A2(new_n1214), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1243), .ZN(new_n1278));
  OAI211_X1 g1078(.A(G378), .B(new_n1216), .C1(new_n1183), .C2(new_n1189), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1273), .B1(new_n1280), .B2(new_n1268), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n1265), .B(new_n1267), .C1(new_n1278), .C2(new_n1279), .ZN(new_n1282));
  OAI21_X1  g1082(.A(KEYINPUT63), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1267), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1265), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT63), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT61), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(G393), .B(G396), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1023), .A2(new_n1025), .A3(new_n1086), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1086), .B1(new_n993), .B2(new_n1021), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1291), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1022), .A2(G390), .ZN(new_n1296));
  NOR3_X1   g1096(.A1(new_n1296), .A2(new_n1293), .A3(new_n1290), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1289), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1298), .B(KEYINPUT124), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1283), .A2(new_n1288), .A3(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(KEYINPUT125), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT62), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1280), .A2(new_n1268), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1273), .ZN(new_n1305));
  AOI22_X1  g1105(.A1(new_n1282), .A2(new_n1303), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT61), .B1(new_n1286), .B2(KEYINPUT62), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1302), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1256), .B1(new_n1300), .B2(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1283), .A2(new_n1299), .A3(new_n1288), .ZN(new_n1310));
  OAI22_X1  g1110(.A1(new_n1286), .A2(KEYINPUT62), .B1(new_n1284), .B2(new_n1273), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1289), .B1(new_n1282), .B2(new_n1303), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  OAI211_X1 g1113(.A(KEYINPUT126), .B(new_n1310), .C1(new_n1313), .C2(new_n1302), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1309), .A2(new_n1314), .ZN(G405));
  AOI21_X1  g1115(.A(G378), .B1(new_n1190), .B2(new_n1216), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1279), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1285), .A2(KEYINPUT127), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(new_n1318), .B(new_n1319), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(new_n1320), .B(new_n1301), .ZN(G402));
endmodule


