//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT73), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G116), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT67), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  XOR2_X1   g009(.A(KEYINPUT2), .B(G113), .Z(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT2), .B(G113), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n193), .A2(new_n198), .A3(new_n194), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(G143), .B(G146), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT0), .B(G128), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT68), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT68), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n206), .B(new_n211), .C1(new_n207), .C2(new_n208), .ZN(new_n212));
  INV_X1    g026(.A(G137), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n213), .A2(G134), .B1(KEYINPUT64), .B2(KEYINPUT11), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n213), .A2(G134), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT65), .B(G131), .ZN(new_n217));
  INV_X1    g031(.A(G134), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(G137), .ZN(new_n219));
  NAND2_X1  g033(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n219), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  AND3_X1   g037(.A1(new_n216), .A2(new_n217), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G131), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n225), .B1(new_n216), .B2(new_n223), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n210), .B(new_n212), .C1(new_n224), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT1), .B1(new_n203), .B2(G146), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n203), .A2(G146), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n201), .A2(G143), .ZN(new_n230));
  OAI211_X1 g044(.A(G128), .B(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G128), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n202), .B(new_n204), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n216), .A2(new_n217), .A3(new_n223), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n213), .A2(G134), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n218), .A2(G137), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n237), .A3(KEYINPUT66), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n238), .B(G131), .C1(KEYINPUT66), .C2(new_n236), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n234), .A2(new_n235), .A3(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n227), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT72), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n200), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n227), .A2(KEYINPUT72), .A3(new_n240), .ZN(new_n244));
  AOI211_X1 g058(.A(new_n188), .B(KEYINPUT28), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n241), .A2(new_n242), .ZN(new_n246));
  INV_X1    g060(.A(new_n200), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(new_n244), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT28), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT73), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n241), .B(new_n200), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT28), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  OR2_X1    g068(.A1(KEYINPUT69), .A2(G953), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT69), .A2(G953), .ZN(new_n256));
  AND2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G237), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(G210), .A3(new_n258), .ZN(new_n259));
  XOR2_X1   g073(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n260));
  XNOR2_X1  g074(.A(new_n259), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT26), .B(G101), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n263), .A2(KEYINPUT29), .ZN(new_n264));
  AOI21_X1  g078(.A(G902), .B1(new_n254), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT30), .ZN(new_n266));
  AND4_X1   g080(.A1(new_n235), .A2(new_n239), .A3(new_n233), .A4(new_n231), .ZN(new_n267));
  INV_X1    g081(.A(new_n222), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n236), .B1(new_n268), .B2(new_n220), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n237), .B1(new_n219), .B2(new_n221), .ZN(new_n270));
  OAI21_X1  g084(.A(G131), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n209), .B1(new_n271), .B2(new_n235), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n266), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n273), .B(new_n200), .C1(new_n241), .C2(new_n266), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n241), .A2(new_n200), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n263), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT29), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n227), .A2(KEYINPUT72), .A3(new_n240), .ZN(new_n280));
  AOI21_X1  g094(.A(KEYINPUT72), .B1(new_n227), .B2(new_n240), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n280), .A2(new_n281), .A3(new_n200), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n188), .B1(new_n282), .B2(KEYINPUT28), .ZN(new_n283));
  INV_X1    g097(.A(new_n272), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n247), .B1(new_n284), .B2(new_n240), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT28), .B1(new_n275), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n248), .A2(KEYINPUT73), .A3(new_n249), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n283), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n263), .B(KEYINPUT71), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n279), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n187), .B1(new_n265), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT32), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n289), .B1(new_n251), .B2(new_n286), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n274), .A2(new_n276), .A3(new_n263), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT31), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n274), .A2(new_n276), .A3(KEYINPUT31), .A4(new_n263), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT74), .B1(new_n295), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n288), .A2(new_n290), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT74), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(new_n300), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT75), .B1(G472), .B2(G902), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NOR3_X1   g122(.A1(KEYINPUT75), .A2(G472), .A3(G902), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n294), .B1(new_n306), .B2(new_n311), .ZN(new_n312));
  AOI221_X4 g126(.A(KEYINPUT74), .B1(new_n298), .B2(new_n299), .C1(new_n288), .C2(new_n290), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n304), .B1(new_n303), .B2(new_n300), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n294), .B(new_n311), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n293), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(KEYINPUT9), .B(G234), .ZN(new_n318));
  OAI21_X1  g132(.A(G221), .B1(new_n318), .B2(G902), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G469), .ZN(new_n321));
  INV_X1    g135(.A(G902), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n271), .A2(new_n235), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT10), .ZN(new_n324));
  INV_X1    g138(.A(G104), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT3), .B1(new_n325), .B2(G107), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n327));
  INV_X1    g141(.A(G107), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n328), .A3(G104), .ZN(new_n329));
  INV_X1    g143(.A(G101), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n325), .A2(G107), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n326), .A2(new_n329), .A3(new_n330), .A4(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n325), .A2(G107), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n328), .A2(G104), .ZN(new_n334));
  OAI21_X1  g148(.A(G101), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n231), .A2(new_n332), .A3(new_n335), .A4(new_n233), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n324), .B1(new_n336), .B2(KEYINPUT84), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(KEYINPUT84), .A3(new_n324), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n326), .A2(new_n329), .A3(new_n331), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT4), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(new_n342), .A3(G101), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n210), .A2(new_n212), .A3(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT83), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n341), .A2(G101), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n332), .A2(KEYINPUT4), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n341), .A2(G101), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n349), .A2(KEYINPUT83), .A3(KEYINPUT4), .A4(new_n332), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n344), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n323), .B1(new_n340), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(new_n350), .ZN(new_n353));
  INV_X1    g167(.A(new_n344), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AND3_X1   g169(.A1(new_n336), .A2(KEYINPUT84), .A3(new_n324), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(new_n337), .ZN(new_n357));
  INV_X1    g171(.A(new_n323), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n355), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n352), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n257), .A2(G227), .ZN(new_n361));
  XOR2_X1   g175(.A(G110), .B(G140), .Z(new_n362));
  XNOR2_X1  g176(.A(new_n361), .B(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n360), .A2(KEYINPUT88), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n336), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n233), .A2(new_n231), .B1(new_n332), .B2(new_n335), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n323), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT12), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n323), .B(KEYINPUT12), .C1(new_n365), .C2(new_n366), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n363), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n359), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n364), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(KEYINPUT88), .B1(new_n360), .B2(new_n363), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n321), .B(new_n322), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT86), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n359), .A2(new_n371), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT85), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n359), .A2(new_n371), .A3(KEYINPUT85), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n372), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n352), .A2(new_n372), .A3(new_n359), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n378), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n359), .A2(KEYINPUT85), .A3(new_n371), .ZN(new_n387));
  AOI21_X1  g201(.A(KEYINPUT85), .B1(new_n359), .B2(new_n371), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n363), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(KEYINPUT86), .A3(new_n384), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n321), .B1(new_n391), .B2(new_n322), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n377), .B1(new_n392), .B2(KEYINPUT87), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT87), .ZN(new_n394));
  AOI21_X1  g208(.A(G902), .B1(new_n386), .B2(new_n390), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n394), .B1(new_n395), .B2(new_n321), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n320), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G217), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n398), .B1(G234), .B2(new_n322), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n257), .A2(G221), .A3(G234), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n401), .B(KEYINPUT79), .ZN(new_n402));
  XNOR2_X1  g216(.A(KEYINPUT22), .B(G137), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n402), .B(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT23), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n406), .B1(new_n189), .B2(G128), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n189), .A2(G128), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n232), .A2(KEYINPUT23), .A3(G119), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G110), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT76), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n413), .B1(new_n232), .B2(G119), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n189), .A2(KEYINPUT76), .A3(G128), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n414), .B(new_n415), .C1(new_n189), .C2(G128), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT24), .B(G110), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT78), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n419), .B(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(G125), .B(G140), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT16), .ZN(new_n423));
  INV_X1    g237(.A(G140), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G125), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n423), .B(G146), .C1(KEYINPUT16), .C2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n422), .A2(new_n201), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n421), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n416), .A2(new_n417), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(KEYINPUT77), .ZN(new_n430));
  OR2_X1    g244(.A1(new_n410), .A2(new_n411), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n423), .B1(KEYINPUT16), .B2(new_n425), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n201), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n426), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n430), .A2(new_n431), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n428), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT80), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT80), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n428), .A2(new_n438), .A3(new_n435), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n405), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n405), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT81), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n444), .A2(KEYINPUT25), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n443), .A2(new_n322), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(new_n439), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n438), .B1(new_n428), .B2(new_n435), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n404), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(new_n322), .A3(new_n441), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n445), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n400), .B1(new_n447), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n399), .A2(G902), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(KEYINPUT82), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n443), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G110), .B(G122), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n346), .A2(new_n342), .B1(new_n197), .B2(new_n199), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n332), .A2(KEYINPUT4), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT83), .B1(new_n461), .B2(new_n349), .ZN(new_n462));
  AND4_X1   g276(.A1(KEYINPUT83), .A2(new_n349), .A3(KEYINPUT4), .A4(new_n332), .ZN(new_n463));
  OAI211_X1 g277(.A(KEYINPUT89), .B(new_n460), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n190), .A2(new_n192), .A3(KEYINPUT5), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n465), .B(G113), .C1(KEYINPUT5), .C2(new_n190), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n466), .B1(new_n198), .B2(new_n193), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n332), .A2(new_n335), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n464), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n199), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n198), .B1(new_n194), .B2(new_n193), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n343), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(new_n348), .B2(new_n350), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n475), .A2(KEYINPUT89), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n459), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n469), .B1(new_n475), .B2(KEYINPUT89), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT89), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n478), .A2(new_n481), .A3(new_n458), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n477), .A2(KEYINPUT6), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G125), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n234), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(new_n484), .B2(new_n209), .ZN(new_n486));
  INV_X1    g300(.A(G224), .ZN(new_n487));
  OR2_X1    g301(.A1(new_n487), .A2(G953), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT91), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n486), .B(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n458), .A2(KEYINPUT6), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  AOI211_X1 g306(.A(KEYINPUT90), .B(new_n492), .C1(new_n478), .C2(new_n481), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT90), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n478), .A2(new_n481), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n494), .B1(new_n495), .B2(new_n491), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n483), .B(new_n490), .C1(new_n493), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n488), .A2(KEYINPUT7), .ZN(new_n498));
  XOR2_X1   g312(.A(new_n486), .B(new_n498), .Z(new_n499));
  XOR2_X1   g313(.A(new_n458), .B(KEYINPUT8), .Z(new_n500));
  NAND2_X1  g314(.A1(new_n467), .A2(new_n468), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n500), .B1(new_n470), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(G902), .B1(new_n503), .B2(new_n482), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n497), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(G210), .B1(G237), .B2(G902), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n497), .A2(new_n506), .A3(new_n504), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(G214), .B1(G237), .B2(G902), .ZN(new_n511));
  INV_X1    g325(.A(G952), .ZN(new_n512));
  AOI211_X1 g326(.A(G953), .B(new_n512), .C1(G234), .C2(G237), .ZN(new_n513));
  AOI211_X1 g327(.A(new_n322), .B(new_n257), .C1(G234), .C2(G237), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT21), .B(G898), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(KEYINPUT97), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n513), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n510), .A2(new_n511), .A3(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n257), .A2(G143), .A3(G214), .A4(new_n258), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n255), .A2(G214), .A3(new_n258), .A4(new_n256), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n203), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT18), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n520), .B(new_n522), .C1(new_n523), .C2(new_n225), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n422), .B(new_n201), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n520), .A2(new_n522), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n523), .A2(new_n225), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT92), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT92), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n527), .A2(new_n531), .A3(new_n528), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n526), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n217), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n527), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT17), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n520), .A2(new_n217), .A3(new_n522), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n217), .B1(new_n520), .B2(new_n522), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n434), .B1(new_n539), .B2(KEYINPUT17), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n533), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(G113), .B(G122), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(new_n325), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT94), .ZN(new_n544));
  INV_X1    g358(.A(new_n532), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n531), .B1(new_n527), .B2(new_n528), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n524), .B(new_n525), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n535), .A2(new_n537), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n422), .B(KEYINPUT19), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n201), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT93), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT93), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n549), .A2(new_n552), .A3(new_n201), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(new_n426), .A3(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n547), .B1(new_n548), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n543), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n541), .A2(new_n544), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(G475), .A2(G902), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT95), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n540), .A2(new_n538), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(new_n547), .A3(new_n544), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n554), .A2(new_n548), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(new_n533), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n562), .B1(new_n564), .B2(new_n543), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT95), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n566), .A3(new_n558), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n560), .A2(new_n567), .A3(KEYINPUT20), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n566), .B1(new_n565), .B2(new_n558), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT20), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n562), .B1(new_n541), .B2(new_n543), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n322), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n569), .A2(new_n570), .B1(new_n572), .B2(G475), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n203), .A2(G128), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n232), .A2(G143), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(new_n218), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n191), .A2(KEYINPUT14), .A3(G122), .ZN(new_n579));
  XNOR2_X1  g393(.A(G116), .B(G122), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  OAI211_X1 g395(.A(G107), .B(new_n579), .C1(new_n581), .C2(KEYINPUT14), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n578), .B(new_n582), .C1(G107), .C2(new_n581), .ZN(new_n583));
  INV_X1    g397(.A(new_n575), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n584), .A2(KEYINPUT13), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n576), .B1(new_n584), .B2(KEYINPUT13), .ZN(new_n586));
  OAI21_X1  g400(.A(G134), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n577), .A2(new_n218), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n580), .B(new_n328), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n583), .A2(new_n590), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n318), .A2(new_n398), .A3(G953), .ZN(new_n592));
  XOR2_X1   g406(.A(new_n591), .B(new_n592), .Z(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n322), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT15), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n595), .A2(KEYINPUT96), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n595), .A2(KEYINPUT96), .ZN(new_n597));
  OAI21_X1  g411(.A(G478), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(new_n594), .B(new_n598), .Z(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n574), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n519), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n317), .A2(new_n397), .A3(new_n457), .A4(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  NOR3_X1   g418(.A1(new_n383), .A2(new_n378), .A3(new_n385), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT86), .B1(new_n389), .B2(new_n384), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n322), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(KEYINPUT87), .A3(G469), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n396), .A2(new_n608), .A3(new_n376), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n319), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n322), .B1(new_n313), .B2(new_n314), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(G472), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n311), .B1(new_n313), .B2(new_n314), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n457), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n610), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT100), .ZN(new_n617));
  OR2_X1    g431(.A1(new_n616), .A2(KEYINPUT100), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n593), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n591), .B(new_n592), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n620), .A2(KEYINPUT100), .A3(new_n616), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(G478), .A3(new_n322), .ZN(new_n623));
  INV_X1    g437(.A(G478), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n594), .A2(KEYINPUT101), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT101), .B1(new_n594), .B2(new_n624), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n574), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT98), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n508), .A2(new_n630), .A3(new_n509), .ZN(new_n631));
  INV_X1    g445(.A(new_n511), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n506), .B1(new_n497), .B2(new_n504), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n632), .B1(new_n633), .B2(KEYINPUT98), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n631), .A2(KEYINPUT99), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(KEYINPUT99), .B1(new_n631), .B2(new_n634), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n635), .A2(new_n636), .A3(new_n517), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n615), .A2(new_n629), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT34), .B(G104), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  NAND3_X1  g454(.A1(new_n599), .A2(new_n568), .A3(new_n573), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n615), .A2(new_n637), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT35), .B(G107), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  AND2_X1   g459(.A1(new_n612), .A2(new_n613), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n405), .A2(KEYINPUT36), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(new_n436), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n648), .A2(new_n455), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n453), .A2(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n397), .A2(new_n646), .A3(new_n602), .A4(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT37), .B(G110), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  NAND2_X1  g468(.A1(new_n613), .A2(KEYINPUT32), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n315), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n650), .B1(new_n656), .B2(new_n293), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n635), .A2(new_n636), .ZN(new_n658));
  INV_X1    g472(.A(G900), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n513), .B1(new_n514), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n641), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n657), .A2(new_n397), .A3(new_n658), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  NAND2_X1  g477(.A1(new_n290), .A2(new_n252), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n664), .B(KEYINPUT103), .Z(new_n665));
  INV_X1    g479(.A(new_n296), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n322), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G472), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n656), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n510), .B(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n574), .A2(new_n600), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n650), .A3(new_n511), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n670), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n660), .B(KEYINPUT39), .Z(new_n676));
  NAND2_X1  g490(.A1(new_n397), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(KEYINPUT40), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT104), .B(G143), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G45));
  NAND2_X1  g496(.A1(new_n568), .A2(new_n573), .ZN(new_n683));
  INV_X1    g497(.A(new_n660), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n627), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n657), .A2(new_n397), .A3(new_n658), .A4(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  INV_X1    g502(.A(new_n457), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n656), .B2(new_n293), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n374), .A2(new_n375), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n322), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(G469), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n319), .A3(new_n376), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n690), .A2(new_n637), .A3(new_n629), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT41), .B(G113), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G15));
  NAND4_X1  g512(.A1(new_n690), .A2(new_n637), .A3(new_n642), .A4(new_n695), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G116), .ZN(G18));
  NOR3_X1   g514(.A1(new_n635), .A2(new_n636), .A3(new_n694), .ZN(new_n701));
  INV_X1    g515(.A(new_n601), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n657), .A2(new_n701), .A3(new_n702), .A4(new_n518), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  OAI21_X1  g518(.A(new_n300), .B1(new_n254), .B2(new_n289), .ZN(new_n705));
  XOR2_X1   g519(.A(new_n310), .B(KEYINPUT105), .Z(new_n706));
  AOI22_X1  g520(.A1(new_n612), .A2(KEYINPUT106), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n611), .A2(new_n708), .A3(G472), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n694), .A2(new_n517), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n707), .A2(new_n457), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n658), .A2(new_n673), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT107), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(G902), .B1(new_n302), .B2(new_n305), .ZN(new_n714));
  OAI21_X1  g528(.A(KEYINPUT106), .B1(new_n714), .B2(new_n187), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n705), .A2(new_n706), .ZN(new_n716));
  AND4_X1   g530(.A1(new_n457), .A2(new_n715), .A3(new_n709), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n683), .A2(new_n599), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n635), .A2(new_n636), .A3(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n717), .A2(new_n719), .A3(new_n720), .A4(new_n710), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n713), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT108), .B(G122), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G24));
  AND3_X1   g538(.A1(new_n715), .A2(new_n709), .A3(new_n716), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n725), .A2(new_n701), .A3(new_n651), .A4(new_n686), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G125), .ZN(G27));
  NAND3_X1  g541(.A1(new_n389), .A2(G469), .A3(new_n384), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n321), .A2(new_n322), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n319), .B1(new_n377), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT109), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n728), .A2(new_n730), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n320), .B1(new_n735), .B2(new_n376), .ZN(new_n736));
  INV_X1    g550(.A(new_n509), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n633), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT109), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n736), .A2(new_n738), .A3(new_n739), .A4(new_n511), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n734), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n685), .A2(KEYINPUT42), .ZN(new_n742));
  AND4_X1   g556(.A1(new_n457), .A2(new_n317), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n744), .B1(new_n312), .B2(new_n316), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n655), .A2(KEYINPUT110), .A3(new_n315), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n293), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n685), .B1(new_n734), .B2(new_n740), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n457), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n743), .B1(new_n749), .B2(KEYINPUT42), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G131), .ZN(G33));
  NAND3_X1  g565(.A1(new_n690), .A2(new_n661), .A3(new_n741), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G134), .ZN(G36));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n574), .A2(new_n627), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT43), .ZN(new_n756));
  OR2_X1    g570(.A1(new_n756), .A2(new_n650), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n754), .B1(new_n757), .B2(new_n646), .ZN(new_n758));
  OR4_X1    g572(.A1(new_n754), .A2(new_n756), .A3(new_n646), .A4(new_n650), .ZN(new_n759));
  INV_X1    g573(.A(new_n733), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT45), .B1(new_n386), .B2(new_n390), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n389), .A2(KEYINPUT45), .A3(new_n384), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(G469), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n730), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT46), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n377), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n765), .A2(KEYINPUT46), .A3(new_n730), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n320), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n770), .A2(new_n676), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n758), .A2(new_n759), .A3(new_n760), .A4(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G137), .ZN(G39));
  AOI21_X1  g587(.A(new_n292), .B1(new_n655), .B2(new_n315), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(new_n689), .A3(new_n686), .A4(new_n760), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT111), .ZN(new_n776));
  AOI22_X1  g590(.A1(new_n770), .A2(new_n776), .B1(KEYINPUT112), .B2(KEYINPUT47), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n768), .A2(new_n769), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT111), .B1(new_n778), .B2(new_n320), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT47), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n777), .B(new_n779), .C1(KEYINPUT112), .C2(KEYINPUT47), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n775), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(new_n424), .ZN(G42));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n725), .A2(new_n651), .A3(new_n686), .A4(new_n741), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n733), .A2(new_n660), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n609), .A2(new_n319), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n657), .A2(new_n791), .A3(new_n702), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n789), .A2(new_n792), .A3(new_n752), .ZN(new_n793));
  INV_X1    g607(.A(new_n614), .ZN(new_n794));
  AOI22_X1  g608(.A1(new_n641), .A2(KEYINPUT114), .B1(new_n683), .B2(new_n627), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n574), .A2(new_n796), .A3(new_n599), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n519), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n794), .A2(new_n397), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n603), .A2(new_n799), .A3(new_n652), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n793), .A2(new_n800), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n696), .A2(new_n699), .A3(new_n703), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n722), .A3(new_n750), .A4(new_n802), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n651), .A2(new_n660), .A3(new_n732), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n719), .A3(new_n669), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n662), .A2(new_n726), .A3(new_n687), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT52), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n610), .A2(new_n636), .A3(new_n635), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n808), .B(new_n657), .C1(new_n661), .C2(new_n686), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n809), .A2(new_n810), .A3(new_n726), .A4(new_n805), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n788), .B1(new_n803), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n802), .A2(new_n750), .A3(new_n722), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n603), .A2(new_n799), .A3(new_n652), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n317), .A2(new_n457), .A3(new_n741), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n774), .A2(new_n601), .A3(new_n650), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n816), .A2(new_n661), .B1(new_n817), .B2(new_n791), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n815), .A2(new_n818), .A3(KEYINPUT53), .A4(new_n789), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n807), .A2(new_n811), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT117), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT117), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n812), .A2(new_n814), .A3(new_n819), .A4(new_n823), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n787), .B(new_n813), .C1(new_n822), .C2(new_n824), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n793), .A2(new_n788), .A3(new_n800), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n826), .A2(new_n722), .A3(new_n750), .A4(new_n802), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n812), .ZN(new_n828));
  OR2_X1    g642(.A1(new_n828), .A2(KEYINPUT116), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(KEYINPUT116), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n812), .B1(new_n803), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n832), .B1(new_n831), .B2(new_n803), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n829), .A2(new_n830), .B1(new_n833), .B2(new_n788), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n825), .B1(new_n834), .B2(new_n787), .ZN(new_n835));
  INV_X1    g649(.A(new_n513), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n756), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n694), .A2(new_n733), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n457), .A3(new_n747), .A4(new_n838), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT48), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n837), .A2(new_n701), .A3(new_n717), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(KEYINPUT118), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n689), .A2(new_n836), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n670), .A2(new_n838), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  AOI211_X1 g659(.A(new_n512), .B(G953), .C1(new_n845), .C2(new_n629), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n840), .A2(new_n842), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n837), .A2(new_n717), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n733), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n783), .A2(new_n784), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n693), .A2(new_n376), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(new_n319), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n849), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n672), .A2(new_n632), .A3(new_n695), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n848), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT50), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n837), .A2(new_n651), .A3(new_n725), .A4(new_n838), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n845), .A2(new_n574), .A3(new_n628), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n853), .A2(new_n856), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT51), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n847), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n861), .B1(new_n860), .B2(new_n859), .ZN(new_n862));
  OAI22_X1  g676(.A1(new_n835), .A2(new_n862), .B1(G952), .B2(G953), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n457), .A2(new_n319), .A3(new_n511), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n851), .A2(KEYINPUT49), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n851), .A2(KEYINPUT49), .ZN(new_n866));
  NOR4_X1   g680(.A1(new_n864), .A2(new_n865), .A3(new_n866), .A4(new_n755), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n867), .A2(new_n672), .A3(new_n670), .ZN(new_n868));
  XNOR2_X1  g682(.A(new_n868), .B(KEYINPUT113), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n863), .A2(new_n869), .ZN(G75));
  NOR2_X1   g684(.A1(new_n257), .A2(G952), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n823), .B1(new_n827), .B2(new_n812), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n820), .A2(new_n821), .A3(KEYINPUT117), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n322), .B1(new_n875), .B2(new_n813), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT56), .B1(new_n876), .B2(G210), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n483), .B1(new_n496), .B2(new_n493), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(new_n490), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT55), .Z(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n872), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n803), .A2(new_n812), .ZN(new_n883));
  AOI22_X1  g697(.A1(new_n873), .A2(new_n874), .B1(new_n883), .B2(new_n788), .ZN(new_n884));
  INV_X1    g698(.A(G210), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n884), .A2(new_n885), .A3(new_n322), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n886), .A2(KEYINPUT56), .A3(new_n880), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT119), .B1(new_n882), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n880), .B1(new_n886), .B2(KEYINPUT56), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n877), .A2(new_n881), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n889), .A2(new_n890), .A3(new_n891), .A4(new_n872), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n888), .A2(new_n892), .ZN(G51));
  XNOR2_X1  g707(.A(new_n729), .B(KEYINPUT57), .ZN(new_n894));
  INV_X1    g708(.A(new_n825), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n787), .B1(new_n875), .B2(new_n813), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT120), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n899), .B(new_n894), .C1(new_n895), .C2(new_n896), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n898), .A2(new_n691), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n876), .A2(new_n764), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n871), .B1(new_n901), .B2(new_n902), .ZN(G54));
  INV_X1    g717(.A(KEYINPUT58), .ZN(new_n904));
  INV_X1    g718(.A(G475), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n876), .A2(new_n565), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n565), .B1(new_n876), .B2(new_n906), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n907), .A2(new_n908), .A3(new_n871), .ZN(G60));
  NAND2_X1  g723(.A1(G478), .A2(G902), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT59), .Z(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n622), .B1(new_n835), .B2(new_n912), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n622), .B(new_n912), .C1(new_n895), .C2(new_n896), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n872), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n913), .A2(new_n915), .ZN(G63));
  XNOR2_X1  g730(.A(KEYINPUT123), .B(KEYINPUT61), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n875), .A2(new_n813), .ZN(new_n919));
  XNOR2_X1  g733(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n398), .A2(new_n322), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n920), .B(new_n921), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n919), .A2(KEYINPUT122), .A3(new_n648), .A4(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n443), .ZN(new_n924));
  INV_X1    g738(.A(new_n922), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n924), .B1(new_n884), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n923), .A2(new_n926), .A3(new_n872), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n884), .A2(new_n925), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT122), .B1(new_n928), .B2(new_n648), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n918), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n919), .A2(new_n922), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n871), .B1(new_n931), .B2(new_n924), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n919), .A2(new_n648), .A3(new_n922), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT122), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n932), .A2(new_n935), .A3(new_n923), .A4(new_n917), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n930), .A2(new_n936), .ZN(G66));
  OAI21_X1  g751(.A(G953), .B1(new_n516), .B2(new_n487), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n802), .A2(new_n722), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n815), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n257), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n878), .B1(G898), .B2(new_n257), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(G69));
  AOI21_X1  g759(.A(new_n733), .B1(new_n795), .B2(new_n797), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n690), .A2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n772), .B1(new_n677), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n772), .B(KEYINPUT124), .C1(new_n677), .C2(new_n947), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n785), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n809), .A2(new_n726), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n680), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT62), .Z(new_n955));
  AOI21_X1  g769(.A(new_n942), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n273), .B1(new_n241), .B2(new_n266), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(new_n549), .Z(new_n958));
  OR2_X1    g772(.A1(new_n956), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n257), .A2(G900), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n771), .A2(new_n457), .A3(new_n719), .A4(new_n747), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n772), .A2(new_n752), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n953), .A2(new_n750), .ZN(new_n963));
  OR3_X1    g777(.A1(new_n785), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n960), .B1(new_n964), .B2(new_n257), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT125), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n958), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AOI211_X1 g781(.A(KEYINPUT125), .B(new_n960), .C1(new_n964), .C2(new_n257), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n959), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(G227), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n942), .B1(new_n970), .B2(new_n659), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT126), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n969), .A2(new_n973), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n959), .B(new_n972), .C1(new_n967), .C2(new_n968), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(G72));
  NOR2_X1   g790(.A1(new_n277), .A2(new_n263), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT63), .Z(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n964), .B2(new_n940), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n978), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(new_n982), .B2(new_n981), .ZN(new_n984));
  INV_X1    g798(.A(new_n980), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n278), .B1(new_n276), .B2(new_n274), .ZN(new_n986));
  OR4_X1    g800(.A1(new_n834), .A2(new_n977), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n952), .A2(new_n955), .A3(new_n941), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n980), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n871), .B1(new_n989), .B2(new_n986), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n984), .A2(new_n987), .A3(new_n990), .ZN(G57));
endmodule


