//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n526, new_n527, new_n528,
    new_n529, new_n530, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n540, new_n542, new_n543, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n557, new_n558, new_n559, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n595,
    new_n598, new_n600, new_n601, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1133, new_n1134, new_n1135;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT65), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT66), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(new_n455), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n452), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(G2106), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT68), .Z(G319));
  NAND2_X1  g037(.A1(KEYINPUT69), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(KEYINPUT69), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G137), .ZN(new_n468));
  NAND2_X1  g043(.A1(G101), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  XNOR2_X1  g046(.A(KEYINPUT3), .B(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n470), .A2(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n467), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT70), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n478), .A2(new_n479), .A3(G124), .ZN(new_n480));
  INV_X1    g055(.A(G124), .ZN(new_n481));
  OAI21_X1  g056(.A(KEYINPUT70), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  AND3_X1   g057(.A1(KEYINPUT69), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n483));
  AOI21_X1  g058(.A(KEYINPUT3), .B1(KEYINPUT69), .B2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n480), .A2(new_n482), .A3(new_n487), .A4(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND3_X1  g066(.A1(new_n467), .A2(KEYINPUT4), .A3(G138), .ZN(new_n492));
  NAND2_X1  g067(.A1(G102), .A2(G2104), .ZN(new_n493));
  AOI21_X1  g068(.A(G2105), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g069(.A(KEYINPUT71), .B(G114), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n467), .A2(G126), .B1(new_n495), .B2(G2104), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT4), .B1(new_n496), .B2(new_n471), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n472), .A2(G138), .A3(new_n471), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n494), .B1(new_n497), .B2(new_n498), .ZN(G164));
  AND2_X1   g074(.A1(KEYINPUT6), .A2(G651), .ZN(new_n500));
  NOR2_X1   g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G50), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n506), .B(new_n508), .C1(new_n500), .C2(new_n501), .ZN(new_n509));
  XOR2_X1   g084(.A(KEYINPUT72), .B(G88), .Z(new_n510));
  OAI21_X1  g085(.A(new_n505), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n506), .A2(new_n508), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n511), .A2(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  NAND2_X1  g092(.A1(new_n504), .A2(G51), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  INV_X1    g095(.A(new_n502), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n521), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n506), .A2(new_n508), .ZN(new_n523));
  OAI211_X1 g098(.A(new_n518), .B(new_n520), .C1(new_n522), .C2(new_n523), .ZN(G286));
  INV_X1    g099(.A(G286), .ZN(G168));
  NAND2_X1  g100(.A1(new_n504), .A2(G52), .ZN(new_n526));
  INV_X1    g101(.A(G90), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n527), .B2(new_n509), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n529), .A2(new_n514), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n528), .A2(new_n530), .ZN(G301));
  INV_X1    g106(.A(G301), .ZN(G171));
  NAND2_X1  g107(.A1(new_n504), .A2(G43), .ZN(new_n533));
  INV_X1    g108(.A(G81), .ZN(new_n534));
  OAI21_X1  g109(.A(new_n533), .B1(new_n534), .B2(new_n509), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n514), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G860), .ZN(G153));
  AND3_X1   g114(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G36), .ZN(G176));
  NAND2_X1  g116(.A1(G1), .A2(G3), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT8), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n540), .A2(new_n543), .ZN(G188));
  NAND2_X1  g119(.A1(G78), .A2(G543), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT73), .B(G65), .Z(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n546), .B2(new_n523), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G651), .ZN(new_n548));
  INV_X1    g123(.A(new_n509), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G91), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g126(.A(G53), .B(G543), .C1(new_n500), .C2(new_n501), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT9), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(G299));
  NAND2_X1  g131(.A1(new_n549), .A2(G87), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n504), .A2(G49), .ZN(new_n558));
  OAI21_X1  g133(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(G288));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n561));
  INV_X1    g136(.A(G61), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n523), .B2(new_n562), .ZN(new_n563));
  AND2_X1   g138(.A1(G73), .A2(G543), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT75), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT74), .A4(G61), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G651), .ZN(new_n568));
  OAI211_X1 g143(.A(G48), .B(G543), .C1(new_n500), .C2(new_n501), .ZN(new_n569));
  INV_X1    g144(.A(G86), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n509), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(G305));
  NAND2_X1  g148(.A1(new_n504), .A2(G47), .ZN(new_n574));
  INV_X1    g149(.A(G85), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(new_n509), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n514), .B2(new_n578), .ZN(G290));
  INV_X1    g154(.A(G868), .ZN(new_n580));
  NOR2_X1   g155(.A1(G171), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n504), .A2(G54), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n512), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n584), .B2(new_n514), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT77), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n549), .A2(G92), .ZN(new_n587));
  XOR2_X1   g162(.A(new_n587), .B(KEYINPUT10), .Z(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n582), .B1(new_n590), .B2(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(KEYINPUT76), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n592), .B1(KEYINPUT76), .B2(new_n581), .ZN(G321));
  XOR2_X1   g168(.A(G321), .B(KEYINPUT78), .Z(G284));
  NAND2_X1  g169(.A1(G286), .A2(G868), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(new_n555), .B2(G868), .ZN(G297));
  OAI21_X1  g171(.A(new_n595), .B1(new_n555), .B2(G868), .ZN(G280));
  XNOR2_X1  g172(.A(KEYINPUT79), .B(G559), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n590), .B1(G860), .B2(new_n598), .ZN(G148));
  NAND2_X1  g174(.A1(new_n590), .A2(new_n598), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(G868), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(G868), .B2(new_n538), .ZN(G323));
  XNOR2_X1  g177(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g178(.A1(new_n471), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT12), .Z(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT13), .ZN(new_n606));
  INV_X1    g181(.A(G2100), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n478), .A2(G123), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n486), .A2(G135), .ZN(new_n610));
  NOR2_X1   g185(.A1(G99), .A2(G2105), .ZN(new_n611));
  OAI21_X1  g186(.A(G2104), .B1(new_n471), .B2(G111), .ZN(new_n612));
  OAI211_X1 g187(.A(new_n609), .B(new_n610), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G2096), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n608), .A2(new_n615), .ZN(G156));
  XNOR2_X1  g191(.A(G2443), .B(G2446), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2451), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2454), .ZN(new_n621));
  XOR2_X1   g196(.A(KEYINPUT15), .B(G2435), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(G2438), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2427), .B(G2430), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT82), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n623), .B(new_n625), .ZN(new_n626));
  AND2_X1   g201(.A1(new_n626), .A2(KEYINPUT14), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n621), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G1341), .B(G1348), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(G14), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT83), .Z(G401));
  XOR2_X1   g209(.A(G2084), .B(G2090), .Z(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G2067), .B(G2678), .Z(new_n637));
  NOR2_X1   g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2072), .B(G2078), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT18), .Z(new_n642));
  AOI21_X1  g217(.A(new_n638), .B1(KEYINPUT17), .B2(new_n640), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n636), .A2(new_n637), .ZN(new_n644));
  OAI211_X1 g219(.A(new_n643), .B(new_n644), .C1(KEYINPUT17), .C2(new_n640), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n639), .B(KEYINPUT84), .Z(new_n646));
  OAI211_X1 g221(.A(new_n642), .B(new_n645), .C1(new_n644), .C2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(new_n614), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(new_n607), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G227));
  XOR2_X1   g225(.A(G1956), .B(G2474), .Z(new_n651));
  XOR2_X1   g226(.A(G1961), .B(G1966), .Z(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1971), .B(G1976), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT19), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n651), .A2(new_n652), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT20), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n654), .A2(new_n656), .A3(new_n658), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n661), .B(new_n662), .C1(new_n660), .C2(new_n659), .ZN(new_n663));
  XOR2_X1   g238(.A(G1991), .B(G1996), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT86), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n663), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT85), .B(G1986), .ZN(new_n669));
  INV_X1    g244(.A(G1981), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n668), .B(new_n671), .Z(G229));
  INV_X1    g247(.A(G29), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n673), .A2(G32), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n478), .A2(G129), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n471), .A2(G105), .A3(G2104), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n486), .A2(G141), .ZN(new_n677));
  NAND3_X1  g252(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n678), .B(KEYINPUT26), .Z(new_n679));
  NAND4_X1  g254(.A1(new_n675), .A2(new_n676), .A3(new_n677), .A4(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n674), .B1(new_n680), .B2(G29), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT27), .ZN(new_n682));
  NOR2_X1   g257(.A1(G16), .A2(G21), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(G168), .B2(G16), .ZN(new_n684));
  AOI22_X1  g259(.A1(new_n682), .A2(G1996), .B1(G1966), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n673), .A2(G33), .ZN(new_n686));
  AOI22_X1  g261(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n687), .A2(new_n471), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT92), .B(KEYINPUT25), .Z(new_n689));
  NAND3_X1  g264(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n689), .B(new_n690), .Z(new_n691));
  AOI211_X1 g266(.A(new_n688), .B(new_n691), .C1(G139), .C2(new_n486), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n686), .B1(new_n692), .B2(new_n673), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(G2072), .Z(new_n694));
  INV_X1    g269(.A(KEYINPUT31), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n695), .A2(G11), .ZN(new_n696));
  NOR2_X1   g271(.A1(G164), .A2(new_n673), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G27), .B2(new_n673), .ZN(new_n698));
  INV_X1    g273(.A(G2078), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n613), .A2(new_n673), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT93), .Z(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT30), .B(G28), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n702), .B1(new_n673), .B2(new_n703), .ZN(new_n704));
  AND4_X1   g279(.A1(new_n685), .A2(new_n694), .A3(new_n700), .A4(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(G4), .A2(G16), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n590), .B2(G16), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT91), .B(G1348), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  OR2_X1    g284(.A1(new_n682), .A2(G1996), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n698), .A2(new_n699), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n684), .A2(G1966), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT28), .ZN(new_n713));
  INV_X1    g288(.A(G26), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(G29), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n714), .A2(G29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n478), .A2(G128), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n486), .A2(G140), .ZN(new_n718));
  NOR2_X1   g293(.A1(G104), .A2(G2105), .ZN(new_n719));
  OAI21_X1  g294(.A(G2104), .B1(new_n471), .B2(G116), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n717), .B(new_n718), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n716), .B1(new_n721), .B2(G29), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n715), .B1(new_n722), .B2(new_n713), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G2067), .ZN(new_n724));
  NAND4_X1  g299(.A1(new_n710), .A2(new_n711), .A3(new_n712), .A4(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n709), .A2(new_n725), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n705), .B(new_n726), .C1(G2067), .C2(new_n723), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n673), .A2(G35), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G162), .B2(new_n673), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT95), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT29), .ZN(new_n731));
  INV_X1    g306(.A(G2090), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G16), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(G5), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G171), .B2(new_n734), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT94), .B(G1961), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  AND2_X1   g313(.A1(KEYINPUT24), .A2(G34), .ZN(new_n739));
  NOR2_X1   g314(.A1(KEYINPUT24), .A2(G34), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n673), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G160), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(new_n673), .ZN(new_n743));
  INV_X1    g318(.A(G2084), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NOR4_X1   g320(.A1(new_n727), .A2(new_n733), .A3(new_n738), .A4(new_n745), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n734), .A2(KEYINPUT23), .A3(G20), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT23), .ZN(new_n748));
  INV_X1    g323(.A(G20), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n748), .B1(new_n749), .B2(G16), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n747), .B(new_n750), .C1(new_n555), .C2(new_n734), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT96), .B(G1956), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(G16), .A2(G22), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G166), .B2(G16), .ZN(new_n755));
  INV_X1    g330(.A(G1971), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n734), .A2(G23), .ZN(new_n758));
  INV_X1    g333(.A(G288), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(new_n734), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT89), .B(KEYINPUT33), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1976), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n760), .B(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n734), .A2(G6), .ZN(new_n764));
  INV_X1    g339(.A(G305), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(new_n734), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT32), .B(G1981), .Z(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n757), .A2(new_n763), .A3(new_n768), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(KEYINPUT34), .ZN(new_n770));
  NOR2_X1   g345(.A1(G16), .A2(G24), .ZN(new_n771));
  XOR2_X1   g346(.A(G290), .B(KEYINPUT88), .Z(new_n772));
  AOI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(G16), .ZN(new_n773));
  INV_X1    g348(.A(G1986), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n769), .A2(KEYINPUT34), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n673), .A2(G25), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n486), .A2(G131), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT87), .ZN(new_n779));
  INV_X1    g354(.A(G119), .ZN(new_n780));
  NOR2_X1   g355(.A1(G95), .A2(G2105), .ZN(new_n781));
  OAI21_X1  g356(.A(G2104), .B1(new_n471), .B2(G107), .ZN(new_n782));
  OAI22_X1  g357(.A1(new_n477), .A2(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n777), .B1(new_n784), .B2(new_n673), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT35), .B(G1991), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n770), .A2(new_n775), .A3(new_n776), .A4(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT36), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n789), .A2(KEYINPUT90), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n789), .A2(KEYINPUT90), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n788), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n788), .A2(new_n790), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n746), .A2(new_n753), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n734), .A2(G19), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n538), .B2(new_n734), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1341), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n695), .A2(G11), .ZN(new_n798));
  NOR3_X1   g373(.A1(new_n794), .A2(new_n797), .A3(new_n798), .ZN(G311));
  INV_X1    g374(.A(G311), .ZN(G150));
  NAND2_X1  g375(.A1(new_n549), .A2(G93), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n504), .A2(G55), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n801), .B(new_n802), .C1(new_n803), .C2(new_n514), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT97), .ZN(new_n805));
  INV_X1    g380(.A(new_n538), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT38), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n590), .A2(G559), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n812), .A2(KEYINPUT39), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT98), .Z(new_n814));
  AOI21_X1  g389(.A(G860), .B1(new_n812), .B2(KEYINPUT39), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n804), .A2(G860), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT37), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n818), .ZN(G145));
  INV_X1    g394(.A(new_n605), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n478), .A2(G130), .B1(new_n486), .B2(G142), .ZN(new_n821));
  OAI21_X1  g396(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT100), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n824), .B(new_n825), .C1(G118), .C2(new_n471), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n784), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT101), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n828), .A2(KEYINPUT101), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n820), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(new_n831), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n833), .A2(new_n605), .A3(new_n829), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(G126), .B1(new_n483), .B2(new_n484), .ZN(new_n836));
  INV_X1    g411(.A(G114), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(KEYINPUT71), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT71), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G114), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n838), .A2(new_n840), .A3(G2104), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n471), .B1(new_n836), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT4), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n498), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n492), .A2(new_n493), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(new_n471), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n721), .B(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n680), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n692), .A2(KEYINPUT99), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n835), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT102), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n835), .A2(new_n851), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n742), .B(new_n613), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n490), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n835), .A2(new_n851), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n858), .B1(new_n859), .B2(KEYINPUT102), .ZN(new_n860));
  AOI21_X1  g435(.A(G37), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n852), .A2(new_n854), .A3(new_n858), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g439(.A1(new_n804), .A2(new_n580), .ZN(new_n865));
  XOR2_X1   g440(.A(new_n809), .B(new_n600), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n589), .B(new_n555), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n867), .B(KEYINPUT41), .Z(new_n870));
  OAI21_X1  g445(.A(new_n869), .B1(new_n870), .B2(new_n866), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n765), .B(G303), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n873), .ZN(new_n875));
  INV_X1    g450(.A(G290), .ZN(new_n876));
  XNOR2_X1  g451(.A(G288), .B(KEYINPUT103), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n874), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  OR2_X1    g454(.A1(new_n875), .A2(new_n878), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT42), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n871), .B(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n865), .B1(new_n883), .B2(new_n580), .ZN(G295));
  OAI21_X1  g459(.A(new_n865), .B1(new_n883), .B2(new_n580), .ZN(G331));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n886));
  XNOR2_X1  g461(.A(G301), .B(G168), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n809), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n809), .A2(new_n887), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n809), .A2(new_n887), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(KEYINPUT106), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(new_n867), .A3(new_n892), .ZN(new_n893));
  OR2_X1    g468(.A1(new_n888), .A2(new_n889), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(new_n870), .ZN(new_n895));
  INV_X1    g470(.A(new_n881), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(G37), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n890), .A2(new_n892), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n900), .A2(new_n870), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n894), .A2(new_n868), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n881), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT43), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n899), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n897), .A2(new_n898), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n896), .B1(new_n893), .B2(new_n895), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT43), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  XOR2_X1   g484(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n904), .B1(new_n899), .B2(new_n903), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n906), .A2(new_n907), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT44), .B1(new_n913), .B2(KEYINPUT43), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n911), .B1(new_n912), .B2(new_n914), .ZN(G397));
  OAI21_X1  g490(.A(KEYINPUT107), .B1(G164), .B2(G1384), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT45), .ZN(new_n917));
  AOI21_X1  g492(.A(G1384), .B1(new_n844), .B2(new_n846), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n916), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  XOR2_X1   g496(.A(KEYINPUT108), .B(G40), .Z(new_n922));
  NOR3_X1   g497(.A1(new_n470), .A2(new_n475), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n784), .B(new_n786), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n926), .A2(KEYINPUT110), .ZN(new_n927));
  XOR2_X1   g502(.A(new_n721), .B(G2067), .Z(new_n928));
  NAND2_X1  g503(.A1(new_n680), .A2(G1996), .ZN(new_n929));
  OR2_X1    g504(.A1(new_n680), .A2(G1996), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n927), .A2(new_n931), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n926), .A2(KEYINPUT110), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n925), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n925), .A2(new_n774), .A3(new_n876), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT48), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT46), .ZN(new_n938));
  INV_X1    g513(.A(new_n925), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n938), .B1(new_n939), .B2(G1996), .ZN(new_n940));
  INV_X1    g515(.A(new_n928), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n925), .B1(new_n941), .B2(new_n680), .ZN(new_n942));
  INV_X1    g517(.A(G1996), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n925), .A2(KEYINPUT46), .A3(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n940), .A2(new_n942), .A3(new_n944), .ZN(new_n945));
  XOR2_X1   g520(.A(new_n945), .B(KEYINPUT47), .Z(new_n946));
  NAND2_X1  g521(.A1(new_n784), .A2(new_n786), .ZN(new_n947));
  OAI22_X1  g522(.A1(new_n931), .A2(new_n947), .B1(G2067), .B2(new_n721), .ZN(new_n948));
  AOI211_X1 g523(.A(new_n937), .B(new_n946), .C1(new_n925), .C2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(G303), .A2(G8), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT55), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n918), .A2(KEYINPUT45), .ZN(new_n953));
  AOI211_X1 g528(.A(new_n917), .B(G1384), .C1(new_n844), .C2(new_n846), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(G1971), .B1(new_n955), .B2(new_n923), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n918), .A2(KEYINPUT50), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT50), .ZN(new_n958));
  AOI211_X1 g533(.A(new_n958), .B(G1384), .C1(new_n844), .C2(new_n846), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n732), .B(new_n923), .C1(new_n957), .C2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  OAI211_X1 g536(.A(G8), .B(new_n952), .C1(new_n956), .C2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT111), .ZN(new_n963));
  INV_X1    g538(.A(G8), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n917), .B1(G164), .B2(G1384), .ZN(new_n965));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n847), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n923), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n756), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n964), .B1(new_n969), .B2(new_n960), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(new_n971), .A3(new_n952), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n670), .B1(new_n568), .B2(new_n572), .ZN(new_n973));
  AOI211_X1 g548(.A(G1981), .B(new_n571), .C1(new_n567), .C2(G651), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT113), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT49), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n964), .B1(new_n918), .B2(new_n923), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT49), .ZN(new_n978));
  OAI211_X1 g553(.A(KEYINPUT113), .B(new_n978), .C1(new_n973), .C2(new_n974), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n981));
  INV_X1    g556(.A(G1976), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n981), .B1(G288), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n759), .A2(KEYINPUT112), .A3(G1976), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n977), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT52), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT52), .B1(G288), .B2(new_n982), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n977), .A2(new_n983), .A3(new_n984), .A4(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n980), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n963), .A2(new_n972), .A3(new_n990), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n980), .A2(new_n982), .A3(new_n759), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n977), .B1(new_n992), .B2(new_n974), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT114), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n991), .A2(new_n996), .A3(new_n993), .ZN(new_n997));
  OAI21_X1  g572(.A(G8), .B1(new_n956), .B2(new_n961), .ZN(new_n998));
  INV_X1    g573(.A(new_n952), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n989), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n958), .B1(G164), .B2(G1384), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n918), .A2(KEYINPUT50), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n924), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1966), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n744), .A2(new_n1003), .B1(new_n968), .B2(new_n1004), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n1005), .A2(new_n964), .A3(G286), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n970), .A2(new_n971), .A3(new_n952), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n971), .B1(new_n970), .B2(new_n952), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1000), .B(new_n1006), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT63), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n963), .A2(new_n972), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1012), .A2(KEYINPUT63), .A3(new_n1000), .A4(new_n1006), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n995), .A2(new_n997), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(KEYINPUT56), .B(G2072), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n965), .A2(new_n923), .A3(new_n967), .A4(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(new_n1003), .B2(G1956), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT57), .ZN(new_n1018));
  AOI22_X1  g593(.A1(new_n547), .A2(G651), .B1(G91), .B2(new_n549), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n552), .B(KEYINPUT9), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1020), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1018), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT115), .B1(new_n551), .B2(new_n554), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1026), .A2(KEYINPUT57), .A3(new_n1022), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1017), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT118), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1028), .B(new_n1016), .C1(new_n1003), .C2(G1956), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT61), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1017), .A2(KEYINPUT118), .A3(new_n1029), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n965), .A2(new_n943), .A3(new_n923), .A4(new_n967), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n918), .A2(new_n923), .ZN(new_n1038));
  XOR2_X1   g613(.A(KEYINPUT58), .B(G1341), .Z(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1037), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n538), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT59), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1032), .A2(KEYINPUT61), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1041), .A2(KEYINPUT59), .A3(new_n538), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  OAI22_X1  g622(.A1(new_n1003), .A2(G1348), .B1(G2067), .B2(new_n1038), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT60), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1048), .A2(new_n1049), .A3(new_n590), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1038), .A2(G2067), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n923), .B1(new_n957), .B2(new_n959), .ZN(new_n1053));
  INV_X1    g628(.A(G1348), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1052), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n589), .B1(new_n1055), .B2(KEYINPUT60), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1050), .B1(new_n1051), .B2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1036), .A2(new_n1047), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1059), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1025), .A2(new_n1059), .A3(new_n1027), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1017), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT117), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1048), .A2(new_n590), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT117), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1017), .B(new_n1065), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(new_n1032), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1058), .A2(new_n1068), .ZN(new_n1069));
  XNOR2_X1  g644(.A(KEYINPUT121), .B(KEYINPUT51), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1003), .A2(new_n744), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n968), .A2(new_n1004), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n964), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(G286), .A2(G8), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1074), .B(KEYINPUT119), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1075), .B(KEYINPUT122), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1070), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1075), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1078), .B(new_n1079), .C1(new_n1005), .C2(new_n964), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT120), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n1005), .B2(new_n1079), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1083), .A2(KEYINPUT120), .A3(new_n1075), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n1077), .A2(new_n1080), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1000), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n965), .A2(new_n699), .A3(new_n923), .A4(new_n967), .ZN(new_n1089));
  INV_X1    g664(.A(G1961), .ZN(new_n1090));
  AOI22_X1  g665(.A1(new_n1088), .A2(new_n1089), .B1(new_n1053), .B2(new_n1090), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1091), .A2(G301), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1089), .A2(KEYINPUT123), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1089), .A2(KEYINPUT123), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1093), .A2(KEYINPUT53), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT126), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n1098));
  INV_X1    g673(.A(new_n470), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT124), .ZN(new_n1100));
  OAI21_X1  g675(.A(G40), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n954), .A2(new_n475), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(G2078), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1102), .A2(new_n921), .A3(KEYINPUT53), .A4(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1091), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1098), .B1(new_n1105), .B2(G171), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT126), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1092), .A2(new_n1107), .A3(new_n1095), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1097), .A2(new_n1106), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1091), .A2(G301), .A3(new_n1104), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT125), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1091), .A2(KEYINPUT125), .A3(G301), .A4(new_n1104), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(G301), .B1(new_n1095), .B2(new_n1091), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1098), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1069), .A2(new_n1087), .A3(new_n1109), .A4(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT127), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1014), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1118), .B1(new_n1014), .B2(new_n1117), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1085), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n1115), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1085), .A2(new_n1121), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1123), .A2(new_n1124), .A3(new_n1086), .ZN(new_n1125));
  NOR3_X1   g700(.A1(new_n1119), .A2(new_n1120), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n925), .A2(G1986), .A3(G290), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n935), .A2(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1128), .B(KEYINPUT109), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(new_n934), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n949), .B1(new_n1126), .B2(new_n1130), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g706(.A1(new_n633), .A2(new_n649), .ZN(new_n1133));
  AOI21_X1  g707(.A(new_n1133), .B1(new_n861), .B2(new_n862), .ZN(new_n1134));
  INV_X1    g708(.A(G229), .ZN(new_n1135));
  NAND4_X1  g709(.A1(new_n909), .A2(new_n1134), .A3(new_n461), .A4(new_n1135), .ZN(G225));
  INV_X1    g710(.A(G225), .ZN(G308));
endmodule


