//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1232, new_n1233, new_n1234, new_n1236, new_n1237,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n202), .A2(G50), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n208), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n211), .B1(new_n215), .B2(new_n216), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XNOR2_X1  g0033(.A(G50), .B(G68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT64), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G58), .B(G77), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G351));
  INV_X1    g0042(.A(G1), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G20), .ZN(new_n244));
  XOR2_X1   g0044(.A(KEYINPUT8), .B(G58), .Z(new_n245));
  INV_X1    g0045(.A(KEYINPUT71), .ZN(new_n246));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(KEYINPUT69), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT69), .ZN(new_n249));
  NAND4_X1  g0049(.A1(new_n249), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n248), .A2(new_n212), .A3(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT70), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g0053(.A1(new_n248), .A2(new_n250), .A3(KEYINPUT70), .A4(new_n212), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G13), .ZN(new_n256));
  NOR3_X1   g0056(.A1(new_n256), .A2(new_n213), .A3(G1), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n246), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  AOI211_X1 g0059(.A(KEYINPUT71), .B(new_n257), .C1(new_n253), .C2(new_n254), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n244), .B(new_n245), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT16), .ZN(new_n262));
  AND2_X1   g0062(.A1(G58), .A2(G68), .ZN(new_n263));
  OAI21_X1  g0063(.A(G20), .B1(new_n263), .B2(new_n201), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT81), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT81), .ZN(new_n266));
  OAI211_X1 g0066(.A(new_n266), .B(G20), .C1(new_n263), .C2(new_n201), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(G20), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G159), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G68), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT7), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n273), .B1(new_n274), .B2(G20), .ZN(new_n275));
  AND2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n272), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n262), .B1(new_n271), .B2(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(G1), .A2(G13), .ZN(new_n282));
  AND3_X1   g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n282), .B1(new_n283), .B2(new_n249), .ZN(new_n284));
  AOI21_X1  g0084(.A(KEYINPUT70), .B1(new_n284), .B2(new_n248), .ZN(new_n285));
  INV_X1    g0085(.A(new_n254), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(KEYINPUT7), .B1(new_n278), .B2(new_n213), .ZN(new_n288));
  NOR4_X1   g0088(.A1(new_n276), .A2(new_n277), .A3(new_n273), .A4(G20), .ZN(new_n289));
  OAI21_X1  g0089(.A(G68), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n265), .A2(new_n267), .B1(G159), .B2(new_n269), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT16), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n281), .A2(new_n287), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n245), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n257), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n261), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G87), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT82), .ZN(new_n298));
  OAI211_X1 g0098(.A(G226), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n299));
  INV_X1    g0099(.A(G1698), .ZN(new_n300));
  OAI211_X1 g0100(.A(G223), .B(new_n300), .C1(new_n276), .C2(new_n277), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n298), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n303));
  INV_X1    g0103(.A(G33), .ZN(new_n304));
  INV_X1    g0104(.A(G41), .ZN(new_n305));
  OAI211_X1 g0105(.A(G1), .B(G13), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n243), .B1(G41), .B2(G45), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n302), .A2(new_n303), .B1(G232), .B2(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n306), .A2(G274), .ZN(new_n310));
  OR2_X1    g0110(.A1(KEYINPUT66), .A2(G45), .ZN(new_n311));
  NAND2_X1  g0111(.A1(KEYINPUT66), .A2(G45), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(new_n305), .A3(new_n312), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n313), .A2(KEYINPUT67), .A3(new_n243), .ZN(new_n314));
  AOI21_X1  g0114(.A(KEYINPUT67), .B1(new_n313), .B2(new_n243), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n310), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(G169), .B1(new_n309), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G179), .ZN(new_n318));
  AND2_X1   g0118(.A1(new_n309), .A2(new_n316), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n296), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT18), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n296), .A2(KEYINPUT83), .A3(KEYINPUT18), .A4(new_n320), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n309), .A2(new_n316), .A3(new_n318), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(new_n319), .B2(G169), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n290), .A2(new_n291), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n255), .B1(new_n328), .B2(new_n262), .ZN(new_n329));
  AOI22_X1  g0129(.A1(new_n329), .A2(new_n292), .B1(new_n257), .B2(new_n294), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n327), .B1(new_n330), .B2(new_n261), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT83), .B1(new_n331), .B2(KEYINPUT18), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n325), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G190), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n309), .A2(new_n316), .A3(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n319), .B2(G200), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n336), .A2(new_n261), .A3(new_n293), .A4(new_n295), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT17), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n333), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n274), .A2(G232), .A3(G1698), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G33), .A2(G97), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n342), .B(KEYINPUT78), .ZN(new_n343));
  OAI211_X1 g0143(.A(G226), .B(new_n300), .C1(new_n276), .C2(new_n277), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n303), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n308), .A2(G238), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n316), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT13), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT13), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n316), .A2(new_n346), .A3(new_n350), .A4(new_n347), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G190), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n272), .A2(G20), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n213), .A2(G33), .ZN(new_n356));
  INV_X1    g0156(.A(G77), .ZN(new_n357));
  INV_X1    g0157(.A(new_n269), .ZN(new_n358));
  INV_X1    g0158(.A(G50), .ZN(new_n359));
  OAI221_X1 g0159(.A(new_n355), .B1(new_n356), .B2(new_n357), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n287), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT11), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(KEYINPUT79), .B1(new_n257), .B2(new_n272), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT12), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n287), .A2(KEYINPUT11), .A3(new_n360), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n255), .A2(G68), .A3(new_n244), .A4(new_n258), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n363), .A2(new_n365), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n352), .A2(G200), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n354), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G169), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(new_n349), .B2(new_n351), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT14), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n353), .A2(G179), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT80), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT67), .ZN(new_n377));
  AND2_X1   g0177(.A1(KEYINPUT66), .A2(G45), .ZN(new_n378));
  NOR2_X1   g0178(.A1(KEYINPUT66), .A2(G45), .ZN(new_n379));
  NOR3_X1   g0179(.A1(new_n378), .A2(new_n379), .A3(G41), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n377), .B1(new_n380), .B2(G1), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n313), .A2(KEYINPUT67), .A3(new_n243), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n383), .A2(new_n310), .B1(G238), .B2(new_n308), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n350), .B1(new_n384), .B2(new_n346), .ZN(new_n385));
  INV_X1    g0185(.A(new_n351), .ZN(new_n386));
  OAI21_X1  g0186(.A(G169), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n376), .B1(new_n387), .B2(KEYINPUT14), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n373), .A2(KEYINPUT80), .A3(new_n374), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n375), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n371), .B1(new_n390), .B2(new_n368), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n274), .A2(G232), .A3(new_n300), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n274), .A2(G238), .A3(G1698), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n278), .A2(G107), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT72), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT72), .A4(new_n394), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n397), .A2(new_n303), .A3(new_n398), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n383), .A2(new_n310), .B1(G244), .B2(new_n308), .ZN(new_n400));
  AOI21_X1  g0200(.A(G169), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n245), .A2(new_n269), .B1(G20), .B2(G77), .ZN(new_n403));
  XOR2_X1   g0203(.A(KEYINPUT15), .B(G87), .Z(new_n404));
  NAND4_X1  g0204(.A1(new_n404), .A2(KEYINPUT73), .A3(new_n213), .A4(G33), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT73), .ZN(new_n406));
  XNOR2_X1  g0206(.A(KEYINPUT15), .B(G87), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n406), .B1(new_n407), .B2(new_n356), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n403), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n409), .A2(new_n287), .B1(new_n357), .B2(new_n257), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n255), .A2(G77), .A3(new_n244), .A4(new_n258), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n402), .A2(KEYINPUT74), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT74), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n410), .A2(new_n411), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(new_n401), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n399), .A2(new_n400), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n417), .A2(G179), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n413), .A2(new_n416), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(G226), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n306), .A2(new_n307), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n316), .B(KEYINPUT68), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT68), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n306), .A2(G274), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n381), .B2(new_n382), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n422), .A2(new_n421), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n424), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n274), .A2(G222), .A3(new_n300), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n274), .A2(G223), .A3(G1698), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n429), .B(new_n430), .C1(new_n357), .C2(new_n274), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n303), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n423), .A2(new_n428), .A3(new_n432), .ZN(new_n433));
  OR2_X1    g0233(.A1(new_n433), .A2(G179), .ZN(new_n434));
  OAI211_X1 g0234(.A(G50), .B(new_n244), .C1(new_n259), .C2(new_n260), .ZN(new_n435));
  OAI21_X1  g0235(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n436));
  INV_X1    g0236(.A(G150), .ZN(new_n437));
  OAI221_X1 g0237(.A(new_n436), .B1(new_n437), .B2(new_n358), .C1(new_n294), .C2(new_n356), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n438), .A2(new_n287), .B1(new_n359), .B2(new_n257), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n433), .A2(new_n372), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n434), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n417), .A2(new_n334), .ZN(new_n443));
  INV_X1    g0243(.A(G200), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n444), .B1(new_n399), .B2(new_n400), .ZN(new_n445));
  OR3_X1    g0245(.A1(new_n443), .A2(new_n412), .A3(new_n445), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n420), .A2(new_n442), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n340), .A2(new_n391), .A3(new_n447), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n433), .A2(G200), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n433), .A2(new_n334), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n440), .A2(KEYINPUT9), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT9), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n435), .A2(new_n453), .A3(new_n439), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(KEYINPUT10), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n455), .A2(KEYINPUT75), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT75), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n452), .A2(new_n460), .A3(new_n454), .ZN(new_n461));
  XNOR2_X1  g0261(.A(KEYINPUT76), .B(KEYINPUT10), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n449), .A2(new_n450), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n459), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT77), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n459), .A2(new_n461), .A3(KEYINPUT77), .A4(new_n463), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n458), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n448), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n243), .A2(G33), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n258), .B(new_n471), .C1(new_n285), .C2(new_n286), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT87), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n255), .A2(KEYINPUT87), .A3(new_n258), .A4(new_n471), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n474), .A2(G87), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n274), .A2(G244), .A3(G1698), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G116), .ZN(new_n478));
  OAI211_X1 g0278(.A(G238), .B(new_n300), .C1(new_n276), .C2(new_n277), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n303), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n243), .A2(G45), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n306), .A2(G250), .A3(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n425), .B2(new_n482), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n481), .A2(new_n485), .A3(new_n334), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n484), .B1(new_n303), .B2(new_n480), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n486), .B1(G200), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT19), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n213), .B1(new_n343), .B2(new_n489), .ZN(new_n490));
  XNOR2_X1  g0290(.A(KEYINPUT84), .B(G97), .ZN(new_n491));
  INV_X1    g0291(.A(G87), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n491), .A2(new_n492), .A3(new_n205), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n204), .A2(KEYINPUT84), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT84), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G97), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT19), .B1(new_n498), .B2(G33), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n278), .A2(G20), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(G68), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n494), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n502), .A2(new_n287), .B1(new_n257), .B2(new_n407), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n476), .A2(new_n488), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n481), .A2(new_n485), .A3(new_n318), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(G169), .B2(new_n487), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n474), .A2(new_n404), .A3(new_n475), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(G45), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(G1), .ZN(new_n511));
  NAND2_X1  g0311(.A1(KEYINPUT5), .A2(G41), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(KEYINPUT5), .A2(G41), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n515), .A2(G257), .A3(new_n306), .ZN(new_n516));
  OAI211_X1 g0316(.A(G244), .B(new_n300), .C1(new_n276), .C2(new_n277), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT4), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n274), .A2(KEYINPUT4), .A3(G244), .A4(new_n300), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G283), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n274), .A2(G250), .A3(G1698), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n519), .A2(new_n520), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n516), .B1(new_n523), .B2(new_n303), .ZN(new_n524));
  OR2_X1    g0324(.A1(KEYINPUT5), .A2(G41), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n512), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n526), .A2(new_n306), .A3(G274), .A4(new_n511), .ZN(new_n527));
  AOI21_X1  g0327(.A(G169), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n527), .ZN(new_n529));
  AOI211_X1 g0329(.A(new_n529), .B(new_n516), .C1(new_n523), .C2(new_n303), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n528), .B1(new_n318), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n258), .A2(G97), .ZN(new_n532));
  AND2_X1   g0332(.A1(G97), .A2(G107), .ZN(new_n533));
  NOR2_X1   g0333(.A1(G97), .A2(G107), .ZN(new_n534));
  OAI21_X1  g0334(.A(KEYINPUT86), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT86), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G97), .A2(G107), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n206), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT6), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT85), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n498), .A2(new_n541), .A3(KEYINPUT6), .A4(new_n205), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n205), .A2(KEYINPUT6), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT85), .B1(new_n491), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n540), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G20), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n269), .A2(G77), .ZN(new_n547));
  OAI21_X1  g0347(.A(G107), .B1(new_n288), .B2(new_n289), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n532), .B1(new_n549), .B2(new_n287), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n474), .A2(G97), .A3(new_n475), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n531), .A2(new_n552), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n524), .A2(new_n334), .A3(new_n527), .ZN(new_n554));
  AOI21_X1  g0354(.A(G200), .B1(new_n524), .B2(new_n527), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n550), .B(new_n551), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n474), .A2(G107), .A3(new_n475), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n257), .A2(new_n205), .ZN(new_n558));
  XNOR2_X1  g0358(.A(new_n558), .B(KEYINPUT25), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n492), .A2(KEYINPUT89), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n560), .B(new_n213), .C1(new_n277), .C2(new_n276), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT22), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n274), .A2(KEYINPUT22), .A3(new_n213), .A4(new_n560), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n478), .A2(G20), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT23), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n213), .B2(G107), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n205), .A2(KEYINPUT23), .A3(G20), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n565), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n563), .A2(new_n564), .A3(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT24), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n255), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT24), .A4(new_n569), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n559), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n515), .A2(G264), .A3(new_n306), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n527), .ZN(new_n576));
  OAI211_X1 g0376(.A(G257), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n577));
  OAI211_X1 g0377(.A(G250), .B(new_n300), .C1(new_n276), .C2(new_n277), .ZN(new_n578));
  INV_X1    g0378(.A(G294), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n577), .B(new_n578), .C1(new_n304), .C2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n576), .B1(new_n303), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(G190), .ZN(new_n582));
  AND2_X1   g0382(.A1(new_n575), .A2(new_n527), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n580), .A2(new_n303), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G200), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n557), .A2(new_n574), .A3(new_n582), .A4(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n509), .A2(new_n553), .A3(new_n556), .A4(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(G116), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G20), .ZN(new_n590));
  AOI21_X1  g0390(.A(G33), .B1(new_n495), .B2(new_n497), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n521), .A2(new_n213), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n251), .B(new_n590), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT20), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n213), .B(new_n521), .C1(new_n491), .C2(G33), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n596), .A2(KEYINPUT20), .A3(new_n251), .A4(new_n590), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n255), .A2(G116), .A3(new_n258), .A4(new_n471), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n257), .A2(new_n589), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n482), .B1(new_n525), .B2(new_n512), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n602), .A2(new_n303), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n603), .A2(G270), .B1(new_n310), .B2(new_n602), .ZN(new_n604));
  OAI211_X1 g0404(.A(G264), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n605));
  OAI211_X1 g0405(.A(G257), .B(new_n300), .C1(new_n276), .C2(new_n277), .ZN(new_n606));
  INV_X1    g0406(.A(G303), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n605), .B(new_n606), .C1(new_n607), .C2(new_n274), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n303), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n372), .B1(new_n604), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n601), .A2(KEYINPUT21), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT88), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT88), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n601), .A2(new_n613), .A3(KEYINPUT21), .A4(new_n610), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n557), .A2(new_n574), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n581), .A2(G169), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n585), .A2(G179), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n601), .A2(new_n610), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT21), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n604), .A2(G179), .A3(new_n609), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n621), .A2(new_n622), .B1(new_n601), .B2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n601), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n604), .A2(new_n609), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(G200), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n625), .B(new_n627), .C1(new_n334), .C2(new_n626), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n615), .A2(new_n620), .A3(new_n624), .A4(new_n628), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n470), .A2(new_n588), .A3(new_n629), .ZN(G372));
  INV_X1    g0430(.A(new_n442), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n463), .A2(new_n461), .ZN(new_n632));
  AOI21_X1  g0432(.A(KEYINPUT77), .B1(new_n632), .B2(new_n459), .ZN(new_n633));
  INV_X1    g0433(.A(new_n467), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n457), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n331), .A2(KEYINPUT18), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n323), .ZN(new_n637));
  INV_X1    g0437(.A(new_n420), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n354), .A2(new_n369), .A3(new_n370), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n390), .A2(new_n368), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n637), .B1(new_n640), .B2(new_n339), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n631), .B1(new_n635), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n549), .A2(new_n287), .ZN(new_n643));
  INV_X1    g0443(.A(new_n532), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n643), .A2(new_n551), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n524), .A2(new_n318), .A3(new_n527), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n530), .B2(G169), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n556), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n507), .A2(new_n503), .ZN(new_n649));
  INV_X1    g0449(.A(new_n506), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n476), .A2(new_n488), .A3(new_n503), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(new_n652), .A3(new_n587), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT90), .ZN(new_n655));
  AND3_X1   g0455(.A1(new_n616), .A2(new_n619), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n655), .B1(new_n616), .B2(new_n619), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n615), .B(new_n624), .C1(new_n656), .C2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(KEYINPUT91), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n651), .A2(new_n552), .A3(new_n531), .A4(new_n652), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n647), .B1(new_n551), .B2(new_n550), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n509), .A2(KEYINPUT26), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n663), .A2(new_n665), .A3(KEYINPUT93), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT91), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n654), .A2(new_n658), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT93), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n661), .A2(new_n669), .A3(new_n662), .ZN(new_n670));
  XNOR2_X1  g0470(.A(new_n651), .B(KEYINPUT92), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n660), .A2(new_n666), .A3(new_n668), .A4(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n642), .B1(new_n470), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT94), .ZN(G369));
  NAND2_X1  g0476(.A1(new_n615), .A2(new_n624), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n243), .A2(new_n213), .A3(G13), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G213), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n625), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n677), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n615), .A2(new_n624), .A3(new_n628), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n686), .B1(new_n687), .B2(new_n685), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(G330), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n616), .A2(new_n683), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n620), .A2(new_n691), .A3(new_n587), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n693), .B1(new_n620), .B2(new_n684), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n683), .B(KEYINPUT95), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n656), .A2(new_n657), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n683), .B1(new_n615), .B2(new_n624), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n698), .B1(new_n699), .B2(new_n692), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n695), .A2(new_n700), .ZN(G399));
  NOR2_X1   g0501(.A1(new_n493), .A2(G116), .ZN(new_n702));
  INV_X1    g0502(.A(new_n209), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n705), .A3(G1), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n216), .B2(new_n705), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT96), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n615), .A2(new_n620), .A3(new_n624), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n709), .B1(new_n711), .B2(new_n588), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n654), .A2(KEYINPUT96), .A3(new_n710), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n508), .B(KEYINPUT92), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n714), .B1(new_n663), .B2(new_n665), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(KEYINPUT29), .A3(new_n684), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n654), .A2(new_n658), .A3(new_n667), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n667), .B1(new_n654), .B2(new_n658), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n666), .A2(new_n671), .A3(new_n670), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n697), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n717), .B1(new_n722), .B2(KEYINPUT29), .ZN(new_n723));
  INV_X1    g0523(.A(new_n687), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n724), .A2(new_n654), .A3(new_n620), .A4(new_n696), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT31), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n623), .A2(new_n524), .A3(new_n487), .A4(new_n581), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(KEYINPUT30), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n481), .A2(new_n485), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n585), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT30), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n730), .A2(new_n731), .A3(new_n524), .A4(new_n623), .ZN(new_n732));
  INV_X1    g0532(.A(new_n530), .ZN(new_n733));
  AND4_X1   g0533(.A1(new_n318), .A2(new_n626), .A3(new_n729), .A4(new_n585), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n728), .A2(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n726), .B1(new_n735), .B2(new_n684), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n728), .A2(new_n732), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n734), .A2(new_n733), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n697), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n725), .A2(new_n736), .A3(new_n740), .ZN(new_n741));
  AND2_X1   g0541(.A1(new_n741), .A2(G330), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n723), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n708), .B1(new_n745), .B2(G1), .ZN(G364));
  NOR2_X1   g0546(.A1(new_n256), .A2(G20), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n243), .B1(new_n747), .B2(G45), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n704), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n690), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(G330), .B2(new_n688), .ZN(new_n752));
  INV_X1    g0552(.A(new_n750), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT97), .ZN(new_n754));
  NAND2_X1  g0554(.A1(G355), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n206), .A2(KEYINPUT97), .A3(G87), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n755), .A2(new_n209), .A3(new_n274), .A4(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n237), .A2(new_n510), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n703), .A2(new_n274), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n311), .A2(new_n312), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n759), .B1(new_n216), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT98), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n757), .B1(G116), .B2(new_n209), .C1(new_n758), .C2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n212), .B1(G20), .B2(new_n372), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT99), .Z(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AND2_X1   g0570(.A1(new_n763), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(G20), .A2(G179), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n772), .B(KEYINPUT100), .Z(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n334), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n444), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(G200), .ZN(new_n776));
  AOI22_X1  g0576(.A1(G68), .A2(new_n775), .B1(new_n776), .B2(G77), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n773), .A2(G190), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n444), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G58), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n778), .A2(G200), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n777), .B1(new_n359), .B2(new_n780), .C1(new_n781), .C2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n213), .A2(G179), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n785), .A2(new_n334), .A3(G200), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n205), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n785), .A2(new_n334), .A3(new_n444), .ZN(new_n788));
  INV_X1    g0588(.A(G159), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n787), .B1(new_n791), .B2(KEYINPUT32), .ZN(new_n792));
  NOR3_X1   g0592(.A1(new_n334), .A2(G179), .A3(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n213), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n278), .B1(new_n795), .B2(G97), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT32), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n785), .A2(G190), .A3(G200), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n790), .A2(new_n797), .B1(new_n799), .B2(G87), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n792), .A2(new_n796), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n776), .A2(G311), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n795), .A2(G294), .ZN(new_n803));
  INV_X1    g0603(.A(new_n788), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n274), .B1(new_n804), .B2(G329), .ZN(new_n805));
  INV_X1    g0605(.A(new_n786), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n799), .A2(G303), .B1(new_n806), .B2(G283), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n802), .A2(new_n803), .A3(new_n805), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n779), .A2(G326), .ZN(new_n809));
  INV_X1    g0609(.A(G322), .ZN(new_n810));
  INV_X1    g0610(.A(new_n775), .ZN(new_n811));
  XOR2_X1   g0611(.A(KEYINPUT33), .B(G317), .Z(new_n812));
  OAI221_X1 g0612(.A(new_n809), .B1(new_n783), .B2(new_n810), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n784), .A2(new_n801), .B1(new_n808), .B2(new_n813), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n753), .B(new_n771), .C1(new_n767), .C2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n766), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n688), .B2(new_n816), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n752), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(G396));
  NOR2_X1   g0619(.A1(new_n415), .A2(new_n684), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n420), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n820), .B1(new_n420), .B2(new_n446), .ZN(new_n822));
  NOR3_X1   g0622(.A1(new_n821), .A2(new_n822), .A3(new_n697), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n673), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n821), .A2(new_n822), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n722), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n750), .B1(new_n826), .B2(new_n743), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n743), .B2(new_n826), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n767), .A2(new_n764), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n753), .B1(new_n357), .B2(new_n829), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G294), .A2(new_n782), .B1(new_n779), .B2(G303), .ZN(new_n831));
  INV_X1    g0631(.A(G283), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n831), .B1(new_n832), .B2(new_n811), .ZN(new_n833));
  INV_X1    g0633(.A(new_n776), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(new_n589), .ZN(new_n835));
  INV_X1    g0635(.A(G311), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n278), .B1(new_n788), .B2(new_n836), .C1(new_n794), .C2(new_n204), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n492), .A2(new_n786), .B1(new_n798), .B2(new_n205), .ZN(new_n838));
  NOR4_X1   g0638(.A1(new_n833), .A2(new_n835), .A3(new_n837), .A4(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(G143), .A2(new_n782), .B1(new_n776), .B2(G159), .ZN(new_n840));
  INV_X1    g0640(.A(G137), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n840), .B1(new_n841), .B2(new_n780), .C1(new_n437), .C2(new_n811), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT34), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n795), .A2(G58), .B1(new_n799), .B2(G50), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n278), .B1(new_n804), .B2(G132), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n844), .B(new_n845), .C1(new_n272), .C2(new_n786), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n846), .B(KEYINPUT101), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n839), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n767), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n830), .B1(new_n848), .B2(new_n849), .C1(new_n825), .C2(new_n765), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n828), .A2(new_n850), .ZN(G384));
  AOI211_X1 g0651(.A(new_n589), .B(new_n215), .C1(new_n545), .C2(KEYINPUT35), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(KEYINPUT35), .B2(new_n545), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT36), .Z(new_n854));
  OR3_X1    g0654(.A1(new_n216), .A2(new_n357), .A3(new_n263), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n359), .A2(G68), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT102), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n243), .B(G13), .C1(new_n855), .C2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n681), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n296), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n321), .A2(new_n861), .A3(new_n337), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n862), .A2(KEYINPUT37), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(KEYINPUT103), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT103), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n862), .A2(new_n865), .A3(KEYINPUT37), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT37), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n321), .A2(new_n861), .A3(new_n867), .A4(new_n337), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n868), .A2(KEYINPUT104), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(KEYINPUT104), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n864), .B(new_n866), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n861), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n333), .B2(new_n339), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n871), .A2(KEYINPUT38), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT38), .B1(new_n871), .B2(new_n873), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT39), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n374), .B(G169), .C1(new_n385), .C2(new_n386), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n349), .A2(G179), .A3(new_n351), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n387), .A2(new_n376), .A3(KEYINPUT14), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT80), .B1(new_n373), .B2(new_n374), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NOR3_X1   g0683(.A1(new_n883), .A2(new_n369), .A3(new_n683), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n871), .A2(new_n873), .A3(KEYINPUT38), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  AND2_X1   g0687(.A1(new_n321), .A2(new_n337), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT104), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n888), .A2(new_n889), .A3(new_n867), .A4(new_n861), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n868), .A2(KEYINPUT104), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n890), .A2(new_n891), .B1(KEYINPUT37), .B2(new_n862), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n861), .B1(new_n338), .B2(new_n637), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n887), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT39), .B1(new_n886), .B2(new_n894), .ZN(new_n895));
  NOR3_X1   g0695(.A1(new_n877), .A2(new_n885), .A3(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n368), .B(new_n683), .C1(new_n390), .C2(new_n371), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n368), .A2(new_n683), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n639), .B(new_n898), .C1(new_n883), .C2(new_n369), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n825), .A2(new_n696), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n720), .B2(new_n721), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n420), .A2(new_n683), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n874), .A2(new_n875), .ZN(new_n905));
  OAI22_X1  g0705(.A1(new_n904), .A2(new_n905), .B1(new_n637), .B2(new_n860), .ZN(new_n906));
  OR2_X1    g0706(.A1(new_n896), .A2(new_n906), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n469), .B(new_n717), .C1(new_n722), .C2(KEYINPUT29), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n642), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n907), .B(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n725), .A2(new_n736), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n469), .A2(new_n912), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n913), .B(KEYINPUT105), .Z(new_n914));
  NAND3_X1  g0714(.A1(new_n912), .A2(new_n900), .A3(new_n825), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n886), .B2(new_n894), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT40), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n912), .A2(new_n900), .A3(new_n917), .A4(new_n825), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n916), .A2(new_n917), .B1(new_n905), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n914), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n914), .A2(new_n920), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(G330), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n910), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n243), .B2(new_n747), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n910), .A2(new_n923), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n859), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n927), .B(KEYINPUT106), .Z(G367));
  OAI211_X1 g0728(.A(new_n553), .B(new_n556), .C1(new_n645), .C2(new_n696), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n929), .A2(new_n620), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n697), .B1(new_n930), .B2(new_n553), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n664), .A2(new_n697), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n933), .A2(new_n692), .A3(new_n699), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n931), .B1(new_n934), .B2(KEYINPUT42), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(KEYINPUT42), .B2(new_n934), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n476), .A2(new_n503), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n683), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n509), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n671), .B2(new_n938), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n936), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n942), .B(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n933), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n695), .A2(new_n946), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n945), .B(new_n947), .Z(new_n948));
  NAND2_X1  g0748(.A1(new_n700), .A2(new_n933), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT45), .Z(new_n950));
  NOR2_X1   g0750(.A1(new_n700), .A2(new_n933), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT44), .ZN(new_n952));
  AND3_X1   g0752(.A1(new_n950), .A2(new_n695), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n695), .B1(new_n950), .B2(new_n952), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n689), .A2(KEYINPUT107), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n699), .A2(new_n692), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n694), .B2(new_n699), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n956), .B(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n744), .B1(new_n955), .B2(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n704), .B(KEYINPUT41), .Z(new_n961));
  OAI21_X1  g0761(.A(new_n748), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n948), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n759), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n770), .B1(new_n209), .B2(new_n407), .C1(new_n232), .C2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n753), .B1(new_n965), .B2(KEYINPUT108), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(KEYINPUT108), .B2(new_n965), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n799), .A2(G116), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT46), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT109), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n782), .A2(G303), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n971), .B2(new_n970), .C1(new_n832), .C2(new_n834), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n274), .B1(new_n804), .B2(G317), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n491), .B2(new_n786), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G107), .B2(new_n795), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n969), .B2(new_n968), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n579), .A2(new_n811), .B1(new_n780), .B2(new_n836), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n973), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n794), .A2(new_n272), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n274), .B1(new_n788), .B2(new_n841), .C1(new_n357), .C2(new_n786), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n980), .B(new_n981), .C1(G58), .C2(new_n799), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n437), .B2(new_n783), .ZN(new_n983));
  AOI22_X1  g0783(.A1(G143), .A2(new_n779), .B1(new_n775), .B2(G159), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n359), .B2(new_n834), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n979), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT47), .Z(new_n988));
  AOI21_X1  g0788(.A(new_n967), .B1(new_n988), .B2(new_n767), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n940), .B2(new_n816), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n963), .A2(new_n990), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n991), .A2(KEYINPUT110), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(KEYINPUT110), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n992), .A2(new_n993), .ZN(G387));
  OR2_X1    g0794(.A1(new_n694), .A2(new_n816), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n229), .B1(new_n311), .B2(new_n312), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n274), .A2(new_n209), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n996), .A2(new_n964), .B1(new_n702), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(G45), .B1(G68), .B2(G77), .ZN(new_n999));
  AND3_X1   g0799(.A1(new_n245), .A2(KEYINPUT50), .A3(new_n359), .ZN(new_n1000));
  AOI21_X1  g0800(.A(KEYINPUT50), .B1(new_n245), .B2(new_n359), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n702), .B(new_n999), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n998), .A2(new_n1002), .B1(new_n205), .B2(new_n703), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n750), .B1(new_n1003), .B2(new_n769), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(G50), .A2(new_n782), .B1(new_n775), .B2(new_n245), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n776), .A2(G68), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n794), .A2(new_n407), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n274), .B1(new_n788), .B2(new_n437), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n786), .A2(new_n204), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n798), .A2(new_n357), .ZN(new_n1010));
  NOR4_X1   g0810(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n779), .A2(G159), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1005), .A2(new_n1006), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n274), .B1(new_n804), .B2(G326), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n794), .A2(new_n832), .B1(new_n798), .B2(new_n579), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G303), .A2(new_n776), .B1(new_n782), .B2(G317), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n836), .B2(new_n811), .C1(new_n810), .C2(new_n780), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT48), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n1018), .B2(new_n1017), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT49), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1014), .B1(new_n589), .B2(new_n786), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1013), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1004), .B1(new_n1024), .B2(new_n767), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n959), .A2(new_n749), .B1(new_n995), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n745), .A2(new_n959), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n704), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n745), .A2(new_n959), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1026), .B1(new_n1028), .B2(new_n1029), .ZN(G393));
  INV_X1    g0830(.A(new_n1027), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n705), .B1(new_n1031), .B2(new_n955), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n955), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n1027), .ZN(new_n1034));
  AND2_X1   g0834(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n770), .B1(new_n209), .B2(new_n491), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n241), .A2(new_n964), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n750), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n278), .B1(new_n788), .B2(new_n810), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n794), .A2(new_n589), .B1(new_n798), .B2(new_n832), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(G107), .C2(new_n806), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n607), .B2(new_n811), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G311), .A2(new_n782), .B1(new_n779), .B2(G317), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT52), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1042), .B(new_n1044), .C1(G294), .C2(new_n776), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1045), .A2(KEYINPUT113), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(KEYINPUT113), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G150), .A2(new_n779), .B1(new_n782), .B2(G159), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(KEYINPUT111), .B(KEYINPUT51), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n278), .B1(new_n804), .B2(G143), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1051), .B1(new_n272), .B2(new_n798), .C1(new_n492), .C2(new_n786), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT112), .Z(new_n1053));
  OAI22_X1  g0853(.A1(new_n834), .A2(new_n294), .B1(new_n357), .B2(new_n794), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G50), .B2(new_n775), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1050), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1046), .A2(new_n1047), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1038), .B1(new_n1057), .B2(new_n767), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n933), .B2(new_n816), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n1033), .B2(new_n748), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1035), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(G390));
  INV_X1    g0862(.A(KEYINPUT114), .ZN(new_n1063));
  NOR3_X1   g0863(.A1(new_n588), .A2(new_n629), .A3(new_n697), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n740), .A2(new_n736), .ZN(new_n1065));
  OAI211_X1 g0865(.A(G330), .B(new_n825), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  AND2_X1   g0866(.A1(new_n897), .A2(new_n899), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n716), .A2(new_n684), .A3(new_n825), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n903), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n900), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n884), .B1(new_n886), .B2(new_n894), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n886), .A2(new_n894), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n876), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n871), .A2(new_n873), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n887), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1077), .A2(KEYINPUT39), .A3(new_n886), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1075), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n903), .B1(new_n673), .B2(new_n823), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n885), .B1(new_n1080), .B2(new_n1067), .ZN(new_n1081));
  AOI221_X4 g0881(.A(new_n1068), .B1(new_n1072), .B2(new_n1073), .C1(new_n1079), .C2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n912), .A2(new_n900), .A3(G330), .A4(new_n825), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1081), .B1(new_n877), .B2(new_n895), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1083), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1063), .B1(new_n1082), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1068), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n895), .B1(new_n905), .B2(KEYINPUT39), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n824), .A2(new_n1070), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n884), .B1(new_n1090), .B2(new_n900), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1088), .B(new_n1085), .C1(new_n1089), .C2(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n1079), .A2(new_n1081), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1092), .B(KEYINPUT114), .C1(new_n1093), .C2(new_n1083), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n911), .A2(new_n736), .ZN(new_n1095));
  OAI211_X1 g0895(.A(G330), .B(new_n825), .C1(new_n1064), .C2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n1067), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n1097), .A2(new_n1070), .A3(new_n1069), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1083), .A2(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1098), .A2(new_n1088), .B1(new_n1090), .B2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n469), .A2(G330), .A3(new_n912), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n908), .A2(new_n642), .A3(new_n1102), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1087), .A2(new_n1094), .A3(new_n1105), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1104), .B(new_n1092), .C1(new_n1093), .C2(new_n1083), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(KEYINPUT115), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1087), .A2(KEYINPUT115), .A3(new_n1094), .A4(new_n1105), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n704), .A3(new_n1110), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(G283), .A2(new_n779), .B1(new_n776), .B2(new_n498), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n205), .B2(new_n811), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n783), .A2(new_n589), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n278), .B1(new_n788), .B2(new_n579), .C1(new_n492), .C2(new_n798), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n794), .A2(new_n357), .B1(new_n786), .B2(new_n272), .ZN(new_n1116));
  NOR4_X1   g0916(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1118), .A2(KEYINPUT117), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n278), .B1(new_n804), .B2(G125), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n1120), .B1(new_n359), .B2(new_n786), .C1(new_n789), .C2(new_n794), .ZN(new_n1121));
  INV_X1    g0921(.A(G128), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1122), .A2(new_n780), .B1(new_n811), .B2(new_n841), .ZN(new_n1123));
  INV_X1    g0923(.A(G132), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT54), .B(G143), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n1124), .A2(new_n783), .B1(new_n834), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n799), .A2(G150), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1127), .B(KEYINPUT53), .ZN(new_n1128));
  OR4_X1    g0928(.A1(new_n1121), .A2(new_n1123), .A3(new_n1126), .A4(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT117), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1129), .B1(new_n1117), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n767), .B1(new_n1119), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n829), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1132), .B(new_n750), .C1(new_n245), .C2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(new_n1079), .B2(new_n764), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1092), .B1(new_n1093), .B2(new_n1083), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT116), .ZN(new_n1137));
  OR3_X1    g0937(.A1(new_n1136), .A2(new_n1137), .A3(new_n748), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1137), .B1(new_n1136), .B2(new_n748), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1135), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1111), .A2(new_n1140), .ZN(G378));
  NAND2_X1  g0941(.A1(new_n440), .A2(new_n860), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n635), .A2(new_n442), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1142), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n468), .B2(new_n631), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1143), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n919), .B2(G330), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n912), .A2(new_n900), .A3(new_n825), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n917), .B1(new_n1074), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n918), .B1(new_n1077), .B2(new_n886), .ZN(new_n1155));
  OAI21_X1  g0955(.A(G330), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1143), .A2(new_n1145), .A3(new_n1147), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1147), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n907), .B1(new_n1152), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n896), .A2(new_n906), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1151), .A2(new_n919), .A3(G330), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1156), .A2(new_n1159), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1162), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n749), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n305), .B(new_n278), .C1(new_n788), .C2(new_n832), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n786), .A2(new_n781), .ZN(new_n1169));
  OR4_X1    g0969(.A1(new_n980), .A2(new_n1168), .A3(new_n1010), .A4(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G97), .A2(new_n775), .B1(new_n782), .B2(G107), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n589), .B2(new_n780), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(new_n404), .C2(new_n776), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1173), .A2(KEYINPUT58), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(KEYINPUT58), .ZN(new_n1175));
  AOI21_X1  g0975(.A(G50), .B1(new_n304), .B2(new_n305), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n274), .B2(G41), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT118), .Z(new_n1178));
  NAND2_X1  g0978(.A1(new_n1175), .A2(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n779), .A2(G125), .B1(G150), .B2(new_n795), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT119), .Z(new_n1181));
  OAI22_X1  g0981(.A1(new_n834), .A2(new_n841), .B1(new_n798), .B2(new_n1125), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n1122), .A2(new_n783), .B1(new_n811), .B2(new_n1124), .ZN(new_n1183));
  OR3_X1    g0983(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  OR2_X1    g0984(.A1(new_n1184), .A2(KEYINPUT59), .ZN(new_n1185));
  AOI211_X1 g0985(.A(G33), .B(G41), .C1(new_n804), .C2(G124), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n789), .B2(new_n786), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(new_n1184), .B2(KEYINPUT59), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1174), .B(new_n1179), .C1(new_n1185), .C2(new_n1188), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n750), .B1(G50), .B2(new_n1133), .C1(new_n1189), .C2(new_n849), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n1159), .B2(new_n764), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1167), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1103), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1165), .A2(new_n1161), .B1(new_n1107), .B2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n705), .B1(new_n1195), .B2(KEYINPUT57), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1107), .A2(new_n1194), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1166), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT57), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1193), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(G375));
  INV_X1    g1002(.A(new_n1101), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1203), .A2(new_n1194), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT120), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n961), .ZN(new_n1207));
  OAI21_X1  g1007(.A(KEYINPUT120), .B1(new_n1203), .B2(new_n1194), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1206), .A2(new_n1207), .A3(new_n1105), .A4(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1067), .A2(new_n764), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n750), .B1(G68), .B2(new_n1133), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n779), .A2(G132), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT123), .Z(new_n1213));
  INV_X1    g1013(.A(new_n1125), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G137), .A2(new_n782), .B1(new_n775), .B2(new_n1214), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n794), .A2(new_n359), .B1(new_n798), .B2(new_n789), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n274), .B1(new_n788), .B2(new_n1122), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1216), .A2(new_n1169), .A3(new_n1217), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1215), .B(new_n1218), .C1(new_n437), .C2(new_n834), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n278), .B1(new_n786), .B2(new_n357), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT121), .Z(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n205), .B2(new_n834), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G283), .A2(new_n782), .B1(new_n779), .B2(G294), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n798), .A2(new_n204), .B1(new_n788), .B2(new_n607), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT122), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1007), .B1(new_n775), .B2(G116), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1223), .A2(new_n1225), .A3(new_n1226), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n1213), .A2(new_n1219), .B1(new_n1222), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1211), .B1(new_n1228), .B2(new_n767), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1203), .A2(new_n749), .B1(new_n1210), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1209), .A2(new_n1230), .ZN(G381));
  INV_X1    g1031(.A(G384), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1061), .A2(new_n1232), .ZN(new_n1233));
  OR4_X1    g1033(.A1(G396), .A2(new_n1233), .A3(G393), .A4(G381), .ZN(new_n1234));
  OR4_X1    g1034(.A1(G387), .A2(new_n1234), .A3(G378), .A4(G375), .ZN(G407));
  NAND2_X1  g1035(.A1(new_n682), .A2(G213), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(G375), .A2(G378), .A3(new_n1236), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT124), .Z(new_n1238));
  NAND3_X1  g1038(.A1(new_n1238), .A2(G407), .A3(G213), .ZN(G409));
  NAND3_X1  g1039(.A1(new_n1166), .A2(new_n1197), .A3(new_n1207), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1240), .A2(new_n1167), .A3(new_n1192), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1111), .A2(new_n1241), .A3(new_n1140), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT125), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1201), .A2(G378), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT125), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1111), .A2(new_n1241), .A3(new_n1245), .A4(new_n1140), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(KEYINPUT126), .B1(new_n1204), .B2(KEYINPUT60), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1248), .A2(new_n705), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1105), .A2(KEYINPUT60), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1206), .A2(new_n1250), .A3(new_n1208), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1204), .A2(KEYINPUT126), .A3(KEYINPUT60), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1249), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(G384), .B1(new_n1253), .B2(new_n1230), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1253), .A2(G384), .A3(new_n1230), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1247), .A2(new_n1236), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(KEYINPUT62), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1247), .A2(new_n1236), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n682), .A2(G213), .A3(G2897), .ZN(new_n1262));
  AND3_X1   g1062(.A1(new_n1255), .A2(new_n1256), .A3(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1262), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1261), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT61), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT62), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1247), .A2(new_n1268), .A3(new_n1258), .A4(new_n1236), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1260), .A2(new_n1266), .A3(new_n1267), .A4(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n991), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(G390), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n991), .A2(new_n1061), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(G393), .B(G396), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT127), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1274), .A2(KEYINPUT127), .A3(new_n1276), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n992), .A2(new_n993), .A3(new_n1061), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1276), .B1(new_n1271), .B2(G390), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n1278), .A2(new_n1279), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1270), .A2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT61), .B1(new_n1261), .B2(new_n1265), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1274), .A2(KEYINPUT127), .A3(new_n1276), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1285), .B1(new_n1286), .B2(new_n1277), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT63), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1259), .A2(new_n1288), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1247), .A2(KEYINPUT63), .A3(new_n1258), .A4(new_n1236), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1284), .A2(new_n1287), .A3(new_n1289), .A4(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1283), .A2(new_n1291), .ZN(G405));
  OR2_X1    g1092(.A1(new_n1201), .A2(G378), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1244), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1258), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1293), .A2(new_n1257), .A3(new_n1244), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(new_n1282), .B(new_n1297), .ZN(G402));
endmodule


