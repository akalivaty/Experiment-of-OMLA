//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n447, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n569, new_n570, new_n571, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1166,
    new_n1167, new_n1168;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G220));
  XOR2_X1   g013(.A(KEYINPUT67), .B(G96), .Z(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  NAND2_X1  g021(.A1(G94), .A2(G452), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT68), .Z(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n453), .B(new_n454), .Z(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT70), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT70), .ZN(new_n468));
  OAI211_X1 g043(.A(new_n468), .B(G125), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  OAI211_X1 g048(.A(G137), .B(new_n473), .C1(new_n464), .C2(new_n465), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n473), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n472), .A2(new_n477), .ZN(G160));
  OR2_X1    g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n473), .B1(new_n479), .B2(new_n480), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G114), .C2(new_n473), .ZN(new_n490));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(G138), .B(new_n473), .C1(new_n464), .C2(new_n465), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n479), .A2(new_n480), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n473), .A2(G138), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n492), .B1(new_n494), .B2(new_n498), .ZN(G164));
  NAND2_X1  g074(.A1(G75), .A2(G543), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  INV_X1    g077(.A(G543), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT5), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT71), .A3(G543), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n504), .A2(new_n506), .B1(KEYINPUT5), .B2(new_n503), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n501), .B1(new_n507), .B2(G62), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  OAI21_X1  g084(.A(KEYINPUT72), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n503), .A2(KEYINPUT5), .ZN(new_n511));
  AND3_X1   g086(.A1(new_n505), .A2(KEYINPUT71), .A3(G543), .ZN(new_n512));
  AOI21_X1  g087(.A(KEYINPUT71), .B1(new_n505), .B2(G543), .ZN(new_n513));
  OAI211_X1 g088(.A(G62), .B(new_n511), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(new_n500), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(new_n516), .A3(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n504), .A2(new_n506), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT6), .B(G651), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n518), .A2(G88), .A3(new_n511), .A4(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n519), .A2(G50), .A3(G543), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n510), .A2(new_n517), .A3(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  AND2_X1   g099(.A1(new_n519), .A2(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  AND3_X1   g104(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n518), .A2(new_n511), .A3(new_n519), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G89), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(G168));
  AOI22_X1  g110(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n509), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n519), .A2(G543), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT73), .B(G52), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n531), .A2(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n537), .A2(new_n541), .ZN(G171));
  AOI22_X1  g117(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(KEYINPUT74), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(KEYINPUT74), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n544), .A2(G651), .A3(new_n545), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n532), .A2(G81), .B1(G43), .B2(new_n525), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(new_n549));
  XOR2_X1   g124(.A(new_n549), .B(KEYINPUT75), .Z(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT76), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(new_n555));
  XOR2_X1   g130(.A(new_n555), .B(KEYINPUT77), .Z(G188));
  AOI22_X1  g131(.A1(new_n507), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n557), .A2(new_n509), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT78), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n531), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n507), .A2(KEYINPUT78), .A3(new_n519), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n560), .A2(G91), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OR3_X1    g138(.A1(new_n539), .A2(KEYINPUT9), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT9), .B1(new_n539), .B2(new_n563), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n558), .A2(new_n562), .A3(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  NAND3_X1  g143(.A1(new_n530), .A2(KEYINPUT79), .A3(new_n533), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(KEYINPUT79), .B1(new_n530), .B2(new_n533), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n570), .A2(new_n571), .ZN(G286));
  OR2_X1    g147(.A1(new_n507), .A2(G74), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n573), .A2(G651), .B1(G49), .B2(new_n525), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n560), .A2(G87), .A3(new_n561), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(new_n525), .A2(G48), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n507), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n578), .B2(new_n509), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n560), .A2(G86), .A3(new_n561), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT80), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n560), .A2(new_n582), .A3(G86), .A4(new_n561), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n579), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G305));
  AOI22_X1  g160(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n509), .ZN(new_n587));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  INV_X1    g163(.A(G47), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n531), .A2(new_n588), .B1(new_n589), .B2(new_n539), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n587), .A2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(G301), .A2(G868), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT81), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n507), .A2(G66), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(G54), .B2(new_n525), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n560), .A2(KEYINPUT10), .A3(G92), .A4(new_n561), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT10), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n560), .A2(new_n561), .ZN(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n598), .B1(new_n599), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n593), .B1(G868), .B2(new_n604), .ZN(G284));
  OAI21_X1  g180(.A(new_n593), .B1(G868), .B2(new_n604), .ZN(G321));
  AOI21_X1  g181(.A(KEYINPUT82), .B1(G286), .B2(G868), .ZN(new_n607));
  INV_X1    g182(.A(G299), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(G868), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(G286), .A2(KEYINPUT82), .A3(G868), .ZN(new_n610));
  AND2_X1   g185(.A1(new_n609), .A2(new_n610), .ZN(G297));
  XNOR2_X1  g186(.A(G297), .B(KEYINPUT83), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n604), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n603), .A2(new_n599), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(new_n597), .ZN(new_n616));
  OAI21_X1  g191(.A(G868), .B1(new_n616), .B2(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n495), .A2(new_n475), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  INV_X1    g197(.A(G2100), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n481), .A2(G135), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n483), .A2(G123), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n473), .A2(G111), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n626), .B(new_n627), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(G2096), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n624), .A2(new_n625), .A3(new_n632), .ZN(G156));
  XOR2_X1   g208(.A(KEYINPUT15), .B(G2435), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT85), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2427), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT84), .B(G2438), .Z(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(new_n640), .A3(KEYINPUT14), .ZN(new_n641));
  XOR2_X1   g216(.A(G2451), .B(G2454), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n641), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  AND3_X1   g225(.A1(new_n649), .A2(G14), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT86), .Z(G401));
  INV_X1    g227(.A(KEYINPUT18), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n654), .A2(new_n655), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(new_n623), .ZN(new_n660));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n656), .B2(KEYINPUT18), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(new_n631), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(G1971), .B(G1976), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT20), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n668), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n666), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n666), .B2(new_n672), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n675), .B(new_n676), .Z(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1981), .B(G1986), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(G229));
  INV_X1    g257(.A(G16), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n683), .A2(G23), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(G288), .B2(G16), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT33), .ZN(new_n686));
  INV_X1    g261(.A(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n683), .A2(G6), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(new_n584), .B2(new_n683), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT32), .B(G1981), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  NOR2_X1   g268(.A1(G16), .A2(G22), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(G166), .B2(G16), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT89), .B(G1971), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  AND4_X1   g272(.A1(new_n688), .A2(new_n692), .A3(new_n693), .A4(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT34), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  MUX2_X1   g276(.A(G24), .B(G290), .S(G16), .Z(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G1986), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G25), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT87), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n481), .A2(G131), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n483), .A2(G119), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n473), .A2(G107), .ZN(new_n709));
  OAI21_X1  g284(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n710));
  OAI211_X1 g285(.A(new_n707), .B(new_n708), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n706), .B1(new_n711), .B2(G29), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT35), .B(G1991), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT88), .Z(new_n714));
  XOR2_X1   g289(.A(new_n712), .B(new_n714), .Z(new_n715));
  NOR2_X1   g290(.A1(new_n703), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n700), .A2(new_n701), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(KEYINPUT36), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT36), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n700), .A2(new_n719), .A3(new_n701), .A4(new_n716), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n704), .A2(G33), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT25), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n481), .A2(G139), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n495), .A2(G127), .ZN(new_n726));
  NAND2_X1  g301(.A1(G115), .A2(G2104), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n473), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n721), .B1(new_n730), .B2(new_n704), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n731), .A2(G2072), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT94), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n704), .A2(G26), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT92), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT28), .ZN(new_n736));
  AOI22_X1  g311(.A1(G128), .A2(new_n483), .B1(new_n481), .B2(G140), .ZN(new_n737));
  INV_X1    g312(.A(G104), .ZN(new_n738));
  AND3_X1   g313(.A1(new_n738), .A2(new_n473), .A3(KEYINPUT91), .ZN(new_n739));
  AOI21_X1  g314(.A(KEYINPUT91), .B1(new_n738), .B2(new_n473), .ZN(new_n740));
  OAI221_X1 g315(.A(G2104), .B1(G116), .B2(new_n473), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n736), .B1(new_n742), .B2(G29), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT93), .B(G2067), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT100), .B(KEYINPUT29), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G2090), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n704), .A2(G35), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT99), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n487), .B2(G29), .ZN(new_n750));
  OAI22_X1  g325(.A1(new_n743), .A2(new_n744), .B1(new_n747), .B2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G2078), .ZN(new_n752));
  NOR2_X1   g327(.A1(G164), .A2(new_n704), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G27), .B2(new_n704), .ZN(new_n754));
  AOI211_X1 g329(.A(new_n745), .B(new_n751), .C1(new_n752), .C2(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT30), .B(G28), .ZN(new_n756));
  OR2_X1    g331(.A1(KEYINPUT31), .A2(G11), .ZN(new_n757));
  NAND2_X1  g332(.A1(KEYINPUT31), .A2(G11), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n756), .A2(new_n704), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n630), .B2(new_n704), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n750), .A2(new_n747), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n754), .B2(new_n752), .ZN(new_n762));
  AOI211_X1 g337(.A(new_n760), .B(new_n762), .C1(G2072), .C2(new_n731), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n481), .A2(G141), .B1(G105), .B2(new_n475), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n483), .A2(G129), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT26), .Z(new_n767));
  NAND3_X1  g342(.A1(new_n764), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  MUX2_X1   g343(.A(G32), .B(new_n768), .S(G29), .Z(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT27), .B(G1996), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n733), .A2(new_n755), .A3(new_n763), .A4(new_n771), .ZN(new_n772));
  XOR2_X1   g347(.A(KEYINPUT95), .B(KEYINPUT24), .Z(new_n773));
  INV_X1    g348(.A(G34), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n704), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n774), .B2(new_n773), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT96), .Z(new_n777));
  INV_X1    g352(.A(G160), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n704), .B2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(G2084), .ZN(new_n780));
  OR2_X1    g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n683), .A2(G5), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G171), .B2(new_n683), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G1961), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n783), .A2(G1961), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n779), .A2(new_n780), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n781), .A2(new_n784), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n683), .A2(G19), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n548), .B2(new_n683), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1341), .ZN(new_n790));
  NOR3_X1   g365(.A1(new_n772), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n683), .A2(G4), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n604), .B2(new_n683), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT90), .B(G1348), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n683), .A2(G21), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G168), .B2(new_n683), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT97), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT98), .B(G1966), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n798), .B(new_n799), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n683), .A2(G20), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT23), .Z(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G299), .B2(G16), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT101), .B(G1956), .Z(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n791), .A2(new_n795), .A3(new_n800), .A4(new_n805), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(KEYINPUT102), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(KEYINPUT102), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n718), .A2(new_n720), .B1(new_n807), .B2(new_n808), .ZN(G311));
  INV_X1    g384(.A(G311), .ZN(G150));
  AOI22_X1  g385(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(new_n509), .ZN(new_n812));
  INV_X1    g387(.A(G93), .ZN(new_n813));
  INV_X1    g388(.A(G55), .ZN(new_n814));
  OAI22_X1  g389(.A1(new_n531), .A2(new_n813), .B1(new_n814), .B2(new_n539), .ZN(new_n815));
  OAI21_X1  g390(.A(G860), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT37), .Z(new_n817));
  NOR2_X1   g392(.A1(new_n616), .A2(new_n613), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT38), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n812), .A2(new_n815), .ZN(new_n820));
  AND3_X1   g395(.A1(new_n546), .A2(new_n547), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n820), .B1(new_n546), .B2(new_n547), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n819), .A2(new_n823), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n824), .A2(KEYINPUT39), .A3(new_n825), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT103), .Z(new_n827));
  AOI21_X1  g402(.A(KEYINPUT39), .B1(new_n824), .B2(new_n825), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n828), .A2(G860), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n827), .A2(KEYINPUT104), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(KEYINPUT104), .B1(new_n827), .B2(new_n829), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n817), .B1(new_n830), .B2(new_n831), .ZN(G145));
  NAND2_X1  g407(.A1(new_n483), .A2(G130), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n473), .A2(G118), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(G142), .B2(new_n481), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(new_n621), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n711), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT107), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n742), .B(new_n768), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n494), .A2(new_n498), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n490), .A2(new_n491), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n842), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT106), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n729), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n846), .A2(new_n848), .A3(new_n730), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n841), .B(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n630), .B(KEYINPUT105), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G160), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n487), .ZN(new_n856));
  AOI21_X1  g431(.A(G37), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT108), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n856), .B1(new_n841), .B2(new_n852), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n838), .B(new_n711), .Z(new_n860));
  NAND3_X1  g435(.A1(new_n850), .A2(new_n860), .A3(new_n851), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n858), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n859), .A2(new_n858), .A3(new_n861), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n857), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g440(.A1(new_n616), .A2(G559), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n823), .B(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n616), .A2(new_n608), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT109), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n604), .A2(new_n869), .A3(G299), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n869), .B1(new_n604), .B2(G299), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n868), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n867), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n604), .A2(G299), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT110), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n868), .A2(KEYINPUT110), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n877), .B(new_n878), .C1(new_n871), .C2(new_n872), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT41), .ZN(new_n880));
  INV_X1    g455(.A(new_n872), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n880), .B1(new_n881), .B2(new_n870), .ZN(new_n882));
  AOI22_X1  g457(.A1(new_n879), .A2(new_n880), .B1(new_n882), .B2(new_n868), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n874), .B1(new_n883), .B2(new_n867), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT111), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT42), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n584), .B(G166), .ZN(new_n887));
  INV_X1    g462(.A(G288), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(G290), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n887), .B(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT42), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n890), .B1(KEYINPUT111), .B2(new_n891), .ZN(new_n892));
  OAI221_X1 g467(.A(new_n874), .B1(KEYINPUT111), .B2(new_n891), .C1(new_n883), .C2(new_n867), .ZN(new_n893));
  AND3_X1   g468(.A1(new_n886), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n892), .B1(new_n886), .B2(new_n893), .ZN(new_n895));
  OAI21_X1  g470(.A(G868), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n896), .B1(G868), .B2(new_n820), .ZN(G295));
  OAI21_X1  g472(.A(new_n896), .B1(G868), .B2(new_n820), .ZN(G331));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n899));
  INV_X1    g474(.A(new_n821), .ZN(new_n900));
  INV_X1    g475(.A(new_n822), .ZN(new_n901));
  INV_X1    g476(.A(new_n571), .ZN(new_n902));
  AOI21_X1  g477(.A(G301), .B1(new_n902), .B2(new_n569), .ZN(new_n903));
  NOR2_X1   g478(.A1(G168), .A2(G171), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n900), .B(new_n901), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n904), .ZN(new_n906));
  OAI21_X1  g481(.A(G171), .B1(new_n570), .B2(new_n571), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n906), .B(new_n907), .C1(new_n822), .C2(new_n821), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n873), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT112), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n909), .A2(new_n873), .A3(KEYINPUT112), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n877), .A2(new_n878), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(new_n882), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n873), .A2(new_n880), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n909), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n890), .B1(new_n914), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(G37), .ZN(new_n920));
  INV_X1    g495(.A(new_n890), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n921), .B(new_n910), .C1(new_n883), .C2(new_n909), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n899), .B1(new_n923), .B2(KEYINPUT43), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n922), .A2(new_n920), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n879), .A2(new_n880), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n882), .A2(new_n868), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n909), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n910), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n890), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n926), .A2(KEYINPUT113), .A3(new_n927), .A4(new_n932), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n932), .A2(new_n927), .A3(new_n920), .A4(new_n922), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT113), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n924), .A2(new_n933), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n928), .A2(new_n929), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n905), .A2(new_n908), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n921), .B1(new_n940), .B2(new_n910), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT43), .B1(new_n925), .B2(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n919), .A2(new_n927), .A3(new_n920), .A4(new_n922), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n899), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n937), .A2(new_n945), .ZN(G397));
  AOI22_X1  g521(.A1(new_n466), .A2(KEYINPUT70), .B1(G113), .B2(G2104), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n473), .B1(new_n947), .B2(new_n469), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n474), .A2(new_n476), .A3(G40), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT114), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT114), .ZN(new_n951));
  INV_X1    g526(.A(new_n949), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n472), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n955));
  INV_X1    g530(.A(G1384), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n845), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT115), .ZN(new_n959));
  INV_X1    g534(.A(G2067), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n742), .B(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n768), .B(G1996), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XOR2_X1   g539(.A(new_n711), .B(new_n714), .Z(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(G290), .B(G1986), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n959), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT124), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n951), .B1(new_n472), .B2(new_n952), .ZN(new_n970));
  AOI211_X1 g545(.A(KEYINPUT114), .B(new_n949), .C1(new_n471), .C2(G2105), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n955), .B1(G164), .B2(G1384), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n845), .A2(KEYINPUT45), .A3(new_n956), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n799), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(G164), .B2(G1384), .ZN(new_n978));
  XOR2_X1   g553(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n845), .A2(new_n956), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT119), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n982), .A2(new_n954), .A3(new_n983), .A4(new_n780), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n976), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(G2084), .B1(new_n978), .B2(new_n981), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n983), .B1(new_n986), .B2(new_n954), .ZN(new_n987));
  OAI211_X1 g562(.A(KEYINPUT123), .B(G8), .C1(new_n985), .C2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G8), .ZN(new_n989));
  NOR2_X1   g564(.A1(G168), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(KEYINPUT51), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT50), .B1(new_n845), .B2(new_n956), .ZN(new_n993));
  AOI211_X1 g568(.A(G1384), .B(new_n979), .C1(new_n843), .C2(new_n844), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n780), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT119), .B1(new_n995), .B2(new_n972), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n996), .A2(new_n976), .A3(new_n984), .ZN(new_n997));
  AOI21_X1  g572(.A(KEYINPUT123), .B1(new_n997), .B2(G8), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n969), .B1(new_n992), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n997), .A2(G8), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT123), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n1002), .A2(KEYINPUT124), .A3(new_n988), .A4(new_n991), .ZN(new_n1003));
  OAI211_X1 g578(.A(KEYINPUT51), .B(G8), .C1(new_n997), .C2(new_n534), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n999), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT62), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n997), .A2(new_n990), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1006), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1009));
  NAND2_X1  g584(.A1(G303), .A2(G8), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n980), .B1(G164), .B2(G1384), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(new_n970), .B2(new_n971), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G2090), .ZN(new_n1019));
  INV_X1    g594(.A(new_n957), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n977), .ZN(new_n1021));
  OAI211_X1 g596(.A(KEYINPUT118), .B(new_n1015), .C1(new_n970), .C2(new_n971), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n973), .A2(new_n974), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1971), .B1(new_n1024), .B2(new_n954), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1014), .B1(new_n1027), .B2(G8), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT49), .ZN(new_n1029));
  AOI211_X1 g604(.A(G1981), .B(new_n579), .C1(new_n581), .C2(new_n583), .ZN(new_n1030));
  INV_X1    g605(.A(G1981), .ZN(new_n1031));
  INV_X1    g606(.A(new_n579), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n532), .A2(G86), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1029), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n584), .A2(new_n1031), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1034), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1036), .A2(KEYINPUT49), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n957), .B1(new_n950), .B2(new_n953), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1039), .A2(new_n989), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1035), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n982), .A2(new_n954), .A3(new_n1019), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1014), .B(G8), .C1(new_n1025), .C2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n888), .A2(G1976), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(KEYINPUT52), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT52), .B1(G288), .B2(new_n687), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1040), .A2(new_n1044), .A3(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1041), .A2(new_n1043), .A3(new_n1046), .A4(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1028), .A2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n954), .A2(new_n752), .A3(new_n973), .A4(new_n974), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1052), .A2(KEYINPUT125), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1024), .A2(new_n752), .A3(new_n954), .A4(new_n1053), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n982), .A2(new_n954), .ZN(new_n1057));
  INV_X1    g632(.A(G1961), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1055), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  AND3_X1   g635(.A1(new_n1060), .A2(KEYINPUT126), .A3(G171), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT126), .B1(new_n1060), .B2(G171), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1050), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n1008), .A2(new_n1009), .A3(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n752), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1024), .A2(G160), .A3(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1066), .A2(new_n1059), .A3(new_n1068), .ZN(new_n1069));
  OR2_X1    g644(.A1(new_n1069), .A2(G171), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT54), .B1(new_n1065), .B2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1055), .A2(G301), .A3(new_n1056), .A4(new_n1059), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT127), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1051), .A2(new_n1054), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1075), .A2(KEYINPUT127), .A3(G301), .A4(new_n1056), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1078), .B1(new_n1069), .B2(G171), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1050), .A2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1071), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT61), .ZN(new_n1084));
  INV_X1    g659(.A(G1956), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1022), .A2(new_n1021), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT118), .B1(new_n954), .B2(new_n1015), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n972), .A2(new_n975), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n1090), .B(G2072), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  XOR2_X1   g667(.A(G299), .B(KEYINPUT57), .Z(new_n1093));
  AND3_X1   g668(.A1(new_n1088), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1093), .B1(new_n1088), .B2(new_n1092), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1084), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1093), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n950), .A2(new_n953), .B1(new_n957), .B2(new_n980), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1098), .A2(KEYINPUT118), .B1(new_n977), .B2(new_n1020), .ZN(new_n1099));
  AOI21_X1  g674(.A(G1956), .B1(new_n1099), .B2(new_n1018), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1092), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1097), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1088), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n1103), .A3(KEYINPUT61), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n1105));
  XNOR2_X1  g680(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1106), .B(G1341), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1105), .B(new_n1107), .C1(new_n972), .C2(new_n957), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1107), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT122), .B1(new_n1039), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1996), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1024), .A2(new_n1111), .A3(new_n954), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1108), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n548), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT59), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(new_n1116), .A3(new_n548), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1057), .A2(new_n794), .B1(new_n960), .B2(new_n1039), .ZN(new_n1119));
  AND3_X1   g694(.A1(new_n1119), .A2(KEYINPUT60), .A3(new_n616), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n616), .B1(new_n1119), .B2(KEYINPUT60), .ZN(new_n1121));
  OAI22_X1  g696(.A1(new_n1120), .A2(new_n1121), .B1(KEYINPUT60), .B2(new_n1119), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1096), .A2(new_n1104), .A3(new_n1118), .A4(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1119), .A2(new_n616), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1095), .B1(new_n1103), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1082), .A2(new_n1083), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n687), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1128), .B(KEYINPUT117), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1129), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1040), .B1(new_n1130), .B2(new_n1030), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n1041), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1131), .B1(new_n1043), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1000), .A2(G286), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1050), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT63), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(G8), .B1(new_n1025), .B2(new_n1042), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1014), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1137), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1135), .A2(new_n1141), .ZN(new_n1142));
  OR2_X1    g717(.A1(new_n1142), .A2(new_n1049), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1134), .B1(new_n1138), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1127), .A2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n968), .B1(new_n1064), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n959), .B1(new_n768), .B2(new_n962), .ZN(new_n1147));
  INV_X1    g722(.A(new_n959), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1148), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT46), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1150), .B1(new_n959), .B2(new_n1111), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1147), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  XOR2_X1   g727(.A(new_n1152), .B(KEYINPUT47), .Z(new_n1153));
  NOR2_X1   g728(.A1(G290), .A2(G1986), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n959), .A2(KEYINPUT48), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n959), .A2(new_n966), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT48), .B1(new_n959), .B2(new_n1154), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n742), .A2(G2067), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n711), .A2(new_n714), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1159), .B1(new_n964), .B2(new_n1160), .ZN(new_n1161));
  OAI22_X1  g736(.A1(new_n1157), .A2(new_n1158), .B1(new_n1148), .B2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1153), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1146), .A2(new_n1163), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g739(.A1(new_n462), .A2(G227), .ZN(new_n1166));
  NAND2_X1  g740(.A1(new_n681), .A2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g741(.A1(new_n651), .A2(new_n1167), .ZN(new_n1168));
  AND3_X1   g742(.A1(new_n1168), .A2(new_n944), .A3(new_n864), .ZN(G308));
  NAND3_X1  g743(.A1(new_n1168), .A2(new_n944), .A3(new_n864), .ZN(G225));
endmodule


