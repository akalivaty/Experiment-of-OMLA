

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U551 ( .A1(n522), .A2(G2104), .ZN(n527) );
  NOR2_X2 U552 ( .A1(n973), .A2(n617), .ZN(n626) );
  NOR2_X2 U553 ( .A1(n638), .A2(n945), .ZN(n622) );
  NOR2_X1 U554 ( .A1(G164), .A2(G1384), .ZN(n709) );
  INV_X1 U555 ( .A(KEYINPUT17), .ZN(n518) );
  NOR2_X1 U556 ( .A1(G2105), .A2(G2104), .ZN(n519) );
  NOR2_X1 U557 ( .A1(n674), .A2(n648), .ZN(n650) );
  NAND2_X1 U558 ( .A1(n889), .A2(G137), .ZN(n531) );
  INV_X1 U559 ( .A(KEYINPUT23), .ZN(n528) );
  NOR2_X2 U560 ( .A1(n526), .A2(n525), .ZN(G164) );
  XOR2_X1 U561 ( .A(G543), .B(KEYINPUT0), .Z(n516) );
  INV_X1 U562 ( .A(G2105), .ZN(n522) );
  XNOR2_X1 U563 ( .A(n645), .B(KEYINPUT93), .ZN(n620) );
  INV_X1 U564 ( .A(KEYINPUT30), .ZN(n649) );
  BUF_X1 U565 ( .A(n645), .Z(n664) );
  XNOR2_X1 U566 ( .A(KEYINPUT29), .B(KEYINPUT100), .ZN(n635) );
  INV_X1 U567 ( .A(KEYINPUT92), .ZN(n646) );
  NOR2_X2 U568 ( .A1(n537), .A2(n575), .ZN(n799) );
  XNOR2_X1 U569 ( .A(KEYINPUT5), .B(KEYINPUT73), .ZN(n548) );
  NOR2_X2 U570 ( .A1(G651), .A2(n575), .ZN(n796) );
  XNOR2_X1 U571 ( .A(n549), .B(n548), .ZN(n554) );
  XNOR2_X1 U572 ( .A(n529), .B(n528), .ZN(n530) );
  NAND2_X1 U573 ( .A1(n527), .A2(G102), .ZN(n517) );
  XNOR2_X1 U574 ( .A(n517), .B(KEYINPUT88), .ZN(n521) );
  XNOR2_X2 U575 ( .A(n519), .B(n518), .ZN(n889) );
  NAND2_X1 U576 ( .A1(G138), .A2(n889), .ZN(n520) );
  NAND2_X1 U577 ( .A1(n521), .A2(n520), .ZN(n526) );
  NOR2_X2 U578 ( .A1(G2104), .A2(n522), .ZN(n885) );
  NAND2_X1 U579 ( .A1(G126), .A2(n885), .ZN(n524) );
  AND2_X1 U580 ( .A1(G2105), .A2(G2104), .ZN(n886) );
  NAND2_X1 U581 ( .A1(G114), .A2(n886), .ZN(n523) );
  NAND2_X1 U582 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U583 ( .A1(G101), .A2(n527), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n531), .A2(n530), .ZN(n535) );
  NAND2_X1 U585 ( .A1(G125), .A2(n885), .ZN(n533) );
  NAND2_X1 U586 ( .A1(G113), .A2(n886), .ZN(n532) );
  NAND2_X1 U587 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X2 U588 ( .A1(n535), .A2(n534), .ZN(G160) );
  INV_X1 U589 ( .A(G651), .ZN(n537) );
  NOR2_X1 U590 ( .A1(G543), .A2(n537), .ZN(n536) );
  XOR2_X1 U591 ( .A(KEYINPUT1), .B(n536), .Z(n795) );
  NAND2_X1 U592 ( .A1(G65), .A2(n795), .ZN(n539) );
  XNOR2_X1 U593 ( .A(KEYINPUT64), .B(n516), .ZN(n575) );
  NAND2_X1 U594 ( .A1(G78), .A2(n799), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n539), .A2(n538), .ZN(n543) );
  NOR2_X1 U596 ( .A1(G651), .A2(G543), .ZN(n800) );
  NAND2_X1 U597 ( .A1(G91), .A2(n800), .ZN(n541) );
  NAND2_X1 U598 ( .A1(G53), .A2(n796), .ZN(n540) );
  NAND2_X1 U599 ( .A1(n541), .A2(n540), .ZN(n542) );
  OR2_X1 U600 ( .A1(n543), .A2(n542), .ZN(G299) );
  XNOR2_X1 U601 ( .A(KEYINPUT7), .B(KEYINPUT74), .ZN(n556) );
  NAND2_X1 U602 ( .A1(n800), .A2(G89), .ZN(n544) );
  XOR2_X1 U603 ( .A(KEYINPUT4), .B(n544), .Z(n547) );
  NAND2_X1 U604 ( .A1(n799), .A2(G76), .ZN(n545) );
  XOR2_X1 U605 ( .A(KEYINPUT72), .B(n545), .Z(n546) );
  NOR2_X1 U606 ( .A1(n547), .A2(n546), .ZN(n549) );
  NAND2_X1 U607 ( .A1(G63), .A2(n795), .ZN(n551) );
  NAND2_X1 U608 ( .A1(G51), .A2(n796), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U610 ( .A(KEYINPUT6), .B(n552), .Z(n553) );
  NAND2_X1 U611 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U612 ( .A(n556), .B(n555), .ZN(G168) );
  NAND2_X1 U613 ( .A1(G64), .A2(n795), .ZN(n558) );
  NAND2_X1 U614 ( .A1(G52), .A2(n796), .ZN(n557) );
  NAND2_X1 U615 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U616 ( .A(KEYINPUT65), .B(n559), .Z(n564) );
  NAND2_X1 U617 ( .A1(G77), .A2(n799), .ZN(n561) );
  NAND2_X1 U618 ( .A1(G90), .A2(n800), .ZN(n560) );
  NAND2_X1 U619 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U620 ( .A(KEYINPUT9), .B(n562), .Z(n563) );
  NOR2_X1 U621 ( .A1(n564), .A2(n563), .ZN(G171) );
  XOR2_X1 U622 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U623 ( .A1(G75), .A2(n799), .ZN(n566) );
  NAND2_X1 U624 ( .A1(G88), .A2(n800), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U626 ( .A(KEYINPUT80), .B(n567), .ZN(n571) );
  NAND2_X1 U627 ( .A1(G62), .A2(n795), .ZN(n569) );
  NAND2_X1 U628 ( .A1(G50), .A2(n796), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U630 ( .A1(n571), .A2(n570), .ZN(G166) );
  XNOR2_X1 U631 ( .A(KEYINPUT89), .B(G166), .ZN(G303) );
  NAND2_X1 U632 ( .A1(G49), .A2(n796), .ZN(n573) );
  NAND2_X1 U633 ( .A1(G74), .A2(G651), .ZN(n572) );
  NAND2_X1 U634 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U635 ( .A1(n795), .A2(n574), .ZN(n578) );
  NAND2_X1 U636 ( .A1(n575), .A2(G87), .ZN(n576) );
  XOR2_X1 U637 ( .A(KEYINPUT79), .B(n576), .Z(n577) );
  NAND2_X1 U638 ( .A1(n578), .A2(n577), .ZN(G288) );
  NAND2_X1 U639 ( .A1(G61), .A2(n795), .ZN(n580) );
  NAND2_X1 U640 ( .A1(G86), .A2(n800), .ZN(n579) );
  NAND2_X1 U641 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U642 ( .A1(n799), .A2(G73), .ZN(n581) );
  XOR2_X1 U643 ( .A(KEYINPUT2), .B(n581), .Z(n582) );
  NOR2_X1 U644 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U645 ( .A1(n796), .A2(G48), .ZN(n584) );
  NAND2_X1 U646 ( .A1(n585), .A2(n584), .ZN(G305) );
  AND2_X1 U647 ( .A1(n795), .A2(G60), .ZN(n589) );
  NAND2_X1 U648 ( .A1(G72), .A2(n799), .ZN(n587) );
  NAND2_X1 U649 ( .A1(G85), .A2(n800), .ZN(n586) );
  NAND2_X1 U650 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U651 ( .A1(n589), .A2(n588), .ZN(n591) );
  NAND2_X1 U652 ( .A1(n796), .A2(G47), .ZN(n590) );
  NAND2_X1 U653 ( .A1(n591), .A2(n590), .ZN(G290) );
  NAND2_X1 U654 ( .A1(G160), .A2(G40), .ZN(n708) );
  INV_X1 U655 ( .A(n708), .ZN(n592) );
  NAND2_X1 U656 ( .A1(n592), .A2(n709), .ZN(n645) );
  NAND2_X1 U657 ( .A1(G2067), .A2(n620), .ZN(n594) );
  NAND2_X1 U658 ( .A1(G1348), .A2(n664), .ZN(n593) );
  NAND2_X1 U659 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U660 ( .A(n595), .B(KEYINPUT98), .ZN(n619) );
  NAND2_X1 U661 ( .A1(G92), .A2(n800), .ZN(n602) );
  NAND2_X1 U662 ( .A1(G66), .A2(n795), .ZN(n597) );
  NAND2_X1 U663 ( .A1(G79), .A2(n799), .ZN(n596) );
  NAND2_X1 U664 ( .A1(n597), .A2(n596), .ZN(n600) );
  NAND2_X1 U665 ( .A1(G54), .A2(n796), .ZN(n598) );
  XNOR2_X1 U666 ( .A(KEYINPUT71), .B(n598), .ZN(n599) );
  NOR2_X1 U667 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U668 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X2 U669 ( .A(n603), .B(KEYINPUT15), .ZN(n969) );
  NAND2_X1 U670 ( .A1(G56), .A2(n795), .ZN(n604) );
  XOR2_X1 U671 ( .A(KEYINPUT14), .B(n604), .Z(n611) );
  NAND2_X1 U672 ( .A1(n799), .A2(G68), .ZN(n605) );
  XNOR2_X1 U673 ( .A(KEYINPUT69), .B(n605), .ZN(n608) );
  NAND2_X1 U674 ( .A1(n800), .A2(G81), .ZN(n606) );
  XOR2_X1 U675 ( .A(KEYINPUT12), .B(n606), .Z(n607) );
  NOR2_X1 U676 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U677 ( .A(n609), .B(KEYINPUT13), .ZN(n610) );
  NOR2_X1 U678 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U679 ( .A1(n796), .A2(G43), .ZN(n612) );
  NAND2_X1 U680 ( .A1(n613), .A2(n612), .ZN(n973) );
  INV_X1 U681 ( .A(G1996), .ZN(n947) );
  NOR2_X1 U682 ( .A1(n664), .A2(n947), .ZN(n614) );
  XOR2_X1 U683 ( .A(n614), .B(KEYINPUT26), .Z(n616) );
  NAND2_X1 U684 ( .A1(n664), .A2(G1341), .ZN(n615) );
  NAND2_X1 U685 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U686 ( .A1(n969), .A2(n626), .ZN(n618) );
  NOR2_X1 U687 ( .A1(n619), .A2(n618), .ZN(n630) );
  INV_X1 U688 ( .A(n620), .ZN(n638) );
  INV_X1 U689 ( .A(G2072), .ZN(n945) );
  XOR2_X1 U690 ( .A(KEYINPUT97), .B(KEYINPUT27), .Z(n621) );
  XNOR2_X1 U691 ( .A(n622), .B(n621), .ZN(n624) );
  NAND2_X1 U692 ( .A1(n638), .A2(G1956), .ZN(n623) );
  NAND2_X1 U693 ( .A1(n624), .A2(n623), .ZN(n631) );
  NOR2_X2 U694 ( .A1(n631), .A2(G299), .ZN(n625) );
  XNOR2_X1 U695 ( .A(n625), .B(KEYINPUT99), .ZN(n628) );
  NAND2_X1 U696 ( .A1(n626), .A2(n969), .ZN(n627) );
  NAND2_X1 U697 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U698 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U699 ( .A1(G299), .A2(n631), .ZN(n632) );
  XOR2_X1 U700 ( .A(KEYINPUT28), .B(n632), .Z(n633) );
  NOR2_X1 U701 ( .A1(n634), .A2(n633), .ZN(n636) );
  XNOR2_X1 U702 ( .A(n636), .B(n635), .ZN(n644) );
  XOR2_X1 U703 ( .A(G2078), .B(KEYINPUT25), .Z(n637) );
  XNOR2_X1 U704 ( .A(KEYINPUT94), .B(n637), .ZN(n944) );
  NOR2_X1 U705 ( .A1(n638), .A2(n944), .ZN(n639) );
  XNOR2_X1 U706 ( .A(n639), .B(KEYINPUT95), .ZN(n641) );
  INV_X1 U707 ( .A(G1961), .ZN(n994) );
  NAND2_X1 U708 ( .A1(n994), .A2(n664), .ZN(n640) );
  NAND2_X1 U709 ( .A1(n641), .A2(n640), .ZN(n652) );
  NAND2_X1 U710 ( .A1(G171), .A2(n652), .ZN(n642) );
  XNOR2_X1 U711 ( .A(KEYINPUT96), .B(n642), .ZN(n643) );
  NAND2_X1 U712 ( .A1(n644), .A2(n643), .ZN(n662) );
  NOR2_X1 U713 ( .A1(G2084), .A2(n664), .ZN(n674) );
  NAND2_X1 U714 ( .A1(G8), .A2(n645), .ZN(n704) );
  NOR2_X1 U715 ( .A1(G1966), .A2(n704), .ZN(n647) );
  XNOR2_X1 U716 ( .A(n647), .B(n646), .ZN(n676) );
  NAND2_X1 U717 ( .A1(n676), .A2(G8), .ZN(n648) );
  XNOR2_X1 U718 ( .A(n650), .B(n649), .ZN(n651) );
  NOR2_X1 U719 ( .A1(n651), .A2(G168), .ZN(n654) );
  NOR2_X1 U720 ( .A1(G171), .A2(n652), .ZN(n653) );
  NOR2_X2 U721 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U722 ( .A1(KEYINPUT101), .A2(n655), .ZN(n659) );
  INV_X1 U723 ( .A(n655), .ZN(n657) );
  INV_X1 U724 ( .A(KEYINPUT101), .ZN(n656) );
  NAND2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U727 ( .A(n660), .B(KEYINPUT31), .ZN(n661) );
  NAND2_X1 U728 ( .A1(n662), .A2(n661), .ZN(n678) );
  AND2_X1 U729 ( .A1(G286), .A2(G8), .ZN(n663) );
  NAND2_X1 U730 ( .A1(n678), .A2(n663), .ZN(n671) );
  INV_X1 U731 ( .A(G8), .ZN(n669) );
  NOR2_X1 U732 ( .A1(G1971), .A2(n704), .ZN(n666) );
  NOR2_X1 U733 ( .A1(G2090), .A2(n664), .ZN(n665) );
  NOR2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U735 ( .A1(n667), .A2(G303), .ZN(n668) );
  OR2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n673) );
  INV_X1 U738 ( .A(KEYINPUT32), .ZN(n672) );
  XNOR2_X1 U739 ( .A(n673), .B(n672), .ZN(n694) );
  NAND2_X1 U740 ( .A1(G8), .A2(n674), .ZN(n675) );
  AND2_X1 U741 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U742 ( .A1(n678), .A2(n677), .ZN(n695) );
  NAND2_X1 U743 ( .A1(G1976), .A2(G288), .ZN(n978) );
  AND2_X1 U744 ( .A1(n695), .A2(n978), .ZN(n679) );
  NAND2_X1 U745 ( .A1(n694), .A2(n679), .ZN(n684) );
  INV_X1 U746 ( .A(n978), .ZN(n682) );
  NOR2_X1 U747 ( .A1(G1976), .A2(G288), .ZN(n976) );
  NOR2_X1 U748 ( .A1(G1971), .A2(G303), .ZN(n680) );
  NOR2_X1 U749 ( .A1(n976), .A2(n680), .ZN(n681) );
  OR2_X1 U750 ( .A1(n682), .A2(n681), .ZN(n683) );
  AND2_X1 U751 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U752 ( .A1(n685), .A2(n704), .ZN(n686) );
  NOR2_X1 U753 ( .A1(KEYINPUT33), .A2(n686), .ZN(n688) );
  INV_X1 U754 ( .A(KEYINPUT102), .ZN(n687) );
  XNOR2_X1 U755 ( .A(n688), .B(n687), .ZN(n692) );
  NAND2_X1 U756 ( .A1(n976), .A2(KEYINPUT33), .ZN(n689) );
  OR2_X1 U757 ( .A1(n704), .A2(n689), .ZN(n690) );
  XOR2_X1 U758 ( .A(G1981), .B(G305), .Z(n985) );
  AND2_X1 U759 ( .A1(n690), .A2(n985), .ZN(n691) );
  NAND2_X1 U760 ( .A1(n692), .A2(n691), .ZN(n700) );
  NOR2_X1 U761 ( .A1(G2090), .A2(G303), .ZN(n693) );
  NAND2_X1 U762 ( .A1(G8), .A2(n693), .ZN(n697) );
  NAND2_X1 U763 ( .A1(n694), .A2(n695), .ZN(n696) );
  NAND2_X1 U764 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U765 ( .A1(n698), .A2(n704), .ZN(n699) );
  NAND2_X1 U766 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U767 ( .A(n701), .B(KEYINPUT103), .ZN(n707) );
  NOR2_X1 U768 ( .A1(G1981), .A2(G305), .ZN(n702) );
  XNOR2_X1 U769 ( .A(n702), .B(KEYINPUT91), .ZN(n703) );
  XNOR2_X1 U770 ( .A(n703), .B(KEYINPUT24), .ZN(n705) );
  OR2_X1 U771 ( .A1(n705), .A2(n704), .ZN(n706) );
  AND2_X1 U772 ( .A1(n707), .A2(n706), .ZN(n727) );
  NOR2_X1 U773 ( .A1(n709), .A2(n708), .ZN(n752) );
  NAND2_X1 U774 ( .A1(G129), .A2(n885), .ZN(n711) );
  NAND2_X1 U775 ( .A1(G141), .A2(n889), .ZN(n710) );
  NAND2_X1 U776 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U777 ( .A1(n527), .A2(G105), .ZN(n712) );
  XOR2_X1 U778 ( .A(KEYINPUT38), .B(n712), .Z(n713) );
  NOR2_X1 U779 ( .A1(n714), .A2(n713), .ZN(n716) );
  NAND2_X1 U780 ( .A1(n886), .A2(G117), .ZN(n715) );
  NAND2_X1 U781 ( .A1(n716), .A2(n715), .ZN(n884) );
  NAND2_X1 U782 ( .A1(G1996), .A2(n884), .ZN(n724) );
  NAND2_X1 U783 ( .A1(G119), .A2(n885), .ZN(n718) );
  NAND2_X1 U784 ( .A1(G131), .A2(n889), .ZN(n717) );
  NAND2_X1 U785 ( .A1(n718), .A2(n717), .ZN(n722) );
  NAND2_X1 U786 ( .A1(G95), .A2(n527), .ZN(n720) );
  NAND2_X1 U787 ( .A1(G107), .A2(n886), .ZN(n719) );
  NAND2_X1 U788 ( .A1(n720), .A2(n719), .ZN(n721) );
  OR2_X1 U789 ( .A1(n722), .A2(n721), .ZN(n872) );
  NAND2_X1 U790 ( .A1(G1991), .A2(n872), .ZN(n723) );
  NAND2_X1 U791 ( .A1(n724), .A2(n723), .ZN(n928) );
  NAND2_X1 U792 ( .A1(n752), .A2(n928), .ZN(n740) );
  XNOR2_X1 U793 ( .A(G1986), .B(G290), .ZN(n968) );
  NAND2_X1 U794 ( .A1(n752), .A2(n968), .ZN(n725) );
  NAND2_X1 U795 ( .A1(n740), .A2(n725), .ZN(n726) );
  NOR2_X1 U796 ( .A1(n727), .A2(n726), .ZN(n738) );
  XNOR2_X1 U797 ( .A(G2067), .B(KEYINPUT37), .ZN(n749) );
  NAND2_X1 U798 ( .A1(G104), .A2(n527), .ZN(n729) );
  NAND2_X1 U799 ( .A1(G140), .A2(n889), .ZN(n728) );
  NAND2_X1 U800 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U801 ( .A(KEYINPUT34), .B(n730), .ZN(n736) );
  NAND2_X1 U802 ( .A1(n886), .A2(G116), .ZN(n731) );
  XNOR2_X1 U803 ( .A(n731), .B(KEYINPUT90), .ZN(n733) );
  NAND2_X1 U804 ( .A1(G128), .A2(n885), .ZN(n732) );
  NAND2_X1 U805 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U806 ( .A(KEYINPUT35), .B(n734), .Z(n735) );
  NOR2_X1 U807 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U808 ( .A(KEYINPUT36), .B(n737), .ZN(n901) );
  NOR2_X1 U809 ( .A1(n749), .A2(n901), .ZN(n932) );
  NAND2_X1 U810 ( .A1(n752), .A2(n932), .ZN(n747) );
  NAND2_X1 U811 ( .A1(n738), .A2(n747), .ZN(n739) );
  XNOR2_X1 U812 ( .A(n739), .B(KEYINPUT104), .ZN(n754) );
  NOR2_X1 U813 ( .A1(G1996), .A2(n884), .ZN(n920) );
  INV_X1 U814 ( .A(n740), .ZN(n743) );
  NOR2_X1 U815 ( .A1(G1991), .A2(n872), .ZN(n926) );
  NOR2_X1 U816 ( .A1(G1986), .A2(G290), .ZN(n741) );
  NOR2_X1 U817 ( .A1(n926), .A2(n741), .ZN(n742) );
  NOR2_X1 U818 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U819 ( .A(KEYINPUT105), .B(n744), .Z(n745) );
  NOR2_X1 U820 ( .A1(n920), .A2(n745), .ZN(n746) );
  XNOR2_X1 U821 ( .A(n746), .B(KEYINPUT39), .ZN(n748) );
  NAND2_X1 U822 ( .A1(n748), .A2(n747), .ZN(n750) );
  NAND2_X1 U823 ( .A1(n749), .A2(n901), .ZN(n923) );
  NAND2_X1 U824 ( .A1(n750), .A2(n923), .ZN(n751) );
  NAND2_X1 U825 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U826 ( .A1(n754), .A2(n753), .ZN(n756) );
  XNOR2_X1 U827 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n755) );
  XNOR2_X1 U828 ( .A(n756), .B(n755), .ZN(G329) );
  XOR2_X1 U829 ( .A(G2443), .B(G2446), .Z(n758) );
  XNOR2_X1 U830 ( .A(G2427), .B(G2451), .ZN(n757) );
  XNOR2_X1 U831 ( .A(n758), .B(n757), .ZN(n764) );
  XOR2_X1 U832 ( .A(G2430), .B(G2454), .Z(n760) );
  XNOR2_X1 U833 ( .A(G1341), .B(G1348), .ZN(n759) );
  XNOR2_X1 U834 ( .A(n760), .B(n759), .ZN(n762) );
  XOR2_X1 U835 ( .A(G2435), .B(G2438), .Z(n761) );
  XNOR2_X1 U836 ( .A(n762), .B(n761), .ZN(n763) );
  XOR2_X1 U837 ( .A(n764), .B(n763), .Z(n765) );
  AND2_X1 U838 ( .A1(G14), .A2(n765), .ZN(G401) );
  AND2_X1 U839 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U840 ( .A(G120), .ZN(G236) );
  INV_X1 U841 ( .A(G69), .ZN(G235) );
  INV_X1 U842 ( .A(G57), .ZN(G237) );
  INV_X1 U843 ( .A(G132), .ZN(G219) );
  INV_X1 U844 ( .A(G82), .ZN(G220) );
  XOR2_X1 U845 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n767) );
  NAND2_X1 U846 ( .A1(G7), .A2(G661), .ZN(n766) );
  XNOR2_X1 U847 ( .A(n767), .B(n766), .ZN(n768) );
  XNOR2_X1 U848 ( .A(KEYINPUT66), .B(n768), .ZN(G223) );
  XOR2_X1 U849 ( .A(KEYINPUT11), .B(KEYINPUT68), .Z(n770) );
  INV_X1 U850 ( .A(G223), .ZN(n836) );
  NAND2_X1 U851 ( .A1(n836), .A2(G567), .ZN(n769) );
  XNOR2_X1 U852 ( .A(n770), .B(n769), .ZN(G234) );
  INV_X1 U853 ( .A(G860), .ZN(n794) );
  OR2_X1 U854 ( .A1(n973), .A2(n794), .ZN(G153) );
  XOR2_X1 U855 ( .A(G171), .B(KEYINPUT70), .Z(G301) );
  NAND2_X1 U856 ( .A1(G868), .A2(G301), .ZN(n772) );
  OR2_X1 U857 ( .A1(n969), .A2(G868), .ZN(n771) );
  NAND2_X1 U858 ( .A1(n772), .A2(n771), .ZN(G284) );
  INV_X1 U859 ( .A(G868), .ZN(n773) );
  NAND2_X1 U860 ( .A1(G299), .A2(n773), .ZN(n775) );
  NAND2_X1 U861 ( .A1(G868), .A2(G286), .ZN(n774) );
  NAND2_X1 U862 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U863 ( .A(KEYINPUT75), .B(n776), .Z(G297) );
  NAND2_X1 U864 ( .A1(n794), .A2(G559), .ZN(n777) );
  NAND2_X1 U865 ( .A1(n777), .A2(n969), .ZN(n778) );
  XNOR2_X1 U866 ( .A(n778), .B(KEYINPUT76), .ZN(n779) );
  XNOR2_X1 U867 ( .A(KEYINPUT16), .B(n779), .ZN(G148) );
  NOR2_X1 U868 ( .A1(G868), .A2(n973), .ZN(n782) );
  NAND2_X1 U869 ( .A1(G868), .A2(n969), .ZN(n780) );
  NOR2_X1 U870 ( .A1(G559), .A2(n780), .ZN(n781) );
  NOR2_X1 U871 ( .A1(n782), .A2(n781), .ZN(G282) );
  NAND2_X1 U872 ( .A1(G123), .A2(n885), .ZN(n783) );
  XNOR2_X1 U873 ( .A(n783), .B(KEYINPUT18), .ZN(n786) );
  NAND2_X1 U874 ( .A1(G135), .A2(n889), .ZN(n784) );
  XOR2_X1 U875 ( .A(KEYINPUT77), .B(n784), .Z(n785) );
  NAND2_X1 U876 ( .A1(n786), .A2(n785), .ZN(n790) );
  NAND2_X1 U877 ( .A1(G99), .A2(n527), .ZN(n788) );
  NAND2_X1 U878 ( .A1(G111), .A2(n886), .ZN(n787) );
  NAND2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U880 ( .A1(n790), .A2(n789), .ZN(n925) );
  XOR2_X1 U881 ( .A(G2096), .B(n925), .Z(n791) );
  NOR2_X1 U882 ( .A1(G2100), .A2(n791), .ZN(n792) );
  XOR2_X1 U883 ( .A(KEYINPUT78), .B(n792), .Z(G156) );
  NAND2_X1 U884 ( .A1(G559), .A2(n969), .ZN(n793) );
  XOR2_X1 U885 ( .A(n973), .B(n793), .Z(n814) );
  NAND2_X1 U886 ( .A1(n794), .A2(n814), .ZN(n805) );
  NAND2_X1 U887 ( .A1(G67), .A2(n795), .ZN(n798) );
  NAND2_X1 U888 ( .A1(G55), .A2(n796), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n804) );
  NAND2_X1 U890 ( .A1(G80), .A2(n799), .ZN(n802) );
  NAND2_X1 U891 ( .A1(G93), .A2(n800), .ZN(n801) );
  NAND2_X1 U892 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U893 ( .A1(n804), .A2(n803), .ZN(n809) );
  XOR2_X1 U894 ( .A(n805), .B(n809), .Z(G145) );
  OR2_X1 U895 ( .A1(G868), .A2(n809), .ZN(n806) );
  XNOR2_X1 U896 ( .A(n806), .B(KEYINPUT82), .ZN(n817) );
  XOR2_X1 U897 ( .A(KEYINPUT19), .B(KEYINPUT81), .Z(n807) );
  XNOR2_X1 U898 ( .A(G290), .B(n807), .ZN(n808) );
  XNOR2_X1 U899 ( .A(n809), .B(n808), .ZN(n811) );
  XNOR2_X1 U900 ( .A(G305), .B(G166), .ZN(n810) );
  XNOR2_X1 U901 ( .A(n811), .B(n810), .ZN(n812) );
  XNOR2_X1 U902 ( .A(n812), .B(G299), .ZN(n813) );
  XNOR2_X1 U903 ( .A(n813), .B(G288), .ZN(n905) );
  XNOR2_X1 U904 ( .A(n905), .B(n814), .ZN(n815) );
  NAND2_X1 U905 ( .A1(G868), .A2(n815), .ZN(n816) );
  NAND2_X1 U906 ( .A1(n817), .A2(n816), .ZN(G295) );
  NAND2_X1 U907 ( .A1(G2078), .A2(G2084), .ZN(n818) );
  XNOR2_X1 U908 ( .A(n818), .B(KEYINPUT20), .ZN(n819) );
  XNOR2_X1 U909 ( .A(n819), .B(KEYINPUT83), .ZN(n820) );
  NAND2_X1 U910 ( .A1(n820), .A2(G2090), .ZN(n821) );
  XNOR2_X1 U911 ( .A(KEYINPUT21), .B(n821), .ZN(n822) );
  NAND2_X1 U912 ( .A1(n822), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U913 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U914 ( .A1(G220), .A2(G219), .ZN(n823) );
  XOR2_X1 U915 ( .A(KEYINPUT22), .B(n823), .Z(n824) );
  NOR2_X1 U916 ( .A1(G218), .A2(n824), .ZN(n825) );
  XNOR2_X1 U917 ( .A(KEYINPUT84), .B(n825), .ZN(n826) );
  NAND2_X1 U918 ( .A1(n826), .A2(G96), .ZN(n841) );
  NAND2_X1 U919 ( .A1(n841), .A2(G2106), .ZN(n832) );
  NOR2_X1 U920 ( .A1(G235), .A2(G236), .ZN(n827) );
  XNOR2_X1 U921 ( .A(n827), .B(KEYINPUT85), .ZN(n828) );
  NOR2_X1 U922 ( .A1(G237), .A2(n828), .ZN(n829) );
  XNOR2_X1 U923 ( .A(KEYINPUT86), .B(n829), .ZN(n830) );
  NAND2_X1 U924 ( .A1(n830), .A2(G108), .ZN(n840) );
  NAND2_X1 U925 ( .A1(G567), .A2(n840), .ZN(n831) );
  NAND2_X1 U926 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U927 ( .A(n833), .B(KEYINPUT87), .ZN(G319) );
  INV_X1 U928 ( .A(G319), .ZN(n835) );
  NAND2_X1 U929 ( .A1(G661), .A2(G483), .ZN(n834) );
  NOR2_X1 U930 ( .A1(n835), .A2(n834), .ZN(n839) );
  NAND2_X1 U931 ( .A1(n839), .A2(G36), .ZN(G176) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n836), .ZN(G217) );
  AND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U934 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U936 ( .A1(n839), .A2(n838), .ZN(G188) );
  INV_X1 U938 ( .A(G108), .ZN(G238) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  NOR2_X1 U940 ( .A1(n841), .A2(n840), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  XOR2_X1 U942 ( .A(G2096), .B(G2072), .Z(n843) );
  XNOR2_X1 U943 ( .A(G2067), .B(G2090), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n853) );
  XOR2_X1 U945 ( .A(KEYINPUT110), .B(G2678), .Z(n845) );
  XNOR2_X1 U946 ( .A(KEYINPUT109), .B(KEYINPUT107), .ZN(n844) );
  XNOR2_X1 U947 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U948 ( .A(G2100), .B(KEYINPUT43), .Z(n847) );
  XNOR2_X1 U949 ( .A(KEYINPUT42), .B(KEYINPUT108), .ZN(n846) );
  XNOR2_X1 U950 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U951 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U952 ( .A(G2078), .B(G2084), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U954 ( .A(n853), .B(n852), .Z(G227) );
  XOR2_X1 U955 ( .A(G1976), .B(G1971), .Z(n855) );
  XNOR2_X1 U956 ( .A(G1966), .B(G1956), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U958 ( .A(G1981), .B(G1986), .Z(n857) );
  XNOR2_X1 U959 ( .A(G1996), .B(G1991), .ZN(n856) );
  XNOR2_X1 U960 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U961 ( .A(n859), .B(n858), .Z(n861) );
  XNOR2_X1 U962 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n860) );
  XNOR2_X1 U963 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U964 ( .A(G2474), .B(n862), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n863), .B(n994), .ZN(G229) );
  NAND2_X1 U966 ( .A1(G100), .A2(n527), .ZN(n865) );
  NAND2_X1 U967 ( .A1(G112), .A2(n886), .ZN(n864) );
  NAND2_X1 U968 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U969 ( .A(KEYINPUT112), .B(n866), .ZN(n871) );
  NAND2_X1 U970 ( .A1(n885), .A2(G124), .ZN(n867) );
  XNOR2_X1 U971 ( .A(n867), .B(KEYINPUT44), .ZN(n869) );
  NAND2_X1 U972 ( .A1(G136), .A2(n889), .ZN(n868) );
  NAND2_X1 U973 ( .A1(n869), .A2(n868), .ZN(n870) );
  NOR2_X1 U974 ( .A1(n871), .A2(n870), .ZN(G162) );
  XNOR2_X1 U975 ( .A(KEYINPUT48), .B(KEYINPUT114), .ZN(n874) );
  XNOR2_X1 U976 ( .A(n872), .B(KEYINPUT46), .ZN(n873) );
  XNOR2_X1 U977 ( .A(n874), .B(n873), .ZN(n900) );
  NAND2_X1 U978 ( .A1(G103), .A2(n527), .ZN(n876) );
  NAND2_X1 U979 ( .A1(G139), .A2(n889), .ZN(n875) );
  NAND2_X1 U980 ( .A1(n876), .A2(n875), .ZN(n882) );
  NAND2_X1 U981 ( .A1(n885), .A2(G127), .ZN(n877) );
  XOR2_X1 U982 ( .A(KEYINPUT113), .B(n877), .Z(n879) );
  NAND2_X1 U983 ( .A1(n886), .A2(G115), .ZN(n878) );
  NAND2_X1 U984 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U985 ( .A(KEYINPUT47), .B(n880), .Z(n881) );
  NOR2_X1 U986 ( .A1(n882), .A2(n881), .ZN(n915) );
  XOR2_X1 U987 ( .A(n915), .B(G162), .Z(n883) );
  XNOR2_X1 U988 ( .A(n884), .B(n883), .ZN(n896) );
  NAND2_X1 U989 ( .A1(G130), .A2(n885), .ZN(n888) );
  NAND2_X1 U990 ( .A1(G118), .A2(n886), .ZN(n887) );
  NAND2_X1 U991 ( .A1(n888), .A2(n887), .ZN(n894) );
  NAND2_X1 U992 ( .A1(G106), .A2(n527), .ZN(n891) );
  NAND2_X1 U993 ( .A1(G142), .A2(n889), .ZN(n890) );
  NAND2_X1 U994 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U995 ( .A(KEYINPUT45), .B(n892), .Z(n893) );
  NOR2_X1 U996 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U997 ( .A(n896), .B(n895), .Z(n898) );
  XNOR2_X1 U998 ( .A(G164), .B(G160), .ZN(n897) );
  XNOR2_X1 U999 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U1000 ( .A(n900), .B(n899), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(n901), .B(n925), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n904), .ZN(G395) );
  XNOR2_X1 U1004 ( .A(G286), .B(n905), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n969), .B(G171), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(n908), .B(n973), .ZN(n909) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n909), .ZN(G397) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1011 ( .A1(G401), .A2(n911), .ZN(n912) );
  AND2_X1 U1012 ( .A1(G319), .A2(n912), .ZN(n914) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1016 ( .A(G164), .B(G2078), .Z(n917) );
  XNOR2_X1 U1017 ( .A(n945), .B(n915), .ZN(n916) );
  NOR2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1019 ( .A(KEYINPUT50), .B(n918), .Z(n938) );
  XOR2_X1 U1020 ( .A(G2090), .B(G162), .Z(n919) );
  NOR2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1022 ( .A(KEYINPUT51), .B(n921), .Z(n922) );
  XNOR2_X1 U1023 ( .A(n922), .B(KEYINPUT116), .ZN(n924) );
  NAND2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n935) );
  NOR2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n930) );
  XOR2_X1 U1026 ( .A(G160), .B(G2084), .Z(n927) );
  NOR2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(n933), .B(KEYINPUT115), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(KEYINPUT117), .B(n936), .ZN(n937) );
  NOR2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1034 ( .A(KEYINPUT52), .B(n939), .ZN(n941) );
  INV_X1 U1035 ( .A(KEYINPUT55), .ZN(n940) );
  NAND2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1037 ( .A1(n942), .A2(G29), .ZN(n1028) );
  XOR2_X1 U1038 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n943) );
  XNOR2_X1 U1039 ( .A(KEYINPUT120), .B(n943), .ZN(n958) );
  XNOR2_X1 U1040 ( .A(G27), .B(n944), .ZN(n956) );
  XNOR2_X1 U1041 ( .A(G33), .B(n945), .ZN(n946) );
  NAND2_X1 U1042 ( .A1(n946), .A2(G28), .ZN(n950) );
  XOR2_X1 U1043 ( .A(G32), .B(n947), .Z(n948) );
  XNOR2_X1 U1044 ( .A(KEYINPUT118), .B(n948), .ZN(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(G2067), .B(G26), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(G25), .B(G1991), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(n958), .B(n957), .ZN(n964) );
  XOR2_X1 U1052 ( .A(G2090), .B(G35), .Z(n962) );
  XNOR2_X1 U1053 ( .A(KEYINPUT54), .B(G34), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(n959), .B(KEYINPUT121), .ZN(n960) );
  XNOR2_X1 U1055 ( .A(n960), .B(G2084), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n1020) );
  NAND2_X1 U1058 ( .A1(KEYINPUT55), .A2(n1020), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(G11), .A2(n965), .ZN(n1026) );
  INV_X1 U1060 ( .A(G16), .ZN(n1016) );
  XOR2_X1 U1061 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n966) );
  XNOR2_X1 U1062 ( .A(n1016), .B(n966), .ZN(n993) );
  XOR2_X1 U1063 ( .A(G171), .B(G1961), .Z(n967) );
  NOR2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n972) );
  XOR2_X1 U1065 ( .A(n969), .B(G1348), .Z(n970) );
  XNOR2_X1 U1066 ( .A(KEYINPUT123), .B(n970), .ZN(n971) );
  NAND2_X1 U1067 ( .A1(n972), .A2(n971), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(G1341), .B(n973), .ZN(n974) );
  NOR2_X1 U1069 ( .A1(n975), .A2(n974), .ZN(n991) );
  INV_X1 U1070 ( .A(n976), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  XOR2_X1 U1072 ( .A(KEYINPUT124), .B(n979), .Z(n983) );
  XNOR2_X1 U1073 ( .A(G1971), .B(G303), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(G1956), .B(G299), .ZN(n980) );
  NOR2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1077 ( .A(KEYINPUT125), .B(n984), .Z(n989) );
  XNOR2_X1 U1078 ( .A(G1966), .B(G168), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1080 ( .A(KEYINPUT57), .B(n987), .Z(n988) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n1018) );
  XNOR2_X1 U1084 ( .A(G5), .B(n994), .ZN(n1011) );
  XOR2_X1 U1085 ( .A(G1348), .B(KEYINPUT59), .Z(n995) );
  XNOR2_X1 U1086 ( .A(G4), .B(n995), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(G20), .B(G1956), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(G1981), .B(G6), .ZN(n999) );
  XNOR2_X1 U1090 ( .A(G19), .B(G1341), .ZN(n998) );
  NOR2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(n1002), .B(KEYINPUT60), .ZN(n1009) );
  XNOR2_X1 U1094 ( .A(G1971), .B(G22), .ZN(n1004) );
  XNOR2_X1 U1095 ( .A(G23), .B(G1976), .ZN(n1003) );
  NOR2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XOR2_X1 U1097 ( .A(G1986), .B(G24), .Z(n1005) );
  NAND2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1099 ( .A(KEYINPUT58), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(G21), .B(G1966), .ZN(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XNOR2_X1 U1104 ( .A(KEYINPUT61), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1107 ( .A(KEYINPUT126), .B(n1019), .Z(n1024) );
  INV_X1 U1108 ( .A(n1020), .ZN(n1022) );
  NOR2_X1 U1109 ( .A1(G29), .A2(KEYINPUT55), .ZN(n1021) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1113 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1114 ( .A(n1029), .B(KEYINPUT62), .ZN(n1030) );
  XNOR2_X1 U1115 ( .A(KEYINPUT127), .B(n1030), .ZN(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

