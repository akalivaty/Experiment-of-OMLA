

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737;

  AND2_X1 U372 ( .A1(n363), .A2(n609), .ZN(n679) );
  BUF_X1 U373 ( .A(n586), .Z(n596) );
  XNOR2_X2 U374 ( .A(KEYINPUT93), .B(n596), .ZN(n598) );
  XNOR2_X2 U375 ( .A(n572), .B(KEYINPUT32), .ZN(n734) );
  XOR2_X2 U376 ( .A(KEYINPUT4), .B(G101), .Z(n506) );
  XNOR2_X2 U377 ( .A(n441), .B(n400), .ZN(n455) );
  XNOR2_X2 U378 ( .A(n401), .B(G128), .ZN(n441) );
  XNOR2_X2 U379 ( .A(G140), .B(KEYINPUT69), .ZN(n478) );
  AND2_X1 U380 ( .A1(n396), .A2(n394), .ZN(n609) );
  AND2_X1 U381 ( .A1(n594), .A2(n582), .ZN(n585) );
  NOR2_X1 U382 ( .A1(n570), .A2(n523), .ZN(n503) );
  INV_X1 U383 ( .A(KEYINPUT16), .ZN(n424) );
  NOR2_X2 U384 ( .A1(n610), .A2(n679), .ZN(n693) );
  NOR2_X1 U385 ( .A1(n575), .A2(n574), .ZN(n576) );
  AND2_X1 U386 ( .A1(n669), .A2(KEYINPUT34), .ZN(n382) );
  XOR2_X1 U387 ( .A(n476), .B(KEYINPUT106), .Z(n631) );
  NAND2_X1 U388 ( .A1(n415), .A2(n413), .ZN(n567) );
  NAND2_X1 U389 ( .A1(n414), .A2(n351), .ZN(n413) );
  AND2_X1 U390 ( .A1(n417), .A2(n416), .ZN(n415) );
  BUF_X1 U391 ( .A(n532), .Z(n547) );
  NOR2_X1 U392 ( .A1(G902), .A2(n690), .ZN(n448) );
  NAND2_X1 U393 ( .A1(n656), .A2(KEYINPUT19), .ZN(n416) );
  XNOR2_X1 U394 ( .A(KEYINPUT87), .B(n436), .ZN(n608) );
  XNOR2_X1 U395 ( .A(n467), .B(n424), .ZN(n423) );
  BUF_X1 U396 ( .A(n693), .Z(n699) );
  XNOR2_X1 U397 ( .A(n581), .B(KEYINPUT75), .ZN(n594) );
  XOR2_X1 U398 ( .A(G146), .B(G125), .Z(n462) );
  XNOR2_X1 U399 ( .A(n462), .B(n369), .ZN(n479) );
  XNOR2_X1 U400 ( .A(KEYINPUT10), .B(KEYINPUT67), .ZN(n369) );
  INV_X1 U401 ( .A(G143), .ZN(n401) );
  XNOR2_X1 U402 ( .A(n430), .B(n429), .ZN(n445) );
  XOR2_X1 U403 ( .A(n704), .B(KEYINPUT72), .Z(n430) );
  AND2_X1 U404 ( .A1(n551), .A2(n552), .ZN(n657) );
  XNOR2_X1 U405 ( .A(n426), .B(n425), .ZN(n428) );
  NOR2_X1 U406 ( .A1(KEYINPUT47), .A2(n542), .ZN(n543) );
  INV_X1 U407 ( .A(n410), .ZN(n406) );
  XNOR2_X1 U408 ( .A(n465), .B(n354), .ZN(n466) );
  INV_X1 U409 ( .A(KEYINPUT17), .ZN(n433) );
  XNOR2_X1 U410 ( .A(n432), .B(n431), .ZN(n422) );
  NOR2_X1 U411 ( .A1(n733), .A2(n395), .ZN(n394) );
  INV_X1 U412 ( .A(n638), .ZN(n395) );
  XOR2_X1 U413 ( .A(n475), .B(n474), .Z(n551) );
  NOR2_X1 U414 ( .A1(G902), .A2(n611), .ZN(n475) );
  XOR2_X1 U415 ( .A(G122), .B(G104), .Z(n467) );
  XNOR2_X1 U416 ( .A(KEYINPUT96), .B(KEYINPUT23), .ZN(n482) );
  XNOR2_X1 U417 ( .A(G119), .B(G128), .ZN(n480) );
  INV_X1 U418 ( .A(G134), .ZN(n400) );
  XNOR2_X1 U419 ( .A(G107), .B(KEYINPUT100), .ZN(n374) );
  XNOR2_X1 U420 ( .A(n512), .B(n392), .ZN(n690) );
  XNOR2_X1 U421 ( .A(n393), .B(n445), .ZN(n392) );
  XNOR2_X1 U422 ( .A(n583), .B(KEYINPUT85), .ZN(n584) );
  NOR2_X1 U423 ( .A1(n516), .A2(n515), .ZN(n537) );
  NOR2_X1 U424 ( .A1(n669), .A2(KEYINPUT34), .ZN(n385) );
  XNOR2_X1 U425 ( .A(n492), .B(n355), .ZN(n577) );
  XNOR2_X1 U426 ( .A(n461), .B(G478), .ZN(n552) );
  XNOR2_X1 U427 ( .A(n366), .B(n512), .ZN(n616) );
  XNOR2_X1 U428 ( .A(n511), .B(n513), .ZN(n366) );
  NAND2_X1 U429 ( .A1(n388), .A2(n387), .ZN(n391) );
  NOR2_X1 U430 ( .A1(n679), .A2(n412), .ZN(n388) );
  INV_X1 U431 ( .A(n610), .ZN(n387) );
  AND2_X1 U432 ( .A1(n561), .A2(n631), .ZN(n550) );
  INV_X1 U433 ( .A(KEYINPUT44), .ZN(n378) );
  NOR2_X1 U434 ( .A1(n558), .A2(n559), .ZN(n397) );
  XOR2_X1 U435 ( .A(G902), .B(KEYINPUT15), .Z(n436) );
  NAND2_X1 U436 ( .A1(G234), .A2(G237), .ZN(n495) );
  XOR2_X1 U437 ( .A(KEYINPUT14), .B(KEYINPUT91), .Z(n496) );
  OR2_X1 U438 ( .A1(G237), .A2(G902), .ZN(n439) );
  NOR2_X1 U439 ( .A1(n656), .A2(n655), .ZN(n659) );
  XOR2_X1 U440 ( .A(KEYINPUT38), .B(n547), .Z(n655) );
  INV_X1 U441 ( .A(n403), .ZN(n407) );
  NOR2_X1 U442 ( .A1(n656), .A2(n406), .ZN(n405) );
  NAND2_X1 U443 ( .A1(n412), .A2(G902), .ZN(n410) );
  NAND2_X1 U444 ( .A1(n616), .A2(n412), .ZN(n411) );
  OR2_X1 U445 ( .A1(n616), .A2(n408), .ZN(n403) );
  NAND2_X1 U446 ( .A1(G472), .A2(n409), .ZN(n408) );
  INV_X1 U447 ( .A(G902), .ZN(n409) );
  NOR2_X1 U448 ( .A1(n577), .A2(n570), .ZN(n643) );
  XNOR2_X1 U449 ( .A(n514), .B(n649), .ZN(n582) );
  NOR2_X1 U450 ( .A1(G953), .A2(G237), .ZN(n508) );
  XNOR2_X1 U451 ( .A(G953), .B(KEYINPUT64), .ZN(n499) );
  INV_X1 U452 ( .A(n609), .ZN(n726) );
  XNOR2_X1 U453 ( .A(n472), .B(n370), .ZN(n611) );
  XNOR2_X1 U454 ( .A(n473), .B(n471), .ZN(n370) );
  XNOR2_X1 U455 ( .A(n421), .B(n420), .ZN(n685) );
  XNOR2_X1 U456 ( .A(n706), .B(n422), .ZN(n421) );
  XNOR2_X1 U457 ( .A(n434), .B(n433), .ZN(n435) );
  AND2_X1 U458 ( .A1(n710), .A2(KEYINPUT2), .ZN(n363) );
  XNOR2_X1 U459 ( .A(n399), .B(n398), .ZN(n561) );
  INV_X1 U460 ( .A(KEYINPUT39), .ZN(n398) );
  NOR2_X1 U461 ( .A1(n548), .A2(n655), .ZN(n399) );
  NAND2_X1 U462 ( .A1(n403), .A2(n402), .ZN(n573) );
  AND2_X1 U463 ( .A1(n411), .A2(n410), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n361), .B(KEYINPUT22), .ZN(n575) );
  AND2_X1 U465 ( .A1(n657), .A2(n639), .ZN(n365) );
  INV_X1 U466 ( .A(n573), .ZN(n649) );
  XNOR2_X1 U467 ( .A(n719), .B(n486), .ZN(n487) );
  XNOR2_X1 U468 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U469 ( .A(n459), .B(n373), .ZN(n697) );
  XNOR2_X1 U470 ( .A(n458), .B(n460), .ZN(n373) );
  XNOR2_X1 U471 ( .A(n455), .B(n374), .ZN(n456) );
  INV_X1 U472 ( .A(G953), .ZN(n709) );
  NAND2_X1 U473 ( .A1(n385), .A2(n386), .ZN(n383) );
  NOR2_X1 U474 ( .A1(n534), .A2(n552), .ZN(n633) );
  NAND2_X1 U475 ( .A1(n552), .A2(n534), .ZN(n476) );
  XNOR2_X1 U476 ( .A(n362), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U477 ( .A1(n390), .A2(n389), .ZN(n362) );
  XNOR2_X1 U478 ( .A(n391), .B(n353), .ZN(n390) );
  XNOR2_X1 U479 ( .A(n694), .B(n695), .ZN(n372) );
  NOR2_X1 U480 ( .A1(n656), .A2(KEYINPUT19), .ZN(n351) );
  AND2_X1 U481 ( .A1(n372), .A2(n389), .ZN(G54) );
  XOR2_X1 U482 ( .A(n616), .B(n359), .Z(n353) );
  AND2_X1 U483 ( .A1(G214), .A2(n508), .ZN(n354) );
  XOR2_X1 U484 ( .A(n491), .B(n490), .Z(n355) );
  XOR2_X1 U485 ( .A(KEYINPUT45), .B(KEYINPUT65), .Z(n356) );
  OR2_X1 U486 ( .A1(n608), .A2(n675), .ZN(n357) );
  XOR2_X1 U487 ( .A(n611), .B(KEYINPUT59), .Z(n358) );
  XNOR2_X1 U488 ( .A(KEYINPUT62), .B(KEYINPUT86), .ZN(n359) );
  NOR2_X1 U489 ( .A1(n727), .A2(G952), .ZN(n703) );
  INV_X1 U490 ( .A(n703), .ZN(n389) );
  XNOR2_X1 U491 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n360) );
  INV_X1 U492 ( .A(G472), .ZN(n412) );
  XNOR2_X1 U493 ( .A(n443), .B(G104), .ZN(n444) );
  XNOR2_X1 U494 ( .A(n444), .B(n446), .ZN(n393) );
  NAND2_X1 U495 ( .A1(n586), .A2(n365), .ZN(n361) );
  XNOR2_X1 U496 ( .A(n397), .B(KEYINPUT48), .ZN(n396) );
  XNOR2_X2 U497 ( .A(n364), .B(n588), .ZN(n731) );
  NAND2_X1 U498 ( .A1(n380), .A2(n383), .ZN(n364) );
  AND2_X2 U499 ( .A1(n418), .A2(n357), .ZN(n610) );
  XNOR2_X2 U500 ( .A(n569), .B(n568), .ZN(n586) );
  NAND2_X1 U501 ( .A1(n384), .A2(n587), .ZN(n381) );
  NOR2_X1 U502 ( .A1(n575), .A2(n582), .ZN(n590) );
  NAND2_X1 U503 ( .A1(n376), .A2(n604), .ZN(n375) );
  XNOR2_X1 U504 ( .A(n375), .B(n356), .ZN(n605) );
  XNOR2_X1 U505 ( .A(n473), .B(G137), .ZN(n442) );
  XNOR2_X1 U506 ( .A(n442), .B(n455), .ZN(n720) );
  NAND2_X1 U507 ( .A1(n379), .A2(n378), .ZN(n377) );
  NOR2_X1 U508 ( .A1(n382), .A2(n381), .ZN(n380) );
  XNOR2_X1 U509 ( .A(n367), .B(n615), .ZN(G60) );
  NOR2_X2 U510 ( .A1(n613), .A2(n703), .ZN(n367) );
  NAND2_X1 U511 ( .A1(n598), .A2(KEYINPUT34), .ZN(n384) );
  XNOR2_X1 U512 ( .A(n368), .B(n689), .ZN(G51) );
  NOR2_X2 U513 ( .A1(n688), .A2(n703), .ZN(n368) );
  NAND2_X1 U514 ( .A1(n371), .A2(n377), .ZN(n376) );
  NAND2_X1 U515 ( .A1(n589), .A2(n731), .ZN(n371) );
  NAND2_X1 U516 ( .A1(n605), .A2(n606), .ZN(n607) );
  INV_X1 U517 ( .A(n731), .ZN(n379) );
  XNOR2_X2 U518 ( .A(n585), .B(n584), .ZN(n669) );
  INV_X1 U519 ( .A(n598), .ZN(n386) );
  NOR2_X1 U520 ( .A1(G902), .A2(n697), .ZN(n461) );
  XNOR2_X2 U521 ( .A(n448), .B(n447), .ZN(n530) );
  XNOR2_X2 U522 ( .A(n530), .B(KEYINPUT1), .ZN(n642) );
  NAND2_X1 U523 ( .A1(n524), .A2(n525), .ZN(n548) );
  NAND2_X1 U524 ( .A1(n411), .A2(n405), .ZN(n404) );
  NOR2_X1 U525 ( .A1(n407), .A2(n404), .ZN(n521) );
  NOR2_X1 U526 ( .A1(n547), .A2(n656), .ZN(n538) );
  NAND2_X1 U527 ( .A1(n567), .A2(n566), .ZN(n569) );
  INV_X1 U528 ( .A(n532), .ZN(n414) );
  NAND2_X1 U529 ( .A1(n532), .A2(KEYINPUT19), .ZN(n417) );
  XNOR2_X2 U530 ( .A(n438), .B(n437), .ZN(n532) );
  INV_X1 U531 ( .A(n605), .ZN(n676) );
  NAND2_X1 U532 ( .A1(n419), .A2(n609), .ZN(n418) );
  XNOR2_X1 U533 ( .A(n607), .B(KEYINPUT81), .ZN(n419) );
  XNOR2_X1 U534 ( .A(n445), .B(n435), .ZN(n420) );
  XNOR2_X2 U535 ( .A(n513), .B(n423), .ZN(n706) );
  XNOR2_X2 U536 ( .A(n428), .B(n427), .ZN(n513) );
  XNOR2_X1 U537 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U538 ( .A(n479), .B(n466), .ZN(n469) );
  INV_X1 U539 ( .A(G119), .ZN(n425) );
  XNOR2_X1 U540 ( .A(n470), .B(G140), .ZN(n471) );
  XNOR2_X1 U541 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U542 ( .A(n612), .B(n358), .ZN(n613) );
  XNOR2_X1 U543 ( .A(n614), .B(KEYINPUT60), .ZN(n615) );
  INV_X1 U544 ( .A(n499), .ZN(n727) );
  XNOR2_X2 U545 ( .A(KEYINPUT88), .B(KEYINPUT3), .ZN(n426) );
  XOR2_X1 U546 ( .A(G113), .B(G116), .Z(n427) );
  XOR2_X2 U547 ( .A(G107), .B(G110), .Z(n704) );
  XNOR2_X1 U548 ( .A(n506), .B(KEYINPUT73), .ZN(n429) );
  XOR2_X1 U549 ( .A(n441), .B(KEYINPUT18), .Z(n432) );
  NAND2_X1 U550 ( .A1(G224), .A2(n727), .ZN(n431) );
  XNOR2_X1 U551 ( .A(n462), .B(KEYINPUT89), .ZN(n434) );
  NAND2_X1 U552 ( .A1(n685), .A2(n608), .ZN(n438) );
  NAND2_X1 U553 ( .A1(G210), .A2(n439), .ZN(n437) );
  NAND2_X1 U554 ( .A1(n439), .A2(G214), .ZN(n440) );
  XOR2_X1 U555 ( .A(KEYINPUT90), .B(n440), .Z(n656) );
  XNOR2_X1 U556 ( .A(G131), .B(KEYINPUT68), .ZN(n473) );
  XNOR2_X1 U557 ( .A(G146), .B(n720), .ZN(n512) );
  NAND2_X1 U558 ( .A1(G227), .A2(n727), .ZN(n446) );
  XNOR2_X1 U559 ( .A(n478), .B(KEYINPUT94), .ZN(n443) );
  XNOR2_X1 U560 ( .A(KEYINPUT71), .B(G469), .ZN(n447) );
  INV_X1 U561 ( .A(n642), .ZN(n591) );
  XOR2_X1 U562 ( .A(KEYINPUT102), .B(KEYINPUT101), .Z(n450) );
  XNOR2_X1 U563 ( .A(G122), .B(KEYINPUT104), .ZN(n449) );
  XNOR2_X1 U564 ( .A(n450), .B(n449), .ZN(n454) );
  XOR2_X1 U565 ( .A(KEYINPUT9), .B(KEYINPUT103), .Z(n452) );
  XNOR2_X1 U566 ( .A(KEYINPUT105), .B(KEYINPUT7), .ZN(n451) );
  XNOR2_X1 U567 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U568 ( .A(n454), .B(n453), .ZN(n460) );
  XOR2_X1 U569 ( .A(G116), .B(n456), .Z(n459) );
  NAND2_X1 U570 ( .A1(n727), .A2(G234), .ZN(n457) );
  XOR2_X1 U571 ( .A(KEYINPUT8), .B(n457), .Z(n477) );
  NAND2_X1 U572 ( .A1(G217), .A2(n477), .ZN(n458) );
  XOR2_X1 U573 ( .A(KEYINPUT11), .B(KEYINPUT99), .Z(n464) );
  XNOR2_X1 U574 ( .A(KEYINPUT98), .B(KEYINPUT12), .ZN(n463) );
  XNOR2_X1 U575 ( .A(n464), .B(n463), .ZN(n465) );
  INV_X1 U576 ( .A(n467), .ZN(n468) );
  XNOR2_X1 U577 ( .A(n469), .B(n468), .ZN(n472) );
  XNOR2_X1 U578 ( .A(G113), .B(G143), .ZN(n470) );
  XNOR2_X1 U579 ( .A(KEYINPUT13), .B(G475), .ZN(n474) );
  INV_X1 U580 ( .A(n551), .ZN(n534) );
  INV_X1 U581 ( .A(n631), .ZN(n516) );
  NAND2_X1 U582 ( .A1(n477), .A2(G221), .ZN(n488) );
  XNOR2_X1 U583 ( .A(n479), .B(n478), .ZN(n719) );
  XOR2_X1 U584 ( .A(G110), .B(G137), .Z(n481) );
  XNOR2_X1 U585 ( .A(n481), .B(n480), .ZN(n485) );
  XOR2_X1 U586 ( .A(KEYINPUT95), .B(KEYINPUT24), .Z(n483) );
  XNOR2_X1 U587 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U588 ( .A(n488), .B(n487), .ZN(n701) );
  NOR2_X1 U589 ( .A1(n701), .A2(G902), .ZN(n492) );
  XOR2_X1 U590 ( .A(KEYINPUT77), .B(KEYINPUT25), .Z(n491) );
  NAND2_X1 U591 ( .A1(n608), .A2(G234), .ZN(n489) );
  XNOR2_X1 U592 ( .A(n489), .B(KEYINPUT20), .ZN(n493) );
  NAND2_X1 U593 ( .A1(n493), .A2(G217), .ZN(n490) );
  INV_X1 U594 ( .A(n577), .ZN(n505) );
  NAND2_X1 U595 ( .A1(n493), .A2(G221), .ZN(n494) );
  XOR2_X1 U596 ( .A(n494), .B(KEYINPUT21), .Z(n639) );
  INV_X1 U597 ( .A(n639), .ZN(n570) );
  XNOR2_X1 U598 ( .A(n496), .B(n495), .ZN(n498) );
  NAND2_X1 U599 ( .A1(n498), .A2(G952), .ZN(n497) );
  XOR2_X1 U600 ( .A(KEYINPUT92), .B(n497), .Z(n668) );
  NAND2_X1 U601 ( .A1(n709), .A2(n668), .ZN(n564) );
  NAND2_X1 U602 ( .A1(G902), .A2(n498), .ZN(n562) );
  NOR2_X1 U603 ( .A1(G900), .A2(n562), .ZN(n500) );
  NAND2_X1 U604 ( .A1(n500), .A2(n499), .ZN(n501) );
  NAND2_X1 U605 ( .A1(n564), .A2(n501), .ZN(n502) );
  XOR2_X1 U606 ( .A(KEYINPUT78), .B(n502), .Z(n523) );
  XOR2_X1 U607 ( .A(KEYINPUT70), .B(n503), .Z(n504) );
  NOR2_X1 U608 ( .A1(n505), .A2(n504), .ZN(n528) );
  INV_X1 U609 ( .A(KEYINPUT6), .ZN(n514) );
  XNOR2_X1 U610 ( .A(n506), .B(KEYINPUT76), .ZN(n507) );
  XOR2_X1 U611 ( .A(n507), .B(KEYINPUT5), .Z(n510) );
  NAND2_X1 U612 ( .A1(n508), .A2(G210), .ZN(n509) );
  NAND2_X1 U613 ( .A1(n528), .A2(n582), .ZN(n515) );
  NAND2_X1 U614 ( .A1(n591), .A2(n537), .ZN(n517) );
  NOR2_X1 U615 ( .A1(n656), .A2(n517), .ZN(n518) );
  XNOR2_X1 U616 ( .A(n518), .B(KEYINPUT43), .ZN(n519) );
  NOR2_X1 U617 ( .A1(n414), .A2(n519), .ZN(n520) );
  XNOR2_X1 U618 ( .A(KEYINPUT110), .B(n520), .ZN(n733) );
  NAND2_X1 U619 ( .A1(n530), .A2(n643), .ZN(n600) );
  XNOR2_X1 U620 ( .A(KEYINPUT111), .B(n600), .ZN(n525) );
  XOR2_X1 U621 ( .A(KEYINPUT30), .B(n521), .Z(n522) );
  NOR2_X1 U622 ( .A1(n523), .A2(n522), .ZN(n524) );
  NOR2_X1 U623 ( .A1(n547), .A2(n548), .ZN(n526) );
  XNOR2_X1 U624 ( .A(KEYINPUT112), .B(n526), .ZN(n527) );
  NOR2_X1 U625 ( .A1(n552), .A2(n551), .ZN(n587) );
  NAND2_X1 U626 ( .A1(n527), .A2(n587), .ZN(n628) );
  AND2_X1 U627 ( .A1(n528), .A2(n649), .ZN(n529) );
  XNOR2_X1 U628 ( .A(KEYINPUT28), .B(n529), .ZN(n531) );
  NAND2_X1 U629 ( .A1(n531), .A2(n530), .ZN(n555) );
  INV_X1 U630 ( .A(n567), .ZN(n533) );
  NOR2_X1 U631 ( .A1(n555), .A2(n533), .ZN(n629) );
  XOR2_X1 U632 ( .A(KEYINPUT107), .B(n633), .Z(n560) );
  NOR2_X1 U633 ( .A1(n631), .A2(n560), .ZN(n602) );
  INV_X1 U634 ( .A(n602), .ZN(n660) );
  NAND2_X1 U635 ( .A1(n629), .A2(n660), .ZN(n542) );
  NAND2_X1 U636 ( .A1(KEYINPUT47), .A2(n542), .ZN(n535) );
  NAND2_X1 U637 ( .A1(n628), .A2(n535), .ZN(n536) );
  XNOR2_X1 U638 ( .A(n536), .B(KEYINPUT79), .ZN(n546) );
  XOR2_X1 U639 ( .A(KEYINPUT36), .B(KEYINPUT115), .Z(n540) );
  NAND2_X1 U640 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U641 ( .A(n540), .B(n539), .ZN(n541) );
  NOR2_X1 U642 ( .A1(n591), .A2(n541), .ZN(n636) );
  XNOR2_X1 U643 ( .A(KEYINPUT74), .B(n543), .ZN(n544) );
  NOR2_X1 U644 ( .A1(n636), .A2(n544), .ZN(n545) );
  NAND2_X1 U645 ( .A1(n546), .A2(n545), .ZN(n559) );
  XNOR2_X1 U646 ( .A(KEYINPUT113), .B(KEYINPUT40), .ZN(n549) );
  XNOR2_X1 U647 ( .A(n550), .B(n549), .ZN(n737) );
  XOR2_X1 U648 ( .A(KEYINPUT114), .B(KEYINPUT41), .Z(n554) );
  NAND2_X1 U649 ( .A1(n659), .A2(n657), .ZN(n553) );
  XNOR2_X1 U650 ( .A(n554), .B(n553), .ZN(n670) );
  NOR2_X1 U651 ( .A1(n670), .A2(n555), .ZN(n556) );
  XOR2_X1 U652 ( .A(KEYINPUT42), .B(n556), .Z(n735) );
  NAND2_X1 U653 ( .A1(n737), .A2(n735), .ZN(n557) );
  XNOR2_X1 U654 ( .A(n557), .B(KEYINPUT46), .ZN(n558) );
  NAND2_X1 U655 ( .A1(n561), .A2(n560), .ZN(n638) );
  INV_X1 U656 ( .A(n608), .ZN(n606) );
  NOR2_X1 U657 ( .A1(KEYINPUT44), .A2(KEYINPUT83), .ZN(n580) );
  NOR2_X1 U658 ( .A1(G898), .A2(n709), .ZN(n708) );
  INV_X1 U659 ( .A(n562), .ZN(n563) );
  NAND2_X1 U660 ( .A1(n708), .A2(n563), .ZN(n565) );
  NAND2_X1 U661 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U662 ( .A(KEYINPUT84), .B(KEYINPUT0), .Z(n568) );
  XOR2_X1 U663 ( .A(KEYINPUT108), .B(n577), .Z(n640) );
  NOR2_X1 U664 ( .A1(n591), .A2(n640), .ZN(n571) );
  NAND2_X1 U665 ( .A1(n590), .A2(n571), .ZN(n572) );
  NAND2_X1 U666 ( .A1(n591), .A2(n573), .ZN(n574) );
  XNOR2_X1 U667 ( .A(KEYINPUT66), .B(n576), .ZN(n578) );
  NAND2_X1 U668 ( .A1(n578), .A2(n577), .ZN(n622) );
  NAND2_X1 U669 ( .A1(n734), .A2(n622), .ZN(n579) );
  XNOR2_X1 U670 ( .A(n580), .B(n579), .ZN(n589) );
  NAND2_X1 U671 ( .A1(n642), .A2(n643), .ZN(n581) );
  INV_X1 U672 ( .A(KEYINPUT33), .ZN(n583) );
  INV_X1 U673 ( .A(KEYINPUT35), .ZN(n588) );
  AND2_X1 U674 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U675 ( .A1(n640), .A2(n592), .ZN(n593) );
  XNOR2_X1 U676 ( .A(KEYINPUT109), .B(n593), .ZN(n732) );
  NAND2_X1 U677 ( .A1(n649), .A2(n594), .ZN(n595) );
  XNOR2_X1 U678 ( .A(KEYINPUT97), .B(n595), .ZN(n651) );
  NAND2_X1 U679 ( .A1(n651), .A2(n596), .ZN(n597) );
  XNOR2_X1 U680 ( .A(n597), .B(KEYINPUT31), .ZN(n634) );
  OR2_X1 U681 ( .A1(n598), .A2(n649), .ZN(n599) );
  NOR2_X1 U682 ( .A1(n600), .A2(n599), .ZN(n618) );
  NOR2_X1 U683 ( .A1(n634), .A2(n618), .ZN(n601) );
  NOR2_X1 U684 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U685 ( .A1(n732), .A2(n603), .ZN(n604) );
  INV_X1 U686 ( .A(KEYINPUT2), .ZN(n675) );
  INV_X1 U687 ( .A(n676), .ZN(n710) );
  NAND2_X1 U688 ( .A1(n693), .A2(G475), .ZN(n612) );
  INV_X1 U689 ( .A(KEYINPUT123), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n618), .A2(n631), .ZN(n617) );
  XNOR2_X1 U691 ( .A(G104), .B(n617), .ZN(G6) );
  XOR2_X1 U692 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n620) );
  NAND2_X1 U693 ( .A1(n618), .A2(n633), .ZN(n619) );
  XNOR2_X1 U694 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U695 ( .A(G107), .B(n621), .ZN(G9) );
  XNOR2_X1 U696 ( .A(n622), .B(G110), .ZN(G12) );
  XOR2_X1 U697 ( .A(KEYINPUT29), .B(KEYINPUT118), .Z(n624) );
  XNOR2_X1 U698 ( .A(G128), .B(KEYINPUT117), .ZN(n623) );
  XNOR2_X1 U699 ( .A(n624), .B(n623), .ZN(n625) );
  XOR2_X1 U700 ( .A(KEYINPUT116), .B(n625), .Z(n627) );
  NAND2_X1 U701 ( .A1(n629), .A2(n633), .ZN(n626) );
  XNOR2_X1 U702 ( .A(n627), .B(n626), .ZN(G30) );
  XNOR2_X1 U703 ( .A(G143), .B(n628), .ZN(G45) );
  NAND2_X1 U704 ( .A1(n631), .A2(n629), .ZN(n630) );
  XNOR2_X1 U705 ( .A(n630), .B(G146), .ZN(G48) );
  NAND2_X1 U706 ( .A1(n631), .A2(n634), .ZN(n632) );
  XNOR2_X1 U707 ( .A(n632), .B(G113), .ZN(G15) );
  NAND2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U709 ( .A(n635), .B(G116), .ZN(G18) );
  XNOR2_X1 U710 ( .A(G125), .B(n636), .ZN(n637) );
  XNOR2_X1 U711 ( .A(n637), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U712 ( .A(G134), .B(n638), .ZN(G36) );
  NOR2_X1 U713 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U714 ( .A(KEYINPUT49), .B(n641), .ZN(n647) );
  NOR2_X1 U715 ( .A1(n643), .A2(n642), .ZN(n645) );
  XNOR2_X1 U716 ( .A(KEYINPUT50), .B(KEYINPUT119), .ZN(n644) );
  XNOR2_X1 U717 ( .A(n645), .B(n644), .ZN(n646) );
  NAND2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U719 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U720 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U721 ( .A(n652), .B(KEYINPUT51), .Z(n653) );
  XNOR2_X1 U722 ( .A(KEYINPUT120), .B(n653), .ZN(n654) );
  NOR2_X1 U723 ( .A1(n670), .A2(n654), .ZN(n665) );
  NAND2_X1 U724 ( .A1(n656), .A2(n655), .ZN(n658) );
  NAND2_X1 U725 ( .A1(n658), .A2(n657), .ZN(n662) );
  NAND2_X1 U726 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U727 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U728 ( .A1(n663), .A2(n669), .ZN(n664) );
  NOR2_X1 U729 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U730 ( .A(KEYINPUT52), .B(n666), .Z(n667) );
  AND2_X1 U731 ( .A1(n668), .A2(n667), .ZN(n672) );
  NOR2_X1 U732 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U733 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U734 ( .A(n673), .B(KEYINPUT121), .ZN(n682) );
  NAND2_X1 U735 ( .A1(n726), .A2(n675), .ZN(n674) );
  XNOR2_X1 U736 ( .A(n674), .B(KEYINPUT80), .ZN(n678) );
  NAND2_X1 U737 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U738 ( .A1(n678), .A2(n677), .ZN(n680) );
  NOR2_X1 U739 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U740 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U741 ( .A1(n709), .A2(n683), .ZN(n684) );
  XOR2_X1 U742 ( .A(KEYINPUT53), .B(n684), .Z(G75) );
  NAND2_X1 U743 ( .A1(n693), .A2(G210), .ZN(n687) );
  XNOR2_X1 U744 ( .A(n685), .B(n360), .ZN(n686) );
  XNOR2_X1 U745 ( .A(KEYINPUT82), .B(KEYINPUT56), .ZN(n689) );
  XNOR2_X1 U746 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n692) );
  XNOR2_X1 U747 ( .A(n690), .B(KEYINPUT57), .ZN(n691) );
  XNOR2_X1 U748 ( .A(n692), .B(n691), .ZN(n695) );
  NAND2_X1 U749 ( .A1(n699), .A2(G469), .ZN(n694) );
  NAND2_X1 U750 ( .A1(n699), .A2(G478), .ZN(n696) );
  XNOR2_X1 U751 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X1 U752 ( .A1(n703), .A2(n698), .ZN(G63) );
  NAND2_X1 U753 ( .A1(n699), .A2(G217), .ZN(n700) );
  XNOR2_X1 U754 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U755 ( .A1(n703), .A2(n702), .ZN(G66) );
  XOR2_X1 U756 ( .A(G101), .B(n704), .Z(n705) );
  XNOR2_X1 U757 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U758 ( .A1(n708), .A2(n707), .ZN(n718) );
  NAND2_X1 U759 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U760 ( .A(n711), .B(KEYINPUT124), .ZN(n715) );
  NAND2_X1 U761 ( .A1(G953), .A2(G224), .ZN(n712) );
  XNOR2_X1 U762 ( .A(KEYINPUT61), .B(n712), .ZN(n713) );
  NAND2_X1 U763 ( .A1(n713), .A2(G898), .ZN(n714) );
  NAND2_X1 U764 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U765 ( .A(n716), .B(KEYINPUT125), .Z(n717) );
  XNOR2_X1 U766 ( .A(n718), .B(n717), .ZN(G69) );
  XNOR2_X1 U767 ( .A(KEYINPUT4), .B(n719), .ZN(n721) );
  XOR2_X1 U768 ( .A(n721), .B(n720), .Z(n725) );
  XOR2_X1 U769 ( .A(KEYINPUT126), .B(n725), .Z(n722) );
  XNOR2_X1 U770 ( .A(G227), .B(n722), .ZN(n723) );
  NAND2_X1 U771 ( .A1(n723), .A2(G900), .ZN(n724) );
  NAND2_X1 U772 ( .A1(n724), .A2(G953), .ZN(n730) );
  XOR2_X1 U773 ( .A(n726), .B(n725), .Z(n728) );
  NAND2_X1 U774 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U775 ( .A1(n730), .A2(n729), .ZN(G72) );
  XNOR2_X1 U776 ( .A(G122), .B(n731), .ZN(G24) );
  XOR2_X1 U777 ( .A(G101), .B(n732), .Z(G3) );
  XOR2_X1 U778 ( .A(G140), .B(n733), .Z(G42) );
  XNOR2_X1 U779 ( .A(n734), .B(G119), .ZN(G21) );
  XOR2_X1 U780 ( .A(n735), .B(G137), .Z(n736) );
  XNOR2_X1 U781 ( .A(KEYINPUT127), .B(n736), .ZN(G39) );
  XNOR2_X1 U782 ( .A(G131), .B(n737), .ZN(G33) );
endmodule

