

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793;

  OR2_X1 U364 ( .A1(n676), .A2(n474), .ZN(n473) );
  XNOR2_X1 U365 ( .A(n368), .B(n525), .ZN(n676) );
  AND2_X2 U366 ( .A1(n556), .A2(n445), .ZN(n587) );
  NAND2_X1 U367 ( .A1(n343), .A2(n659), .ZN(n446) );
  NAND2_X1 U368 ( .A1(n367), .A2(n782), .ZN(n343) );
  XOR2_X1 U369 ( .A(KEYINPUT72), .B(n611), .Z(n344) );
  AND2_X2 U370 ( .A1(n406), .A2(n404), .ZN(n366) );
  AND2_X2 U371 ( .A1(n373), .A2(n350), .ZN(n372) );
  AND2_X2 U372 ( .A1(n364), .A2(n363), .ZN(n612) );
  XNOR2_X2 U373 ( .A(n577), .B(n397), .ZN(n364) );
  NOR2_X2 U374 ( .A1(n747), .A2(n589), .ZN(n583) );
  NOR2_X1 U375 ( .A1(n417), .A2(n452), .ZN(n416) );
  INV_X2 U376 ( .A(n620), .ZN(n345) );
  INV_X1 U377 ( .A(G110), .ZN(n447) );
  AND2_X1 U378 ( .A1(n668), .A2(n696), .ZN(n496) );
  AND2_X1 U379 ( .A1(n697), .A2(n696), .ZN(n495) );
  XNOR2_X1 U380 ( .A(n365), .B(n361), .ZN(n417) );
  AND2_X1 U381 ( .A1(n434), .A2(n433), .ZN(n428) );
  NOR2_X1 U382 ( .A1(n652), .A2(n444), .ZN(n431) );
  XNOR2_X1 U383 ( .A(n587), .B(n399), .ZN(n408) );
  NAND2_X1 U384 ( .A1(n348), .A2(n633), .ZN(n453) );
  NOR2_X2 U385 ( .A1(n793), .A2(n792), .ZN(n427) );
  XNOR2_X1 U386 ( .A(n591), .B(n590), .ZN(n714) );
  OR2_X1 U387 ( .A1(n670), .A2(G902), .ZN(n493) );
  XNOR2_X1 U388 ( .A(n364), .B(n396), .ZN(n727) );
  XNOR2_X1 U389 ( .A(n394), .B(n393), .ZN(n596) );
  XNOR2_X1 U390 ( .A(n542), .B(n504), .ZN(n779) );
  OR2_X1 U391 ( .A1(n694), .A2(G902), .ZN(n490) );
  XNOR2_X1 U392 ( .A(n447), .B(G119), .ZN(n516) );
  XNOR2_X1 U393 ( .A(n513), .B(KEYINPUT10), .ZN(n542) );
  XNOR2_X1 U394 ( .A(n521), .B(n520), .ZN(n549) );
  XNOR2_X1 U395 ( .A(G146), .B(G125), .ZN(n513) );
  INV_X2 U396 ( .A(G953), .ZN(n783) );
  XNOR2_X1 U397 ( .A(G128), .B(KEYINPUT85), .ZN(n505) );
  XNOR2_X1 U398 ( .A(G122), .B(G116), .ZN(n521) );
  NAND2_X1 U399 ( .A1(G237), .A2(G234), .ZN(n532) );
  NOR2_X2 U400 ( .A1(n410), .A2(n416), .ZN(n346) );
  BUF_X1 U401 ( .A(n557), .Z(n347) );
  NOR2_X1 U402 ( .A1(n410), .A2(n416), .ZN(n782) );
  XNOR2_X2 U403 ( .A(n490), .B(n351), .ZN(n597) );
  AND2_X2 U404 ( .A1(n409), .A2(KEYINPUT28), .ZN(n353) );
  NOR2_X4 U405 ( .A1(n643), .A2(n642), .ZN(n647) );
  XNOR2_X2 U406 ( .A(n625), .B(KEYINPUT104), .ZN(n643) );
  NAND2_X1 U407 ( .A1(n475), .A2(n509), .ZN(n474) );
  AND2_X1 U408 ( .A1(n737), .A2(n443), .ZN(n441) );
  XNOR2_X1 U409 ( .A(n463), .B(n461), .ZN(n515) );
  XNOR2_X1 U410 ( .A(n462), .B(KEYINPUT83), .ZN(n461) );
  AND2_X1 U411 ( .A1(n644), .A2(n390), .ZN(n389) );
  INV_X1 U412 ( .A(n702), .ZN(n391) );
  NOR2_X1 U413 ( .A1(G902), .A2(G237), .ZN(n526) );
  NAND2_X1 U414 ( .A1(n403), .A2(n401), .ZN(n400) );
  INV_X1 U415 ( .A(n790), .ZN(n403) );
  NAND2_X1 U416 ( .A1(n592), .A2(KEYINPUT30), .ZN(n437) );
  NAND2_X1 U417 ( .A1(n467), .A2(KEYINPUT30), .ZN(n439) );
  INV_X1 U418 ( .A(n470), .ZN(n464) );
  NAND2_X1 U419 ( .A1(n737), .A2(KEYINPUT19), .ZN(n470) );
  NAND2_X1 U420 ( .A1(n567), .A2(n481), .ZN(n480) );
  NAND2_X1 U421 ( .A1(n413), .A2(n411), .ZN(n410) );
  NOR2_X1 U422 ( .A1(n412), .A2(n720), .ZN(n411) );
  INV_X1 U423 ( .A(KEYINPUT82), .ZN(n522) );
  XNOR2_X1 U424 ( .A(n497), .B(n488), .ZN(n548) );
  INV_X1 U425 ( .A(KEYINPUT8), .ZN(n488) );
  INV_X1 U426 ( .A(KEYINPUT100), .ZN(n424) );
  XNOR2_X1 U427 ( .A(n511), .B(n354), .ZN(n492) );
  AND2_X1 U428 ( .A1(n473), .A2(n531), .ZN(n472) );
  OR2_X1 U429 ( .A1(n774), .A2(G902), .ZN(n394) );
  BUF_X1 U430 ( .A(n727), .Z(n448) );
  NAND2_X1 U431 ( .A1(n430), .A2(n709), .ZN(n653) );
  INV_X1 U432 ( .A(KEYINPUT66), .ZN(n444) );
  INV_X1 U433 ( .A(KEYINPUT94), .ZN(n390) );
  NOR2_X1 U434 ( .A1(n453), .A2(n452), .ZN(n412) );
  NAND2_X1 U435 ( .A1(n417), .A2(n414), .ZN(n413) );
  NOR2_X1 U436 ( .A1(n415), .A2(KEYINPUT76), .ZN(n414) );
  INV_X1 U437 ( .A(n453), .ZN(n415) );
  XNOR2_X1 U438 ( .A(G131), .B(G134), .ZN(n558) );
  NAND2_X1 U439 ( .A1(n383), .A2(n382), .ZN(n601) );
  AND2_X1 U440 ( .A1(n388), .A2(n384), .ZN(n383) );
  XNOR2_X1 U441 ( .A(G110), .B(G101), .ZN(n569) );
  XOR2_X1 U442 ( .A(KEYINPUT70), .B(G107), .Z(n570) );
  XNOR2_X1 U443 ( .A(n572), .B(n355), .ZN(n449) );
  XNOR2_X1 U444 ( .A(n503), .B(n502), .ZN(n573) );
  INV_X1 U445 ( .A(KEYINPUT65), .ZN(n502) );
  INV_X1 U446 ( .A(KEYINPUT1), .ZN(n396) );
  BUF_X1 U447 ( .A(n747), .Z(n420) );
  XNOR2_X1 U448 ( .A(n615), .B(n614), .ZN(n657) );
  NOR2_X1 U449 ( .A1(n436), .A2(n435), .ZN(n613) );
  AND2_X1 U450 ( .A1(n628), .A2(n711), .ZN(n629) );
  XNOR2_X1 U451 ( .A(n612), .B(KEYINPUT102), .ZN(n637) );
  NAND2_X1 U452 ( .A1(n596), .A2(n597), .ZN(n627) );
  NAND2_X1 U453 ( .A1(n372), .A2(n369), .ZN(n593) );
  XNOR2_X1 U454 ( .A(n524), .B(n523), .ZN(n368) );
  XNOR2_X1 U455 ( .A(n549), .B(n486), .ZN(n485) );
  XNOR2_X1 U456 ( .A(n547), .B(n544), .ZN(n486) );
  AND2_X2 U457 ( .A1(n663), .A2(n662), .ZN(n771) );
  XNOR2_X1 U458 ( .A(n446), .B(KEYINPUT64), .ZN(n663) );
  NOR2_X1 U459 ( .A1(n586), .A2(n345), .ZN(n445) );
  INV_X1 U460 ( .A(n683), .ZN(n398) );
  INV_X1 U461 ( .A(KEYINPUT44), .ZN(n407) );
  NOR2_X1 U462 ( .A1(n386), .A2(n385), .ZN(n384) );
  NOR2_X1 U463 ( .A1(n644), .A2(n390), .ZN(n385) );
  NOR2_X1 U464 ( .A1(n391), .A2(n387), .ZN(n386) );
  NAND2_X1 U465 ( .A1(n528), .A2(n658), .ZN(n477) );
  INV_X1 U466 ( .A(G902), .ZN(n481) );
  NAND2_X1 U467 ( .A1(G472), .A2(G902), .ZN(n483) );
  NOR2_X1 U468 ( .A1(G953), .A2(G237), .ZN(n561) );
  XNOR2_X1 U469 ( .A(G137), .B(G119), .ZN(n559) );
  XOR2_X1 U470 ( .A(KEYINPUT5), .B(G116), .Z(n560) );
  XNOR2_X1 U471 ( .A(G140), .B(G113), .ZN(n539) );
  XNOR2_X1 U472 ( .A(n540), .B(n459), .ZN(n458) );
  XNOR2_X1 U473 ( .A(n541), .B(KEYINPUT12), .ZN(n459) );
  XNOR2_X1 U474 ( .A(G143), .B(G131), .ZN(n541) );
  XNOR2_X1 U475 ( .A(n538), .B(n537), .ZN(n457) );
  NAND2_X1 U476 ( .A1(n783), .A2(G224), .ZN(n462) );
  XNOR2_X1 U477 ( .A(n513), .B(n512), .ZN(n463) );
  XNOR2_X1 U478 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n512) );
  NAND2_X1 U479 ( .A1(n738), .A2(n349), .ZN(n435) );
  INV_X1 U480 ( .A(n596), .ZN(n595) );
  OR2_X1 U481 ( .A1(n380), .A2(n494), .ZN(n371) );
  NAND2_X1 U482 ( .A1(n374), .A2(n494), .ZN(n373) );
  INV_X1 U483 ( .A(n378), .ZN(n375) );
  AND2_X1 U484 ( .A1(n601), .A2(n699), .ZN(n602) );
  INV_X1 U485 ( .A(G101), .ZN(n517) );
  XOR2_X1 U486 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n547) );
  INV_X1 U487 ( .A(G107), .ZN(n520) );
  XNOR2_X1 U488 ( .A(n456), .B(n454), .ZN(n694) );
  XNOR2_X1 U489 ( .A(n542), .B(n455), .ZN(n454) );
  XNOR2_X1 U490 ( .A(n458), .B(n457), .ZN(n456) );
  XNOR2_X1 U491 ( .A(n543), .B(n539), .ZN(n455) );
  NAND2_X1 U492 ( .A1(n658), .A2(KEYINPUT2), .ZN(n659) );
  XNOR2_X1 U493 ( .A(n571), .B(n449), .ZN(n574) );
  XNOR2_X1 U494 ( .A(n582), .B(n581), .ZN(n747) );
  NAND2_X1 U495 ( .A1(n440), .A2(n349), .ZN(n438) );
  INV_X1 U496 ( .A(KEYINPUT22), .ZN(n418) );
  XNOR2_X1 U497 ( .A(n779), .B(KEYINPUT24), .ZN(n451) );
  XNOR2_X1 U498 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U499 ( .A(KEYINPUT101), .B(KEYINPUT43), .ZN(n421) );
  NAND2_X1 U500 ( .A1(n423), .A2(n448), .ZN(n422) );
  NOR2_X1 U501 ( .A1(n657), .A2(n627), .ZN(n616) );
  OR2_X1 U502 ( .A1(n731), .A2(n589), .ZN(n591) );
  OR2_X1 U503 ( .A1(n376), .A2(n381), .ZN(n642) );
  INV_X1 U504 ( .A(n468), .ZN(n381) );
  XNOR2_X1 U505 ( .A(n776), .B(n775), .ZN(n777) );
  INV_X1 U506 ( .A(G119), .ZN(n682) );
  INV_X1 U507 ( .A(n408), .ZN(n684) );
  XOR2_X1 U508 ( .A(n422), .B(n421), .Z(n348) );
  AND2_X1 U509 ( .A1(n344), .A2(n439), .ZN(n349) );
  OR2_X1 U510 ( .A1(n468), .A2(n379), .ZN(n350) );
  XOR2_X1 U511 ( .A(KEYINPUT13), .B(G475), .Z(n351) );
  OR2_X1 U512 ( .A1(n536), .A2(n610), .ZN(n352) );
  NAND2_X1 U513 ( .A1(n469), .A2(n466), .ZN(n380) );
  XOR2_X1 U514 ( .A(KEYINPUT69), .B(KEYINPUT25), .Z(n354) );
  AND2_X1 U515 ( .A1(G227), .A2(n783), .ZN(n355) );
  AND2_X1 U516 ( .A1(n548), .A2(G221), .ZN(n356) );
  NOR2_X1 U517 ( .A1(n725), .A2(n409), .ZN(n357) );
  OR2_X1 U518 ( .A1(n530), .A2(n529), .ZN(n737) );
  INV_X1 U519 ( .A(n737), .ZN(n467) );
  AND2_X1 U520 ( .A1(n391), .A2(KEYINPUT94), .ZN(n358) );
  XOR2_X1 U521 ( .A(KEYINPUT81), .B(n667), .Z(n778) );
  XOR2_X1 U522 ( .A(n665), .B(n664), .Z(n359) );
  XOR2_X1 U523 ( .A(n694), .B(n693), .Z(n360) );
  XNOR2_X1 U524 ( .A(KEYINPUT77), .B(KEYINPUT48), .ZN(n361) );
  NOR2_X1 U525 ( .A1(n368), .A2(n690), .ZN(n362) );
  INV_X1 U526 ( .A(KEYINPUT76), .ZN(n452) );
  NAND2_X2 U527 ( .A1(n345), .A2(n722), .ZN(n726) );
  XNOR2_X1 U528 ( .A(n507), .B(n356), .ZN(n450) );
  XNOR2_X1 U529 ( .A(n451), .B(n450), .ZN(n670) );
  INV_X1 U530 ( .A(n726), .ZN(n363) );
  NAND2_X1 U531 ( .A1(n425), .A2(n426), .ZN(n365) );
  NAND2_X1 U532 ( .A1(n366), .A2(n400), .ZN(n603) );
  XNOR2_X2 U533 ( .A(n604), .B(KEYINPUT45), .ZN(n661) );
  NAND2_X1 U534 ( .A1(n790), .A2(n407), .ZN(n406) );
  XNOR2_X2 U535 ( .A(n585), .B(KEYINPUT35), .ZN(n790) );
  XNOR2_X1 U536 ( .A(n605), .B(KEYINPUT75), .ZN(n367) );
  NAND2_X1 U537 ( .A1(n370), .A2(n468), .ZN(n369) );
  NOR2_X1 U538 ( .A1(n378), .A2(n371), .ZN(n370) );
  NAND2_X1 U539 ( .A1(n375), .A2(n377), .ZN(n374) );
  NAND2_X1 U540 ( .A1(n377), .A2(n471), .ZN(n376) );
  INV_X1 U541 ( .A(n380), .ZN(n377) );
  NAND2_X1 U542 ( .A1(n471), .A2(n352), .ZN(n378) );
  INV_X1 U543 ( .A(n494), .ZN(n379) );
  INV_X1 U544 ( .A(n714), .ZN(n392) );
  NAND2_X1 U545 ( .A1(n714), .A2(n389), .ZN(n388) );
  NAND2_X1 U546 ( .A1(n392), .A2(n358), .ZN(n382) );
  INV_X1 U547 ( .A(n389), .ZN(n387) );
  NAND2_X1 U548 ( .A1(n346), .A2(n661), .ZN(n756) );
  INV_X1 U549 ( .A(G478), .ZN(n393) );
  XNOR2_X1 U550 ( .A(n395), .B(n485), .ZN(n774) );
  XNOR2_X1 U551 ( .A(n489), .B(n487), .ZN(n395) );
  XNOR2_X1 U552 ( .A(n453), .B(G140), .ZN(G42) );
  INV_X1 U553 ( .A(G469), .ZN(n397) );
  NAND2_X1 U554 ( .A1(n408), .A2(n398), .ZN(n405) );
  XNOR2_X2 U555 ( .A(n580), .B(n579), .ZN(n683) );
  INV_X1 U556 ( .A(KEYINPUT96), .ZN(n399) );
  AND2_X1 U557 ( .A1(n408), .A2(n402), .ZN(n401) );
  NOR2_X1 U558 ( .A1(n683), .A2(n407), .ZN(n402) );
  NAND2_X1 U559 ( .A1(n405), .A2(n407), .ZN(n404) );
  INV_X1 U560 ( .A(n409), .ZN(n592) );
  NAND2_X1 U561 ( .A1(n409), .A2(n441), .ZN(n440) );
  NAND2_X1 U562 ( .A1(n628), .A2(n409), .ZN(n622) );
  XNOR2_X1 U563 ( .A(n409), .B(n568), .ZN(n630) );
  NAND2_X1 U564 ( .A1(n588), .A2(n409), .ZN(n731) );
  NAND2_X4 U565 ( .A1(n482), .A2(n479), .ZN(n409) );
  INV_X1 U566 ( .A(n556), .ZN(n600) );
  XNOR2_X2 U567 ( .A(n555), .B(n418), .ZN(n556) );
  NAND2_X1 U568 ( .A1(n419), .A2(n623), .ZN(n624) );
  NAND2_X1 U569 ( .A1(n353), .A2(n628), .ZN(n419) );
  NOR2_X1 U570 ( .A1(n765), .A2(G902), .ZN(n577) );
  XNOR2_X1 U571 ( .A(n491), .B(n424), .ZN(n423) );
  XNOR2_X1 U572 ( .A(n427), .B(KEYINPUT46), .ZN(n425) );
  NAND2_X1 U573 ( .A1(n428), .A2(n429), .ZN(n426) );
  NAND2_X1 U574 ( .A1(n431), .A2(n432), .ZN(n429) );
  XNOR2_X1 U575 ( .A(n430), .B(n718), .ZN(n719) );
  NAND2_X1 U576 ( .A1(n635), .A2(n654), .ZN(n430) );
  INV_X1 U577 ( .A(n653), .ZN(n432) );
  NAND2_X1 U578 ( .A1(n652), .A2(n444), .ZN(n433) );
  NAND2_X1 U579 ( .A1(n653), .A2(n444), .ZN(n434) );
  NAND2_X1 U580 ( .A1(n440), .A2(n437), .ZN(n436) );
  INV_X1 U581 ( .A(n437), .ZN(n442) );
  NOR2_X1 U582 ( .A1(n442), .A2(n438), .ZN(n636) );
  INV_X1 U583 ( .A(KEYINPUT30), .ZN(n443) );
  NAND2_X1 U584 ( .A1(n548), .A2(G217), .ZN(n487) );
  NAND2_X1 U585 ( .A1(n665), .A2(G472), .ZN(n484) );
  AND2_X2 U586 ( .A1(n484), .A2(n483), .ZN(n482) );
  XNOR2_X2 U587 ( .A(n627), .B(KEYINPUT97), .ZN(n711) );
  NAND2_X1 U588 ( .A1(n556), .A2(n460), .ZN(n580) );
  AND2_X1 U589 ( .A1(n620), .A2(n578), .ZN(n460) );
  INV_X1 U590 ( .A(n465), .ZN(n476) );
  NAND2_X1 U591 ( .A1(n465), .A2(n464), .ZN(n469) );
  NAND2_X1 U592 ( .A1(n478), .A2(n477), .ZN(n465) );
  NAND2_X1 U593 ( .A1(n476), .A2(n473), .ZN(n655) );
  NAND2_X1 U594 ( .A1(n467), .A2(n531), .ZN(n466) );
  OR2_X1 U595 ( .A1(n473), .A2(n470), .ZN(n468) );
  NAND2_X1 U596 ( .A1(n472), .A2(n476), .ZN(n471) );
  INV_X1 U597 ( .A(n528), .ZN(n475) );
  NAND2_X1 U598 ( .A1(n676), .A2(n528), .ZN(n478) );
  XNOR2_X2 U599 ( .A(n781), .B(G146), .ZN(n576) );
  XNOR2_X2 U600 ( .A(n557), .B(n558), .ZN(n781) );
  XNOR2_X2 U601 ( .A(n546), .B(KEYINPUT4), .ZN(n557) );
  XNOR2_X2 U602 ( .A(n514), .B(G143), .ZN(n546) );
  OR2_X2 U603 ( .A1(n665), .A2(n480), .ZN(n479) );
  XNOR2_X1 U604 ( .A(n546), .B(n545), .ZN(n489) );
  NOR2_X2 U605 ( .A1(n491), .A2(n633), .ZN(n634) );
  NAND2_X1 U606 ( .A1(n632), .A2(n737), .ZN(n491) );
  XNOR2_X2 U607 ( .A(n493), .B(n492), .ZN(n620) );
  XNOR2_X1 U608 ( .A(n774), .B(n773), .ZN(n775) );
  XOR2_X1 U609 ( .A(KEYINPUT78), .B(KEYINPUT0), .Z(n494) );
  XNOR2_X1 U610 ( .A(n516), .B(n505), .ZN(n506) );
  XNOR2_X1 U611 ( .A(KEYINPUT67), .B(KEYINPUT33), .ZN(n581) );
  XNOR2_X1 U612 ( .A(n576), .B(n575), .ZN(n765) );
  NAND2_X1 U613 ( .A1(G234), .A2(n783), .ZN(n497) );
  INV_X1 U614 ( .A(G140), .ZN(n498) );
  NAND2_X1 U615 ( .A1(n498), .A2(G137), .ZN(n501) );
  INV_X1 U616 ( .A(G137), .ZN(n499) );
  NAND2_X1 U617 ( .A1(n499), .A2(G140), .ZN(n500) );
  NAND2_X1 U618 ( .A1(n501), .A2(n500), .ZN(n503) );
  INV_X1 U619 ( .A(n573), .ZN(n504) );
  XOR2_X1 U620 ( .A(n506), .B(KEYINPUT23), .Z(n507) );
  INV_X1 U621 ( .A(KEYINPUT15), .ZN(n508) );
  XNOR2_X1 U622 ( .A(n508), .B(G902), .ZN(n658) );
  INV_X1 U623 ( .A(n658), .ZN(n509) );
  NAND2_X1 U624 ( .A1(n509), .A2(G234), .ZN(n510) );
  XNOR2_X1 U625 ( .A(n510), .B(KEYINPUT20), .ZN(n550) );
  NAND2_X1 U626 ( .A1(G217), .A2(n550), .ZN(n511) );
  XNOR2_X2 U627 ( .A(G128), .B(KEYINPUT71), .ZN(n514) );
  XNOR2_X1 U628 ( .A(n347), .B(n515), .ZN(n525) );
  XNOR2_X1 U629 ( .A(n516), .B(KEYINPUT16), .ZN(n519) );
  XNOR2_X1 U630 ( .A(KEYINPUT3), .B(G113), .ZN(n518) );
  XNOR2_X1 U631 ( .A(n518), .B(n517), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n519), .B(n564), .ZN(n524) );
  XNOR2_X1 U633 ( .A(n522), .B(G104), .ZN(n572) );
  XNOR2_X1 U634 ( .A(n549), .B(n572), .ZN(n523) );
  XNOR2_X1 U635 ( .A(n526), .B(KEYINPUT68), .ZN(n530) );
  INV_X1 U636 ( .A(G210), .ZN(n527) );
  NOR2_X1 U637 ( .A1(n530), .A2(n527), .ZN(n528) );
  INV_X1 U638 ( .A(G214), .ZN(n529) );
  INV_X1 U639 ( .A(KEYINPUT19), .ZN(n531) );
  XNOR2_X1 U640 ( .A(n532), .B(KEYINPUT14), .ZN(n535) );
  NAND2_X1 U641 ( .A1(G902), .A2(n535), .ZN(n533) );
  XOR2_X1 U642 ( .A(KEYINPUT84), .B(n533), .Z(n534) );
  NAND2_X1 U643 ( .A1(G953), .A2(n534), .ZN(n607) );
  NOR2_X1 U644 ( .A1(n607), .A2(G898), .ZN(n536) );
  NAND2_X1 U645 ( .A1(G952), .A2(n535), .ZN(n754) );
  NOR2_X1 U646 ( .A1(n754), .A2(G953), .ZN(n610) );
  XOR2_X1 U647 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n538) );
  XNOR2_X1 U648 ( .A(G122), .B(KEYINPUT11), .ZN(n537) );
  XOR2_X1 U649 ( .A(KEYINPUT90), .B(G104), .Z(n540) );
  NAND2_X1 U650 ( .A1(G214), .A2(n561), .ZN(n543) );
  XOR2_X1 U651 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n545) );
  XNOR2_X1 U652 ( .A(G134), .B(KEYINPUT91), .ZN(n544) );
  NOR2_X1 U653 ( .A1(n597), .A2(n595), .ZN(n617) );
  XOR2_X1 U654 ( .A(KEYINPUT21), .B(KEYINPUT86), .Z(n552) );
  NAND2_X1 U655 ( .A1(n550), .A2(G221), .ZN(n551) );
  XNOR2_X1 U656 ( .A(n552), .B(n551), .ZN(n722) );
  NAND2_X1 U657 ( .A1(n617), .A2(n722), .ZN(n553) );
  XNOR2_X1 U658 ( .A(n553), .B(KEYINPUT95), .ZN(n554) );
  NAND2_X1 U659 ( .A1(n593), .A2(n554), .ZN(n555) );
  XOR2_X1 U660 ( .A(n560), .B(n559), .Z(n563) );
  NAND2_X1 U661 ( .A1(n561), .A2(G210), .ZN(n562) );
  XNOR2_X1 U662 ( .A(n563), .B(n562), .ZN(n565) );
  XNOR2_X1 U663 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X2 U664 ( .A(n576), .B(n566), .ZN(n665) );
  INV_X1 U665 ( .A(G472), .ZN(n567) );
  INV_X1 U666 ( .A(KEYINPUT6), .ZN(n568) );
  XNOR2_X1 U667 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U668 ( .A(n574), .B(n573), .ZN(n575) );
  NOR2_X1 U669 ( .A1(n630), .A2(n448), .ZN(n578) );
  INV_X1 U670 ( .A(KEYINPUT32), .ZN(n579) );
  NOR2_X2 U671 ( .A1(n727), .A2(n726), .ZN(n588) );
  NAND2_X1 U672 ( .A1(n588), .A2(n630), .ZN(n582) );
  INV_X1 U673 ( .A(n593), .ZN(n589) );
  XNOR2_X1 U674 ( .A(n583), .B(KEYINPUT34), .ZN(n584) );
  AND2_X1 U675 ( .A1(n597), .A2(n595), .ZN(n640) );
  NAND2_X1 U676 ( .A1(n584), .A2(n640), .ZN(n585) );
  NAND2_X1 U677 ( .A1(n448), .A2(n592), .ZN(n586) );
  XOR2_X1 U678 ( .A(KEYINPUT87), .B(KEYINPUT31), .Z(n590) );
  AND2_X1 U679 ( .A1(n592), .A2(n612), .ZN(n594) );
  AND2_X1 U680 ( .A1(n593), .A2(n594), .ZN(n702) );
  NOR2_X1 U681 ( .A1(n596), .A2(n597), .ZN(n713) );
  INV_X1 U682 ( .A(n713), .ZN(n656) );
  NAND2_X1 U683 ( .A1(n656), .A2(n627), .ZN(n644) );
  INV_X1 U684 ( .A(n644), .ZN(n743) );
  NAND2_X1 U685 ( .A1(n448), .A2(n345), .ZN(n598) );
  OR2_X1 U686 ( .A1(n598), .A2(n630), .ZN(n599) );
  OR2_X1 U687 ( .A1(n600), .A2(n599), .ZN(n699) );
  NAND2_X1 U688 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U689 ( .A1(n661), .A2(n658), .ZN(n605) );
  INV_X1 U690 ( .A(KEYINPUT38), .ZN(n606) );
  XNOR2_X1 U691 ( .A(n655), .B(n606), .ZN(n738) );
  XNOR2_X1 U692 ( .A(KEYINPUT98), .B(n607), .ZN(n608) );
  NOR2_X1 U693 ( .A1(G900), .A2(n608), .ZN(n609) );
  NOR2_X1 U694 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U695 ( .A1(n613), .A2(n637), .ZN(n615) );
  INV_X1 U696 ( .A(KEYINPUT39), .ZN(n614) );
  XNOR2_X1 U697 ( .A(n616), .B(KEYINPUT40), .ZN(n792) );
  NAND2_X1 U698 ( .A1(n738), .A2(n737), .ZN(n742) );
  INV_X1 U699 ( .A(n617), .ZN(n741) );
  NOR2_X1 U700 ( .A1(n742), .A2(n741), .ZN(n618) );
  XNOR2_X1 U701 ( .A(n618), .B(KEYINPUT41), .ZN(n735) );
  AND2_X1 U702 ( .A1(n722), .A2(n344), .ZN(n619) );
  AND2_X2 U703 ( .A1(n620), .A2(n619), .ZN(n628) );
  INV_X1 U704 ( .A(KEYINPUT28), .ZN(n621) );
  NAND2_X1 U705 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n624), .A2(n364), .ZN(n625) );
  NOR2_X1 U707 ( .A1(n735), .A2(n643), .ZN(n626) );
  XNOR2_X1 U708 ( .A(n626), .B(KEYINPUT42), .ZN(n793) );
  NAND2_X1 U709 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U710 ( .A(n631), .B(KEYINPUT99), .ZN(n632) );
  INV_X1 U711 ( .A(n655), .ZN(n633) );
  XNOR2_X1 U712 ( .A(n634), .B(KEYINPUT36), .ZN(n635) );
  INV_X1 U713 ( .A(n448), .ZN(n654) );
  AND2_X1 U714 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n638), .A2(n655), .ZN(n639) );
  XNOR2_X1 U716 ( .A(n639), .B(KEYINPUT103), .ZN(n641) );
  NAND2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n709) );
  NAND2_X1 U718 ( .A1(n647), .A2(n644), .ZN(n645) );
  NAND2_X1 U719 ( .A1(n645), .A2(KEYINPUT74), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n646), .B(KEYINPUT47), .ZN(n651) );
  INV_X1 U721 ( .A(KEYINPUT74), .ZN(n649) );
  NAND2_X1 U722 ( .A1(n647), .A2(n743), .ZN(n648) );
  NAND2_X1 U723 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U724 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n720) );
  INV_X1 U726 ( .A(KEYINPUT2), .ZN(n755) );
  NOR2_X1 U727 ( .A1(n756), .A2(n755), .ZN(n759) );
  INV_X1 U728 ( .A(n759), .ZN(n662) );
  NAND2_X1 U729 ( .A1(n771), .A2(G472), .ZN(n666) );
  XOR2_X1 U730 ( .A(KEYINPUT62), .B(KEYINPUT105), .Z(n664) );
  XNOR2_X1 U731 ( .A(n666), .B(n359), .ZN(n668) );
  NOR2_X1 U732 ( .A1(n783), .A2(G952), .ZN(n667) );
  XOR2_X1 U733 ( .A(KEYINPUT80), .B(KEYINPUT63), .Z(n669) );
  XNOR2_X1 U734 ( .A(n496), .B(n669), .ZN(G57) );
  NAND2_X1 U735 ( .A1(n771), .A2(G217), .ZN(n671) );
  XNOR2_X1 U736 ( .A(n671), .B(n670), .ZN(n672) );
  NOR2_X2 U737 ( .A1(n672), .A2(n778), .ZN(n673) );
  XNOR2_X1 U738 ( .A(n673), .B(KEYINPUT124), .ZN(G66) );
  NAND2_X1 U739 ( .A1(n771), .A2(G210), .ZN(n678) );
  XNOR2_X1 U740 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n674) );
  XNOR2_X1 U741 ( .A(n674), .B(KEYINPUT117), .ZN(n675) );
  XNOR2_X1 U742 ( .A(n678), .B(n677), .ZN(n679) );
  NOR2_X2 U743 ( .A1(n679), .A2(n778), .ZN(n681) );
  XNOR2_X1 U744 ( .A(KEYINPUT56), .B(KEYINPUT118), .ZN(n680) );
  XNOR2_X1 U745 ( .A(n681), .B(n680), .ZN(G51) );
  XNOR2_X1 U746 ( .A(n683), .B(n682), .ZN(G21) );
  XOR2_X1 U747 ( .A(G110), .B(n684), .Z(G12) );
  NAND2_X1 U748 ( .A1(n661), .A2(n783), .ZN(n685) );
  XOR2_X1 U749 ( .A(KEYINPUT125), .B(n685), .Z(n689) );
  NAND2_X1 U750 ( .A1(G953), .A2(G224), .ZN(n686) );
  XNOR2_X1 U751 ( .A(KEYINPUT61), .B(n686), .ZN(n687) );
  NAND2_X1 U752 ( .A1(n687), .A2(G898), .ZN(n688) );
  NAND2_X1 U753 ( .A1(n689), .A2(n688), .ZN(n691) );
  NOR2_X1 U754 ( .A1(G898), .A2(n783), .ZN(n690) );
  XNOR2_X1 U755 ( .A(n691), .B(n362), .ZN(G69) );
  NAND2_X1 U756 ( .A1(n771), .A2(G475), .ZN(n695) );
  XNOR2_X1 U757 ( .A(KEYINPUT79), .B(KEYINPUT120), .ZN(n692) );
  XNOR2_X1 U758 ( .A(n692), .B(KEYINPUT59), .ZN(n693) );
  XNOR2_X1 U759 ( .A(n695), .B(n360), .ZN(n697) );
  INV_X1 U760 ( .A(n778), .ZN(n696) );
  XOR2_X1 U761 ( .A(KEYINPUT121), .B(KEYINPUT60), .Z(n698) );
  XNOR2_X1 U762 ( .A(n495), .B(n698), .ZN(G60) );
  XNOR2_X1 U763 ( .A(G101), .B(KEYINPUT106), .ZN(n700) );
  XNOR2_X1 U764 ( .A(n700), .B(n699), .ZN(G3) );
  NAND2_X1 U765 ( .A1(n702), .A2(n711), .ZN(n701) );
  XNOR2_X1 U766 ( .A(n701), .B(G104), .ZN(G6) );
  XOR2_X1 U767 ( .A(KEYINPUT107), .B(KEYINPUT27), .Z(n704) );
  NAND2_X1 U768 ( .A1(n702), .A2(n713), .ZN(n703) );
  XNOR2_X1 U769 ( .A(n704), .B(n703), .ZN(n706) );
  XOR2_X1 U770 ( .A(G107), .B(KEYINPUT26), .Z(n705) );
  XNOR2_X1 U771 ( .A(n706), .B(n705), .ZN(G9) );
  XOR2_X1 U772 ( .A(G128), .B(KEYINPUT29), .Z(n708) );
  NAND2_X1 U773 ( .A1(n647), .A2(n713), .ZN(n707) );
  XNOR2_X1 U774 ( .A(n708), .B(n707), .ZN(G30) );
  XNOR2_X1 U775 ( .A(G143), .B(n709), .ZN(G45) );
  NAND2_X1 U776 ( .A1(n647), .A2(n711), .ZN(n710) );
  XNOR2_X1 U777 ( .A(n710), .B(G146), .ZN(G48) );
  NAND2_X1 U778 ( .A1(n714), .A2(n711), .ZN(n712) );
  XNOR2_X1 U779 ( .A(n712), .B(G113), .ZN(G15) );
  XOR2_X1 U780 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n716) );
  NAND2_X1 U781 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U782 ( .A(n716), .B(n715), .ZN(n717) );
  XNOR2_X1 U783 ( .A(G116), .B(n717), .ZN(G18) );
  XOR2_X1 U784 ( .A(KEYINPUT110), .B(KEYINPUT37), .Z(n718) );
  XNOR2_X1 U785 ( .A(G125), .B(n719), .ZN(G27) );
  XOR2_X1 U786 ( .A(G134), .B(n720), .Z(G36) );
  NOR2_X1 U787 ( .A1(n735), .A2(n420), .ZN(n721) );
  NOR2_X1 U788 ( .A1(G953), .A2(n721), .ZN(n763) );
  NOR2_X1 U789 ( .A1(n722), .A2(n345), .ZN(n724) );
  XNOR2_X1 U790 ( .A(KEYINPUT49), .B(KEYINPUT111), .ZN(n723) );
  XNOR2_X1 U791 ( .A(n724), .B(n723), .ZN(n725) );
  XNOR2_X1 U792 ( .A(n357), .B(KEYINPUT112), .ZN(n730) );
  NAND2_X1 U793 ( .A1(n448), .A2(n726), .ZN(n728) );
  XNOR2_X1 U794 ( .A(KEYINPUT50), .B(n728), .ZN(n729) );
  NAND2_X1 U795 ( .A1(n730), .A2(n729), .ZN(n732) );
  NAND2_X1 U796 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U797 ( .A(KEYINPUT51), .B(n733), .ZN(n734) );
  NOR2_X1 U798 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U799 ( .A(KEYINPUT113), .B(n736), .Z(n750) );
  NOR2_X1 U800 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U801 ( .A(n739), .B(KEYINPUT114), .ZN(n740) );
  NOR2_X1 U802 ( .A1(n741), .A2(n740), .ZN(n746) );
  NOR2_X1 U803 ( .A1(n743), .A2(n742), .ZN(n744) );
  XOR2_X1 U804 ( .A(KEYINPUT115), .B(n744), .Z(n745) );
  NOR2_X1 U805 ( .A1(n746), .A2(n745), .ZN(n748) );
  NOR2_X1 U806 ( .A1(n748), .A2(n420), .ZN(n749) );
  NOR2_X1 U807 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U808 ( .A(n751), .B(KEYINPUT52), .ZN(n752) );
  XNOR2_X1 U809 ( .A(KEYINPUT116), .B(n752), .ZN(n753) );
  NOR2_X1 U810 ( .A1(n754), .A2(n753), .ZN(n761) );
  NAND2_X1 U811 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U812 ( .A(KEYINPUT73), .B(n757), .ZN(n758) );
  NOR2_X1 U813 ( .A1(n759), .A2(n758), .ZN(n760) );
  NOR2_X1 U814 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U815 ( .A1(n763), .A2(n762), .ZN(n764) );
  XOR2_X1 U816 ( .A(KEYINPUT53), .B(n764), .Z(G75) );
  XOR2_X1 U817 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n767) );
  XNOR2_X1 U818 ( .A(n765), .B(KEYINPUT119), .ZN(n766) );
  XNOR2_X1 U819 ( .A(n767), .B(n766), .ZN(n769) );
  NAND2_X1 U820 ( .A1(n771), .A2(G469), .ZN(n768) );
  XOR2_X1 U821 ( .A(n769), .B(n768), .Z(n770) );
  NOR2_X1 U822 ( .A1(n778), .A2(n770), .ZN(G54) );
  BUF_X1 U823 ( .A(n771), .Z(n772) );
  NAND2_X1 U824 ( .A1(n772), .A2(G478), .ZN(n776) );
  XOR2_X1 U825 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n773) );
  NOR2_X1 U826 ( .A1(n778), .A2(n777), .ZN(G63) );
  XOR2_X1 U827 ( .A(n779), .B(KEYINPUT126), .Z(n780) );
  XOR2_X1 U828 ( .A(n781), .B(n780), .Z(n785) );
  XOR2_X1 U829 ( .A(n785), .B(n346), .Z(n784) );
  NAND2_X1 U830 ( .A1(n784), .A2(n783), .ZN(n789) );
  XNOR2_X1 U831 ( .A(G227), .B(n785), .ZN(n786) );
  NAND2_X1 U832 ( .A1(n786), .A2(G900), .ZN(n787) );
  NAND2_X1 U833 ( .A1(G953), .A2(n787), .ZN(n788) );
  NAND2_X1 U834 ( .A1(n789), .A2(n788), .ZN(G72) );
  BUF_X1 U835 ( .A(n790), .Z(n791) );
  XOR2_X1 U836 ( .A(G122), .B(n791), .Z(G24) );
  XOR2_X1 U837 ( .A(n792), .B(G131), .Z(G33) );
  XOR2_X1 U838 ( .A(G137), .B(n793), .Z(G39) );
endmodule

