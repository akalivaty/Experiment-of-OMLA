//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1237,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n203), .A2(G50), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(KEYINPUT64), .ZN(new_n216));
  INV_X1    g0016(.A(KEYINPUT64), .ZN(new_n217));
  NAND3_X1  g0017(.A1(new_n217), .A2(G1), .A3(G13), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n214), .A2(G20), .A3(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n202), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n209), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n212), .B(new_n220), .C1(KEYINPUT1), .C2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT1), .B2(new_n229), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XOR2_X1   g0040(.A(G107), .B(G116), .Z(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT65), .ZN(new_n243));
  INV_X1    g0043(.A(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G68), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n202), .A2(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n243), .B(new_n249), .ZN(G351));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  AOI22_X1  g0051(.A1(new_n251), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G20), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G77), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n252), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n216), .A2(new_n218), .A3(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  OR2_X1    g0060(.A1(new_n260), .A2(KEYINPUT11), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n202), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n264), .B(KEYINPUT12), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n260), .A2(KEYINPUT11), .ZN(new_n266));
  NAND4_X1  g0066(.A1(new_n216), .A2(new_n218), .A3(new_n262), .A4(new_n258), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n206), .A2(G20), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(G68), .A3(new_n269), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n261), .A2(new_n265), .A3(new_n266), .A4(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT66), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n215), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(KEYINPUT66), .A2(G33), .A3(G41), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n272), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  INV_X1    g0078(.A(G45), .ZN(new_n279));
  AOI21_X1  g0079(.A(G1), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n275), .A2(new_n276), .ZN(new_n282));
  INV_X1    g0082(.A(new_n280), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n281), .B1(new_n284), .B2(new_n222), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT70), .ZN(new_n287));
  INV_X1    g0087(.A(G1698), .ZN(new_n288));
  AND2_X1   g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NOR2_X1   g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  OAI211_X1 g0090(.A(G226), .B(new_n288), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT69), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT3), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n253), .ZN(new_n295));
  NAND2_X1  g0095(.A1(KEYINPUT3), .A2(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n297), .A2(KEYINPUT69), .A3(G226), .A4(new_n288), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(G232), .B(G1698), .C1(new_n289), .C2(new_n290), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G97), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n219), .A2(new_n274), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n287), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n302), .B1(new_n293), .B2(new_n298), .ZN(new_n308));
  NOR3_X1   g0108(.A1(new_n308), .A2(KEYINPUT70), .A3(new_n305), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n286), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT13), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n304), .A2(new_n287), .A3(new_n306), .ZN(new_n312));
  OAI21_X1  g0112(.A(KEYINPUT70), .B1(new_n308), .B2(new_n305), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT13), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(new_n315), .A3(new_n286), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n311), .A2(G179), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT71), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT71), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n311), .A2(new_n319), .A3(G179), .A4(new_n316), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n315), .B1(new_n314), .B2(new_n286), .ZN(new_n322));
  AOI211_X1 g0122(.A(KEYINPUT13), .B(new_n285), .C1(new_n312), .C2(new_n313), .ZN(new_n323));
  OAI21_X1  g0123(.A(G169), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT14), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n311), .A2(new_n316), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT14), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n327), .A3(G169), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NOR3_X1   g0129(.A1(new_n321), .A2(new_n329), .A3(KEYINPUT72), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT72), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n327), .B1(new_n326), .B2(G169), .ZN(new_n332));
  INV_X1    g0132(.A(G169), .ZN(new_n333));
  AOI211_X1 g0133(.A(KEYINPUT14), .B(new_n333), .C1(new_n311), .C2(new_n316), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n318), .A2(new_n320), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n331), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n271), .B1(new_n330), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n326), .A2(G200), .ZN(new_n340));
  INV_X1    g0140(.A(new_n271), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n311), .A2(G190), .A3(new_n316), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n269), .A2(G50), .ZN(new_n346));
  OAI22_X1  g0146(.A1(new_n267), .A2(new_n346), .B1(G50), .B2(new_n262), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n347), .B(KEYINPUT67), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n251), .A2(G150), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT8), .B(G58), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(new_n255), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n203), .A2(G50), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n352), .A2(new_n207), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n259), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n348), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT9), .ZN(new_n356));
  INV_X1    g0156(.A(new_n284), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G226), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n288), .B1(new_n295), .B2(new_n296), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G223), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n256), .B2(new_n297), .ZN(new_n361));
  AOI21_X1  g0161(.A(G1698), .B1(new_n295), .B2(new_n296), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n361), .B1(G222), .B2(new_n362), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n281), .B(new_n358), .C1(new_n363), .C2(new_n305), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G200), .ZN(new_n365));
  INV_X1    g0165(.A(G190), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n356), .B(new_n365), .C1(new_n366), .C2(new_n364), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n367), .B(KEYINPUT10), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n364), .A2(new_n333), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n369), .B(new_n355), .C1(G179), .C2(new_n364), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(G58), .A2(G68), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n203), .A2(new_n372), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(G20), .B1(G159), .B2(new_n251), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n295), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n296), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT73), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n289), .A2(new_n290), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT73), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(KEYINPUT7), .A4(new_n207), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n295), .A2(new_n207), .A3(new_n296), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT7), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n376), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  AND3_X1   g0183(.A1(new_n383), .A2(KEYINPUT74), .A3(G68), .ZN(new_n384));
  AOI21_X1  g0184(.A(KEYINPUT74), .B1(new_n383), .B2(G68), .ZN(new_n385));
  OAI211_X1 g0185(.A(KEYINPUT16), .B(new_n374), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n259), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n382), .A2(new_n375), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n374), .B1(new_n389), .B2(new_n202), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT16), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n387), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n350), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(new_n269), .ZN(new_n395));
  OAI22_X1  g0195(.A1(new_n395), .A2(new_n267), .B1(new_n262), .B2(new_n394), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT76), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n282), .A2(G232), .A3(new_n283), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n281), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n297), .A2(G226), .A3(G1698), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G87), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT75), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n297), .A2(new_n405), .A3(G223), .A4(new_n288), .ZN(new_n406));
  OAI211_X1 g0206(.A(G223), .B(new_n288), .C1(new_n289), .C2(new_n290), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT75), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n404), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n399), .B(new_n401), .C1(new_n409), .C2(new_n305), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n406), .ZN(new_n411));
  AOI22_X1  g0211(.A1(new_n359), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n305), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n281), .A2(new_n400), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT76), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(G179), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n413), .A2(new_n414), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n416), .A2(new_n333), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n398), .A2(new_n419), .ZN(new_n420));
  XOR2_X1   g0220(.A(new_n420), .B(KEYINPUT18), .Z(new_n421));
  INV_X1    g0221(.A(G200), .ZN(new_n422));
  AOI22_X1  g0222(.A1(new_n416), .A2(new_n422), .B1(new_n366), .B2(new_n418), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n398), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT17), .ZN(new_n425));
  XNOR2_X1  g0225(.A(new_n424), .B(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n421), .A2(new_n426), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n394), .A2(new_n251), .B1(G20), .B2(G77), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT15), .B(G87), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n428), .A2(KEYINPUT68), .B1(new_n254), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(KEYINPUT68), .B2(new_n428), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n259), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n269), .A2(G77), .ZN(new_n434));
  OAI221_X1 g0234(.A(new_n433), .B1(G77), .B2(new_n262), .C1(new_n267), .C2(new_n434), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n359), .A2(G238), .B1(new_n377), .B2(G107), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n297), .A2(G232), .A3(new_n288), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n306), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n357), .A2(G244), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n439), .A2(new_n281), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n435), .B1(G190), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n422), .B2(new_n442), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n417), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n435), .B(new_n445), .C1(G169), .C2(new_n442), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n371), .A2(new_n427), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n345), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G283), .ZN(new_n451));
  XNOR2_X1  g0251(.A(new_n451), .B(KEYINPUT79), .ZN(new_n452));
  OAI211_X1 g0252(.A(G250), .B(G1698), .C1(new_n289), .C2(new_n290), .ZN(new_n453));
  OAI211_X1 g0253(.A(G244), .B(new_n288), .C1(new_n289), .C2(new_n290), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT4), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n452), .B(new_n453), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(KEYINPUT4), .B1(new_n362), .B2(G244), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n306), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n206), .B(G45), .C1(new_n278), .C2(KEYINPUT5), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n278), .A2(KEYINPUT5), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT80), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT80), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n462), .A2(new_n278), .A3(KEYINPUT5), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n459), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n277), .A2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n459), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n466), .A2(new_n460), .B1(new_n275), .B2(new_n276), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G257), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n458), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n333), .ZN(new_n470));
  XOR2_X1   g0270(.A(G97), .B(G107), .Z(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT77), .B(KEYINPUT6), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n472), .A2(KEYINPUT78), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n472), .A2(G97), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n471), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n472), .A2(KEYINPUT78), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n475), .A2(G20), .A3(new_n478), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n388), .A2(G107), .B1(G77), .B2(new_n251), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n387), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n262), .A2(G97), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n267), .B1(new_n206), .B2(G33), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n482), .B1(new_n483), .B2(G97), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  OAI221_X1 g0285(.A(new_n470), .B1(G179), .B2(new_n469), .C1(new_n481), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n469), .A2(G200), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT81), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT81), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n469), .A2(new_n489), .A3(G200), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n458), .A2(G190), .A3(new_n465), .A4(new_n468), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n479), .A2(new_n480), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n484), .B(new_n492), .C1(new_n493), .C2(new_n387), .ZN(new_n494));
  OAI211_X1 g0294(.A(KEYINPUT82), .B(new_n486), .C1(new_n491), .C2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT82), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n494), .B1(new_n490), .B2(new_n488), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n470), .B1(new_n481), .B2(new_n485), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n469), .A2(G179), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n496), .B1(new_n497), .B2(new_n500), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n467), .A2(G270), .B1(new_n277), .B2(new_n464), .ZN(new_n502));
  OAI211_X1 g0302(.A(G264), .B(G1698), .C1(new_n289), .C2(new_n290), .ZN(new_n503));
  OAI211_X1 g0303(.A(G257), .B(new_n288), .C1(new_n289), .C2(new_n290), .ZN(new_n504));
  INV_X1    g0304(.A(G303), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n503), .B(new_n504), .C1(new_n505), .C2(new_n297), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n306), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n502), .A2(KEYINPUT85), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT85), .B1(new_n502), .B2(new_n507), .ZN(new_n509));
  OAI21_X1  g0309(.A(G190), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT85), .ZN(new_n511));
  INV_X1    g0311(.A(new_n507), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n466), .A2(new_n460), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(G270), .A3(new_n282), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n465), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n511), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n502), .A2(KEYINPUT85), .A3(new_n507), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n516), .A2(G200), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(G97), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n207), .B1(new_n519), .B2(G33), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n452), .A2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(G116), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G20), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n522), .A2(KEYINPUT20), .A3(new_n259), .A4(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT20), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n259), .A2(new_n524), .ZN(new_n527));
  OR2_X1    g0327(.A1(new_n451), .A2(KEYINPUT79), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n451), .A2(KEYINPUT79), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n520), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n526), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n262), .A2(G116), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n533), .B1(new_n483), .B2(G116), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n510), .A2(new_n518), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT21), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n516), .A2(new_n517), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n535), .A2(G169), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n508), .A2(new_n509), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n333), .B1(new_n532), .B2(new_n534), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n542), .A2(KEYINPUT21), .A3(new_n543), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n512), .A2(new_n515), .A3(new_n417), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n535), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n537), .A2(new_n541), .A3(new_n544), .A4(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n362), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n297), .A2(G257), .A3(G1698), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n306), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n467), .A2(G264), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n551), .A2(new_n465), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n333), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n465), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n305), .B1(new_n548), .B2(new_n549), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n417), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT86), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n207), .B2(G107), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT23), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT23), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n559), .B(new_n562), .C1(new_n207), .C2(G107), .ZN(new_n563));
  AOI22_X1  g0363(.A1(new_n561), .A2(new_n563), .B1(G116), .B2(new_n254), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n207), .B(G87), .C1(new_n289), .C2(new_n290), .ZN(new_n565));
  AND2_X1   g0365(.A1(new_n565), .A2(KEYINPUT22), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n565), .A2(KEYINPUT22), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT24), .ZN(new_n569));
  XNOR2_X1  g0369(.A(new_n565), .B(KEYINPUT22), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT24), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n570), .A2(new_n571), .A3(new_n564), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n387), .B1(new_n569), .B2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT25), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n262), .B2(G107), .ZN(new_n575));
  INV_X1    g0375(.A(G107), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n263), .A2(KEYINPUT25), .A3(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n483), .A2(G107), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n554), .B(new_n558), .C1(new_n573), .C2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n568), .A2(KEYINPUT24), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n571), .B1(new_n570), .B2(new_n564), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n259), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n551), .A2(G190), .A3(new_n465), .A4(new_n552), .ZN(new_n584));
  OAI21_X1  g0384(.A(G200), .B1(new_n555), .B2(new_n556), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n583), .A2(new_n578), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n362), .A2(G238), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n359), .A2(G244), .ZN(new_n588));
  NAND2_X1  g0388(.A1(G33), .A2(G116), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n306), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT83), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n279), .A2(G1), .A3(G274), .ZN(new_n593));
  AOI21_X1  g0393(.A(G250), .B1(new_n206), .B2(G45), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n592), .B1(new_n282), .B2(new_n595), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n282), .A2(new_n592), .A3(new_n595), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n591), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(G200), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n297), .A2(new_n207), .A3(G68), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT84), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT84), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n297), .A2(new_n602), .A3(new_n207), .A4(G68), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT19), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n254), .A2(new_n604), .A3(G97), .ZN(new_n605));
  NOR2_X1   g0405(.A1(G97), .A2(G107), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n606), .A2(new_n223), .B1(new_n301), .B2(new_n207), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n605), .B1(new_n607), .B2(new_n604), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n601), .A2(new_n603), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n259), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n429), .A2(new_n263), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n483), .A2(G87), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n591), .B(G190), .C1(new_n596), .C2(new_n597), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n599), .A2(new_n612), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n598), .A2(new_n333), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n483), .A2(new_n430), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n610), .A2(new_n611), .A3(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n591), .B(new_n417), .C1(new_n596), .C2(new_n597), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n616), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n580), .A2(new_n586), .A3(new_n615), .A4(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n547), .A2(new_n621), .ZN(new_n622));
  AND4_X1   g0422(.A1(new_n450), .A2(new_n495), .A3(new_n501), .A4(new_n622), .ZN(G372));
  OAI21_X1  g0423(.A(new_n338), .B1(new_n344), .B2(new_n446), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n624), .A2(new_n426), .ZN(new_n625));
  INV_X1    g0425(.A(new_n421), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n368), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n627), .A2(new_n370), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n500), .A2(KEYINPUT88), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n615), .A2(new_n620), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT88), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n486), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n633), .A2(KEYINPUT26), .ZN(new_n634));
  INV_X1    g0434(.A(new_n620), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n630), .A2(new_n500), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n635), .B1(new_n636), .B2(KEYINPUT26), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n580), .B(KEYINPUT87), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n541), .A2(new_n544), .A3(new_n546), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n497), .A2(new_n500), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n641), .A2(new_n586), .A3(new_n630), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n634), .B(new_n637), .C1(new_n640), .C2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n628), .B1(new_n449), .B2(new_n644), .ZN(G369));
  NAND3_X1  g0445(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n646), .A2(KEYINPUT27), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n647), .B(KEYINPUT89), .ZN(new_n648));
  INV_X1    g0448(.A(G213), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n646), .B2(KEYINPUT27), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(G343), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n536), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n639), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(new_n547), .B2(new_n655), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(G330), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(KEYINPUT90), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  AND2_X1   g0460(.A1(new_n580), .A2(new_n586), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n653), .B1(new_n573), .B2(new_n579), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n580), .B2(new_n654), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n638), .A2(new_n654), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n639), .A2(new_n654), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n661), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n665), .A2(new_n666), .A3(new_n668), .ZN(G399));
  INV_X1    g0469(.A(new_n210), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(G41), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n606), .A2(new_n223), .A3(new_n523), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n671), .A2(new_n672), .A3(new_n206), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(new_n214), .B2(new_n671), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT28), .Z(new_n675));
  NOR2_X1   g0475(.A1(new_n644), .A2(new_n653), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n620), .B1(new_n636), .B2(KEYINPUT26), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n677), .B1(KEYINPUT26), .B2(new_n633), .ZN(new_n678));
  INV_X1    g0478(.A(new_n580), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n639), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n678), .B1(new_n642), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n654), .ZN(new_n682));
  MUX2_X1   g0482(.A(new_n676), .B(new_n682), .S(KEYINPUT29), .Z(new_n683));
  NOR2_X1   g0483(.A1(new_n553), .A2(new_n598), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n458), .A2(new_n468), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(new_n685), .A3(new_n545), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT30), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n684), .A2(KEYINPUT30), .A3(new_n685), .A4(new_n545), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n557), .A2(G179), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n542), .A2(new_n690), .A3(new_n469), .A4(new_n598), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n653), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n622), .A2(new_n501), .A3(new_n495), .A4(new_n654), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n694), .B1(new_n695), .B2(KEYINPUT31), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT31), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(G330), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n683), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n675), .B1(new_n701), .B2(G1), .ZN(G364));
  INV_X1    g0502(.A(new_n671), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n207), .A2(G13), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n206), .B1(new_n704), .B2(G45), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n703), .A2(KEYINPUT91), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT91), .ZN(new_n707));
  INV_X1    g0507(.A(new_n705), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n707), .B1(new_n671), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n659), .B(new_n710), .C1(G330), .C2(new_n657), .ZN(new_n711));
  INV_X1    g0511(.A(new_n710), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n670), .A2(new_n297), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n213), .A2(G45), .ZN(new_n715));
  OR3_X1    g0515(.A1(new_n714), .A2(KEYINPUT93), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT93), .B1(new_n714), .B2(new_n715), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n716), .B(new_n717), .C1(new_n279), .C2(new_n249), .ZN(new_n718));
  INV_X1    g0518(.A(G355), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(KEYINPUT92), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n670), .A2(new_n377), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT92), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(G355), .ZN(new_n723));
  OAI221_X1 g0523(.A(new_n718), .B1(G116), .B2(new_n210), .C1(new_n720), .C2(new_n723), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n724), .A2(KEYINPUT94), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n219), .B1(new_n207), .B2(G169), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(G13), .A2(G33), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G20), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(new_n724), .B2(KEYINPUT94), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n712), .B1(new_n725), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n207), .A2(G179), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(new_n366), .A3(G200), .ZN(new_n735));
  INV_X1    g0535(.A(G283), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n734), .A2(new_n366), .A3(new_n422), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI211_X1 g0539(.A(new_n297), .B(new_n737), .C1(G329), .C2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G294), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n366), .A2(G179), .A3(G200), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(new_n207), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n734), .A2(G190), .A3(G200), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT98), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OAI221_X1 g0546(.A(new_n740), .B1(new_n741), .B2(new_n743), .C1(new_n505), .C2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT96), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(new_n366), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT95), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(new_n207), .B2(new_n417), .ZN(new_n752));
  NAND3_X1  g0552(.A1(KEYINPUT95), .A2(G20), .A3(G179), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n752), .A2(new_n422), .A3(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n366), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n750), .A2(G326), .B1(new_n755), .B2(G322), .ZN(new_n756));
  INV_X1    g0556(.A(G311), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n754), .A2(G190), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n749), .A2(G190), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  XOR2_X1   g0561(.A(KEYINPUT33), .B(G317), .Z(new_n762));
  OAI221_X1 g0562(.A(new_n756), .B1(new_n757), .B2(new_n759), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  AOI22_X1  g0563(.A1(new_n760), .A2(G68), .B1(new_n755), .B2(G58), .ZN(new_n764));
  INV_X1    g0564(.A(new_n750), .ZN(new_n765));
  OAI221_X1 g0565(.A(new_n764), .B1(new_n244), .B2(new_n765), .C1(new_n256), .C2(new_n759), .ZN(new_n766));
  XOR2_X1   g0566(.A(KEYINPUT97), .B(G159), .Z(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n738), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT32), .ZN(new_n769));
  INV_X1    g0569(.A(new_n743), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G97), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n735), .A2(new_n576), .ZN(new_n772));
  INV_X1    g0572(.A(new_n744), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n772), .B1(G87), .B2(new_n773), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n769), .A2(new_n297), .A3(new_n771), .A4(new_n774), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n747), .A2(new_n763), .B1(new_n766), .B2(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT99), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n733), .B1(new_n777), .B2(new_n727), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n730), .B(KEYINPUT100), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n778), .B1(new_n657), .B2(new_n779), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n711), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(G396));
  NOR2_X1   g0582(.A1(new_n727), .A2(new_n728), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n712), .B1(G77), .B2(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT101), .ZN(new_n786));
  INV_X1    g0586(.A(new_n767), .ZN(new_n787));
  AOI22_X1  g0587(.A1(G143), .A2(new_n755), .B1(new_n758), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G137), .ZN(new_n789));
  INV_X1    g0589(.A(G150), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n788), .B1(new_n789), .B2(new_n765), .C1(new_n790), .C2(new_n761), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT34), .ZN(new_n792));
  INV_X1    g0592(.A(G132), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n297), .B1(new_n738), .B2(new_n793), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT103), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n735), .A2(new_n202), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(G58), .B2(new_n770), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n795), .B(new_n797), .C1(new_n244), .C2(new_n746), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n377), .B1(new_n738), .B2(new_n757), .C1(new_n223), .C2(new_n735), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G283), .A2(new_n760), .B1(new_n750), .B2(G303), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(new_n523), .B2(new_n759), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n800), .B(new_n802), .C1(G107), .C2(new_n745), .ZN(new_n803));
  INV_X1    g0603(.A(new_n755), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n771), .B1(new_n804), .B2(new_n741), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT102), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n792), .A2(new_n799), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n446), .A2(new_n653), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n435), .A2(new_n653), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n444), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n808), .B1(new_n810), .B2(new_n446), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n786), .B1(new_n726), .B2(new_n807), .C1(new_n811), .C2(new_n729), .ZN(new_n812));
  INV_X1    g0612(.A(new_n811), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n644), .B2(new_n653), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n643), .A2(new_n654), .A3(new_n811), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n712), .B1(new_n817), .B2(new_n699), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n817), .A2(new_n699), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n812), .B1(new_n819), .B2(new_n820), .ZN(G384));
  AND2_X1   g0621(.A1(new_n475), .A2(new_n478), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(KEYINPUT35), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n823), .A2(G20), .A3(G116), .A4(new_n219), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n822), .A2(KEYINPUT35), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT36), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n214), .A2(G77), .A3(new_n372), .ZN(new_n828));
  AOI211_X1 g0628(.A(new_n206), .B(G13), .C1(new_n828), .C2(new_n245), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n683), .A2(new_n450), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n628), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT112), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n338), .A2(new_n653), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT39), .ZN(new_n836));
  INV_X1    g0636(.A(new_n386), .ZN(new_n837));
  INV_X1    g0637(.A(new_n374), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n383), .A2(G68), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT74), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n383), .A2(KEYINPUT74), .A3(G68), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n838), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n259), .B1(new_n843), .B2(KEYINPUT16), .ZN(new_n844));
  INV_X1    g0644(.A(KEYINPUT105), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n837), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n374), .B1(new_n384), .B2(new_n385), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n387), .B1(new_n847), .B2(new_n391), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(KEYINPUT105), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n396), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT106), .B1(new_n850), .B2(new_n651), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n386), .B1(new_n848), .B2(KEYINPUT105), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n845), .B(new_n387), .C1(new_n847), .C2(new_n391), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n397), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n424), .B1(new_n854), .B2(new_n419), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT106), .ZN(new_n856));
  INV_X1    g0656(.A(new_n651), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n851), .A2(new_n855), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(KEYINPUT37), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n416), .A2(new_n333), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n418), .A2(new_n417), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n396), .B1(new_n386), .B2(new_n392), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT107), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n411), .A2(new_n412), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n306), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n399), .B1(new_n867), .B2(new_n401), .ZN(new_n868));
  NOR3_X1   g0668(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT76), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n422), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n418), .A2(new_n366), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT37), .B1(new_n872), .B2(new_n864), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT107), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n398), .A2(new_n419), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n865), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT108), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n398), .A2(new_n877), .A3(new_n857), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT108), .B1(new_n864), .B2(new_n651), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(KEYINPUT109), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT37), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n398), .B2(new_n423), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n874), .B1(new_n398), .B2(new_n419), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT109), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n878), .A2(new_n879), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n885), .A2(new_n886), .A3(new_n887), .A4(new_n875), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n881), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n860), .A2(new_n889), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n421), .A2(new_n426), .B1(new_n851), .B2(new_n858), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n890), .A2(KEYINPUT38), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n859), .A2(KEYINPUT37), .B1(new_n888), .B2(new_n881), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n894), .B1(new_n895), .B2(new_n891), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n836), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT110), .ZN(new_n898));
  NOR3_X1   g0698(.A1(new_n895), .A2(new_n894), .A3(new_n891), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT111), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n424), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT111), .B1(new_n398), .B2(new_n423), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(new_n420), .A3(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT37), .B1(new_n903), .B2(new_n880), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n889), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n427), .A2(new_n880), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT38), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n899), .A2(new_n907), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n897), .A2(new_n898), .B1(new_n908), .B2(new_n836), .ZN(new_n909));
  AOI21_X1  g0709(.A(KEYINPUT38), .B1(new_n890), .B2(new_n892), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT39), .B1(new_n910), .B2(new_n899), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(KEYINPUT110), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n835), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n893), .A2(new_n896), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n271), .A2(new_n653), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n338), .A2(new_n343), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT72), .B1(new_n321), .B2(new_n329), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n335), .A2(new_n331), .A3(new_n336), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n271), .B(new_n653), .C1(new_n919), .C2(new_n344), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n808), .B(KEYINPUT104), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  AOI22_X1  g0722(.A1(new_n916), .A2(new_n920), .B1(new_n815), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n914), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n626), .A2(new_n651), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n913), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n833), .B(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(KEYINPUT113), .B1(new_n693), .B2(new_n697), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT113), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n692), .A2(new_n930), .A3(KEYINPUT31), .A4(new_n653), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n811), .B1(new_n696), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n916), .B2(new_n920), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n914), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT40), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n936), .B(new_n933), .C1(new_n916), .C2(new_n920), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n905), .A2(new_n906), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n893), .B1(new_n938), .B2(KEYINPUT38), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n935), .A2(new_n936), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n696), .A2(new_n932), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n940), .A2(new_n450), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(G330), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n940), .B1(new_n450), .B2(new_n941), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n928), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n206), .B2(new_n704), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n928), .A2(new_n945), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n830), .B1(new_n947), .B2(new_n948), .ZN(G367));
  OAI221_X1 g0749(.A(new_n731), .B1(new_n210), .B2(new_n429), .C1(new_n714), .C2(new_n238), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n712), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n612), .A2(new_n613), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n653), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n630), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n635), .A2(new_n952), .A3(new_n653), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n745), .A2(KEYINPUT46), .A3(G116), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n957), .B1(new_n505), .B2(new_n804), .C1(new_n757), .C2(new_n765), .ZN(new_n958));
  AOI21_X1  g0758(.A(KEYINPUT46), .B1(new_n773), .B2(G116), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n297), .B1(new_n739), .B2(G317), .ZN(new_n960));
  OAI221_X1 g0760(.A(new_n960), .B1(new_n519), .B2(new_n735), .C1(new_n576), .C2(new_n743), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n761), .A2(new_n741), .B1(new_n759), .B2(new_n736), .ZN(new_n962));
  NOR4_X1   g0762(.A1(new_n958), .A2(new_n959), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n743), .A2(new_n202), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n377), .B(new_n964), .C1(G137), .C2(new_n739), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n750), .A2(G143), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n755), .A2(G150), .ZN(new_n967));
  INV_X1    g0767(.A(new_n735), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n773), .A2(G58), .B1(new_n968), .B2(G77), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n965), .A2(new_n966), .A3(new_n967), .A4(new_n969), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n760), .A2(new_n787), .B1(new_n758), .B2(G50), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(KEYINPUT118), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n971), .A2(KEYINPUT118), .ZN(new_n973));
  NOR3_X1   g0773(.A1(new_n970), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n963), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n951), .B1(new_n779), .B2(new_n956), .C1(new_n976), .C2(new_n726), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n653), .B1(new_n481), .B2(new_n485), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n641), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n500), .A2(new_n653), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n668), .A2(new_n666), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT44), .Z(new_n984));
  NOR2_X1   g0784(.A1(new_n981), .A2(new_n982), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT45), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(KEYINPUT116), .ZN(new_n988));
  INV_X1    g0788(.A(new_n665), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n987), .A2(KEYINPUT116), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT117), .ZN(new_n993));
  INV_X1    g0793(.A(new_n701), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n668), .B1(new_n664), .B2(new_n667), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n659), .B(new_n995), .Z(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n993), .B(new_n998), .C1(new_n989), .C2(new_n987), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n701), .ZN(new_n1000));
  XOR2_X1   g0800(.A(KEYINPUT115), .B(KEYINPUT41), .Z(new_n1001));
  XNOR2_X1  g0801(.A(new_n671), .B(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n708), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n981), .A2(new_n668), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT42), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n979), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n500), .B1(new_n1006), .B2(new_n679), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1005), .B1(new_n653), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n956), .A2(KEYINPUT43), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n956), .ZN(new_n1010));
  XOR2_X1   g0810(.A(KEYINPUT114), .B(KEYINPUT43), .Z(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1008), .A2(new_n1009), .A3(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n665), .A2(new_n981), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n977), .B1(new_n1003), .B2(new_n1016), .ZN(G387));
  AOI22_X1  g0817(.A1(new_n721), .A2(new_n672), .B1(new_n576), .B2(new_n670), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n235), .A2(new_n279), .ZN(new_n1019));
  AOI211_X1 g0819(.A(G45), .B(new_n672), .C1(G68), .C2(G77), .ZN(new_n1020));
  AND3_X1   g0820(.A1(new_n394), .A2(KEYINPUT50), .A3(new_n244), .ZN(new_n1021));
  AOI21_X1  g0821(.A(KEYINPUT50), .B1(new_n394), .B2(new_n244), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n713), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1018), .B1(new_n1019), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n710), .B1(new_n1025), .B2(new_n731), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G311), .A2(new_n760), .B1(new_n750), .B2(G322), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G303), .A2(new_n758), .B1(new_n755), .B2(G317), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1029), .A2(KEYINPUT48), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1027), .A2(KEYINPUT48), .A3(new_n1028), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n770), .A2(G283), .B1(new_n773), .B2(G294), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT49), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n735), .A2(new_n523), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n297), .B(new_n1037), .C1(G326), .C2(new_n739), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(G159), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n765), .A2(new_n1040), .B1(new_n759), .B2(new_n202), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G50), .B2(new_n755), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n744), .A2(new_n256), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n297), .B1(new_n738), .B2(new_n790), .C1(new_n519), .C2(new_n735), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1043), .B(new_n1044), .C1(new_n430), .C2(new_n770), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1042), .B(new_n1045), .C1(new_n350), .C2(new_n761), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1039), .A2(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT119), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1026), .B1(new_n664), .B2(new_n779), .C1(new_n1048), .C2(new_n726), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n671), .B1(new_n994), .B2(new_n997), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n701), .A2(new_n996), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n1049), .B1(new_n705), .B2(new_n997), .C1(new_n1050), .C2(new_n1051), .ZN(G393));
  XNOR2_X1  g0852(.A(new_n987), .B(new_n665), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n708), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n981), .A2(new_n730), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n297), .B(new_n772), .C1(G322), .C2(new_n739), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n770), .A2(G116), .B1(new_n773), .B2(G283), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n741), .B2(new_n759), .C1(new_n505), .C2(new_n761), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n750), .A2(G317), .B1(new_n755), .B2(G311), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT52), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n743), .A2(new_n256), .B1(new_n744), .B2(new_n202), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n377), .B1(new_n739), .B2(G143), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n223), .B2(new_n735), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n1062), .B(new_n1064), .C1(G50), .C2(new_n760), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n350), .B2(new_n759), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n750), .A2(G150), .B1(new_n755), .B2(G159), .ZN(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT51), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n1059), .A2(new_n1061), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n727), .ZN(new_n1070));
  OAI221_X1 g0870(.A(new_n731), .B1(new_n519), .B2(new_n210), .C1(new_n714), .C2(new_n242), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1055), .A2(new_n712), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n1054), .A2(KEYINPUT120), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(KEYINPUT120), .B1(new_n1054), .B2(new_n1072), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n671), .B1(new_n998), .B2(new_n1053), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1075), .B1(new_n999), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(G390));
  NAND2_X1  g0879(.A1(new_n934), .A2(G330), .ZN(new_n1080));
  OAI21_X1  g0880(.A(KEYINPUT121), .B1(new_n923), .B2(new_n834), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n916), .A2(new_n920), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n815), .A2(new_n922), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT121), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1084), .A2(new_n1085), .A3(new_n835), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n909), .A2(new_n912), .A3(new_n1081), .A4(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n922), .B1(new_n682), .B2(new_n813), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n834), .B1(new_n1088), .B2(new_n1082), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n939), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1080), .B1(new_n1087), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1082), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n700), .A2(new_n811), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1094), .B1(new_n939), .B2(new_n1089), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n908), .A2(new_n836), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n897), .A2(new_n898), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n912), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1081), .A2(new_n1086), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1095), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(KEYINPUT122), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT122), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1102), .B(new_n1095), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1091), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n909), .A2(new_n728), .A3(new_n912), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n784), .A2(new_n394), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n297), .B(new_n796), .C1(G294), .C2(new_n739), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1107), .B1(new_n256), .B2(new_n743), .C1(new_n576), .C2(new_n761), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n750), .A2(G283), .B1(new_n755), .B2(G116), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n1109), .B1(new_n519), .B2(new_n759), .C1(new_n223), .C2(new_n746), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n735), .A2(new_n244), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n377), .B(new_n1111), .C1(G125), .C2(new_n739), .ZN(new_n1112));
  INV_X1    g0912(.A(G128), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n1112), .B1(new_n1040), .B2(new_n743), .C1(new_n1113), .C2(new_n765), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n744), .A2(new_n790), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT53), .ZN(new_n1116));
  XOR2_X1   g0916(.A(KEYINPUT54), .B(G143), .Z(new_n1117));
  AOI22_X1  g0917(.A1(G132), .A2(new_n755), .B1(new_n758), .B2(new_n1117), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1116), .B(new_n1118), .C1(new_n789), .C2(new_n761), .ZN(new_n1119));
  OAI22_X1  g0919(.A1(new_n1108), .A2(new_n1110), .B1(new_n1114), .B2(new_n1119), .ZN(new_n1120));
  AOI211_X1 g0920(.A(new_n710), .B(new_n1106), .C1(new_n1120), .C2(new_n727), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1104), .A2(new_n708), .B1(new_n1105), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT123), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n941), .A2(G330), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n450), .A2(new_n1124), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n831), .A2(new_n370), .A3(new_n627), .A4(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1082), .B1(new_n1124), .B2(new_n811), .ZN(new_n1127));
  OR3_X1    g0927(.A1(new_n1094), .A2(new_n1127), .A3(new_n1088), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1080), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1082), .B1(new_n700), .B2(new_n811), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1083), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1126), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n671), .B1(new_n1104), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n1129), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1103), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1102), .B1(new_n1087), .B2(new_n1095), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1135), .B(new_n1132), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1122), .B(new_n1123), .C1(new_n1133), .C2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1126), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1142), .A2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1146), .A2(new_n671), .A3(new_n1138), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1123), .B1(new_n1147), .B2(new_n1122), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1141), .A2(new_n1148), .ZN(G378));
  NAND2_X1  g0949(.A1(new_n355), .A2(new_n857), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT124), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n371), .B(new_n1151), .ZN(new_n1152));
  XOR2_X1   g0952(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1153));
  XNOR2_X1  g0953(.A(new_n1152), .B(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n728), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n712), .B1(G50), .B2(new_n784), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n770), .A2(G150), .B1(new_n773), .B2(new_n1117), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n761), .B2(new_n793), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n1113), .A2(new_n804), .B1(new_n759), .B2(new_n789), .ZN(new_n1160));
  AOI211_X1 g0960(.A(new_n1159), .B(new_n1160), .C1(G125), .C2(new_n750), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  OR2_X1    g0962(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n787), .A2(new_n968), .ZN(new_n1165));
  AOI211_X1 g0965(.A(G33), .B(G41), .C1(new_n739), .C2(G124), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n765), .A2(new_n523), .B1(new_n804), .B2(new_n576), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n278), .B(new_n377), .C1(new_n738), .C2(new_n736), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n735), .A2(new_n201), .ZN(new_n1170));
  NOR4_X1   g0970(.A1(new_n1169), .A2(new_n964), .A3(new_n1043), .A4(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n429), .B2(new_n759), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1168), .B(new_n1172), .C1(G97), .C2(new_n760), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(KEYINPUT58), .ZN(new_n1174));
  OR2_X1    g0974(.A1(new_n1173), .A2(KEYINPUT58), .ZN(new_n1175));
  AOI21_X1  g0975(.A(G50), .B1(new_n253), .B2(new_n278), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n297), .B2(G41), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1167), .A2(new_n1174), .A3(new_n1175), .A4(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1157), .B1(new_n1178), .B2(new_n727), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1156), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n935), .A2(new_n936), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n937), .A2(new_n939), .ZN(new_n1183));
  AND4_X1   g0983(.A1(G330), .A2(new_n1182), .A3(new_n1183), .A4(new_n1154), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1154), .B1(new_n940), .B2(G330), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n1184), .A2(new_n1185), .B1(new_n913), .B2(new_n926), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT125), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1182), .A2(G330), .A3(new_n1183), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n1155), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1098), .A2(new_n834), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n926), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n940), .A2(G330), .A3(new_n1154), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1186), .A2(new_n1187), .A3(new_n1193), .ZN(new_n1194));
  OAI221_X1 g0994(.A(KEYINPUT125), .B1(new_n913), .B2(new_n926), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1181), .B1(new_n1196), .B2(new_n708), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1138), .A2(new_n1144), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT57), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1126), .B1(new_n1104), .B2(new_n1132), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1186), .A2(new_n1193), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(KEYINPUT57), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n671), .B1(new_n1200), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1197), .B1(new_n1199), .B2(new_n1203), .ZN(G375));
  NAND3_X1  g1004(.A1(new_n1126), .A2(new_n1128), .A3(new_n1131), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1145), .A2(new_n1002), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1092), .A2(new_n728), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n712), .B1(G68), .B2(new_n784), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1170), .A2(new_n377), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1209), .B(KEYINPUT127), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n790), .B2(new_n759), .C1(new_n1040), .C2(new_n746), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n760), .A2(new_n1117), .B1(new_n755), .B2(G137), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n770), .A2(G50), .B1(new_n739), .B2(G128), .ZN(new_n1213));
  OAI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(new_n793), .C2(new_n765), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n377), .B1(new_n735), .B2(new_n256), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n745), .A2(G97), .B1(KEYINPUT126), .B2(new_n1215), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n770), .A2(new_n430), .B1(new_n739), .B2(G303), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(KEYINPUT126), .C2(new_n1215), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n750), .A2(G294), .B1(new_n758), .B2(G107), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(new_n523), .B2(new_n761), .C1(new_n736), .C2(new_n804), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n1211), .A2(new_n1214), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1208), .B1(new_n1221), .B2(new_n727), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1143), .A2(new_n708), .B1(new_n1207), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1206), .A2(new_n1223), .ZN(G381));
  OR4_X1    g1024(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1225), .A2(G387), .A3(G381), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1122), .B1(new_n1133), .B2(new_n1139), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1180), .B1(new_n1229), .B2(new_n705), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1202), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n703), .B1(new_n1231), .B2(new_n1198), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT57), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n1200), .B2(new_n1229), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1230), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1226), .A2(new_n1228), .A3(new_n1235), .ZN(G407));
  NOR2_X1   g1036(.A1(new_n649), .A2(G343), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1235), .A2(new_n1228), .A3(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(G407), .A2(G213), .A3(new_n1238), .ZN(G409));
  NAND3_X1  g1039(.A1(new_n1196), .A2(new_n1002), .A3(new_n1198), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1181), .B1(new_n1201), .B2(new_n708), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1228), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1227), .A2(KEYINPUT123), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1140), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1243), .B1(new_n1245), .B2(G375), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1237), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1205), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1248), .A2(new_n1145), .A3(KEYINPUT60), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n671), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1248), .B1(KEYINPUT60), .B2(new_n1145), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1223), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(G384), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  OAI211_X1 g1054(.A(G384), .B(new_n1223), .C1(new_n1250), .C2(new_n1251), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1246), .A2(new_n1247), .A3(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(KEYINPUT62), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT61), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1237), .A2(G2897), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1254), .A2(new_n1255), .A3(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1260), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(G378), .A2(new_n1235), .B1(new_n1228), .B2(new_n1242), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1263), .B1(new_n1264), .B2(new_n1237), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT62), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1246), .A2(new_n1266), .A3(new_n1247), .A4(new_n1256), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1258), .A2(new_n1259), .A3(new_n1265), .A4(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(G387), .A2(new_n1078), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(G387), .A2(new_n1078), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(G393), .B(new_n781), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n1270), .A2(new_n1271), .A3(new_n1273), .ZN(new_n1274));
  OR2_X1    g1074(.A1(G387), .A2(new_n1078), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1272), .B1(new_n1275), .B2(new_n1269), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1268), .A2(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT63), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1257), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT61), .B1(new_n1282), .B2(new_n1263), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1246), .A2(KEYINPUT63), .A3(new_n1247), .A4(new_n1256), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1279), .A2(new_n1281), .A3(new_n1283), .A4(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1278), .A2(new_n1285), .ZN(G405));
  NAND2_X1  g1086(.A1(G378), .A2(new_n1235), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(G375), .A2(new_n1228), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  OR2_X1    g1089(.A1(new_n1289), .A2(new_n1256), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1256), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n1277), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1279), .A2(new_n1291), .A3(new_n1290), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(G402));
endmodule


