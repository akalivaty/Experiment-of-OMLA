

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738;

  OR2_X1 U371 ( .A1(n597), .A2(n513), .ZN(n515) );
  XNOR2_X2 U372 ( .A(G143), .B(G128), .ZN(n458) );
  AND2_X1 U373 ( .A1(n381), .A2(n380), .ZN(n379) );
  NAND2_X1 U374 ( .A1(n379), .A2(n376), .ZN(n606) );
  NAND2_X1 U375 ( .A1(n378), .A2(n377), .ZN(n376) );
  AND2_X1 U376 ( .A1(n383), .A2(n382), .ZN(n381) );
  NOR2_X1 U377 ( .A1(n677), .A2(n676), .ZN(n592) );
  OR2_X1 U378 ( .A1(G902), .A2(n698), .ZN(n421) );
  XNOR2_X1 U379 ( .A(n726), .B(G146), .ZN(n451) );
  XNOR2_X1 U380 ( .A(n408), .B(n481), .ZN(n356) );
  XNOR2_X1 U381 ( .A(KEYINPUT15), .B(G902), .ZN(n604) );
  BUF_X2 U382 ( .A(n540), .Z(n680) );
  XNOR2_X1 U383 ( .A(n452), .B(G472), .ZN(n540) );
  AND2_X1 U384 ( .A1(n592), .A2(n589), .ZN(n582) );
  XNOR2_X1 U385 ( .A(G146), .B(G125), .ZN(n481) );
  XNOR2_X1 U386 ( .A(n399), .B(n505), .ZN(n537) );
  NOR2_X1 U387 ( .A1(n560), .A2(n519), .ZN(n399) );
  AND2_X1 U388 ( .A1(n359), .A2(n357), .ZN(n571) );
  XNOR2_X1 U389 ( .A(n358), .B(KEYINPUT76), .ZN(n357) );
  XNOR2_X1 U390 ( .A(n444), .B(n374), .ZN(n492) );
  XNOR2_X1 U391 ( .A(KEYINPUT69), .B(KEYINPUT3), .ZN(n444) );
  XNOR2_X1 U392 ( .A(n375), .B(G119), .ZN(n374) );
  INV_X1 U393 ( .A(G101), .ZN(n375) );
  XOR2_X1 U394 ( .A(G116), .B(G107), .Z(n494) );
  NOR2_X1 U395 ( .A1(n604), .A2(n385), .ZN(n384) );
  NAND2_X1 U396 ( .A1(n650), .A2(n384), .ZN(n383) );
  XNOR2_X1 U397 ( .A(n484), .B(n409), .ZN(n726) );
  XNOR2_X1 U398 ( .A(n413), .B(G137), .ZN(n409) );
  XNOR2_X1 U399 ( .A(G134), .B(G131), .ZN(n413) );
  XNOR2_X1 U400 ( .A(n469), .B(n468), .ZN(n519) );
  INV_X1 U401 ( .A(G478), .ZN(n468) );
  XNOR2_X1 U402 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n422) );
  XNOR2_X1 U403 ( .A(G119), .B(G128), .ZN(n426) );
  XNOR2_X1 U404 ( .A(n395), .B(n394), .ZN(n425) );
  XNOR2_X1 U405 ( .A(G110), .B(KEYINPUT95), .ZN(n394) );
  XNOR2_X1 U406 ( .A(n396), .B(KEYINPUT94), .ZN(n395) );
  XNOR2_X1 U407 ( .A(KEYINPUT93), .B(G137), .ZN(n396) );
  XNOR2_X1 U408 ( .A(n412), .B(G140), .ZN(n408) );
  XNOR2_X1 U409 ( .A(KEYINPUT68), .B(KEYINPUT10), .ZN(n412) );
  XNOR2_X1 U410 ( .A(n471), .B(n407), .ZN(n406) );
  XNOR2_X1 U411 ( .A(n470), .B(n472), .ZN(n407) );
  INV_X1 U412 ( .A(KEYINPUT11), .ZN(n472) );
  XNOR2_X1 U413 ( .A(n373), .B(G122), .ZN(n491) );
  XNOR2_X1 U414 ( .A(G113), .B(G104), .ZN(n373) );
  XNOR2_X1 U415 ( .A(n400), .B(n355), .ZN(n575) );
  XNOR2_X1 U416 ( .A(n434), .B(n433), .ZN(n529) );
  XNOR2_X1 U417 ( .A(n432), .B(KEYINPUT25), .ZN(n433) );
  XNOR2_X1 U418 ( .A(n476), .B(n477), .ZN(n560) );
  XNOR2_X1 U419 ( .A(n386), .B(KEYINPUT0), .ZN(n597) );
  OR2_X1 U420 ( .A1(n567), .A2(n566), .ZN(n358) );
  NAND2_X1 U421 ( .A1(n360), .A2(n372), .ZN(n368) );
  NAND2_X1 U422 ( .A1(n361), .A2(n370), .ZN(n369) );
  NOR2_X1 U423 ( .A1(n573), .A2(KEYINPUT48), .ZN(n370) );
  INV_X1 U424 ( .A(KEYINPUT80), .ZN(n392) );
  INV_X1 U425 ( .A(G902), .ZN(n454) );
  XNOR2_X1 U426 ( .A(KEYINPUT100), .B(KEYINPUT12), .ZN(n470) );
  XNOR2_X1 U427 ( .A(n458), .B(KEYINPUT4), .ZN(n484) );
  NAND2_X1 U428 ( .A1(n368), .A2(n392), .ZN(n367) );
  INV_X1 U429 ( .A(n368), .ZN(n371) );
  XOR2_X1 U430 ( .A(KEYINPUT73), .B(KEYINPUT14), .Z(n438) );
  XNOR2_X1 U431 ( .A(n451), .B(n450), .ZN(n608) );
  XNOR2_X1 U432 ( .A(n492), .B(n491), .ZN(n496) );
  INV_X1 U433 ( .A(n655), .ZN(n378) );
  NAND2_X1 U434 ( .A1(n604), .A2(n385), .ZN(n382) );
  XNOR2_X1 U435 ( .A(G101), .B(G104), .ZN(n415) );
  INV_X2 U436 ( .A(G953), .ZN(n479) );
  AND2_X1 U437 ( .A1(n402), .A2(n401), .ZN(n548) );
  XNOR2_X1 U438 ( .A(n506), .B(KEYINPUT19), .ZN(n563) );
  AND2_X1 U439 ( .A1(n543), .A2(n581), .ZN(n546) );
  BUF_X1 U440 ( .A(n580), .Z(n587) );
  XNOR2_X1 U441 ( .A(n356), .B(n410), .ZN(n428) );
  XNOR2_X1 U442 ( .A(n467), .B(n466), .ZN(n704) );
  XNOR2_X1 U443 ( .A(n460), .B(n349), .ZN(n467) );
  XNOR2_X1 U444 ( .A(n405), .B(n403), .ZN(n618) );
  XNOR2_X1 U445 ( .A(n491), .B(n404), .ZN(n403) );
  XNOR2_X1 U446 ( .A(n475), .B(n473), .ZN(n404) );
  AND2_X1 U447 ( .A1(n611), .A2(G953), .ZN(n712) );
  XNOR2_X1 U448 ( .A(n550), .B(n549), .ZN(n738) );
  INV_X1 U449 ( .A(KEYINPUT40), .ZN(n549) );
  NOR2_X1 U450 ( .A1(n575), .A2(n641), .ZN(n550) );
  AND2_X1 U451 ( .A1(n459), .A2(G217), .ZN(n349) );
  XOR2_X1 U452 ( .A(KEYINPUT104), .B(KEYINPUT102), .Z(n350) );
  XNOR2_X1 U453 ( .A(n456), .B(KEYINPUT110), .ZN(n351) );
  AND2_X1 U454 ( .A1(n567), .A2(n568), .ZN(n352) );
  AND2_X1 U455 ( .A1(n546), .A2(n661), .ZN(n353) );
  AND2_X1 U456 ( .A1(n369), .A2(n363), .ZN(n354) );
  INV_X1 U457 ( .A(n574), .ZN(n393) );
  XOR2_X1 U458 ( .A(KEYINPUT82), .B(KEYINPUT39), .Z(n355) );
  XNOR2_X1 U459 ( .A(n356), .B(n406), .ZN(n405) );
  XNOR2_X1 U460 ( .A(n726), .B(n356), .ZN(n730) );
  NOR2_X1 U461 ( .A1(n569), .A2(n352), .ZN(n359) );
  NAND2_X1 U462 ( .A1(n572), .A2(KEYINPUT48), .ZN(n360) );
  INV_X1 U463 ( .A(n572), .ZN(n361) );
  NAND2_X1 U464 ( .A1(n364), .A2(n362), .ZN(n391) );
  NAND2_X1 U465 ( .A1(n354), .A2(n371), .ZN(n362) );
  NOR2_X1 U466 ( .A1(n574), .A2(n392), .ZN(n363) );
  AND2_X1 U467 ( .A1(n367), .A2(n365), .ZN(n364) );
  NAND2_X1 U468 ( .A1(n366), .A2(n392), .ZN(n365) );
  NAND2_X1 U469 ( .A1(n369), .A2(n393), .ZN(n366) );
  NAND2_X1 U470 ( .A1(n573), .A2(KEYINPUT48), .ZN(n372) );
  NAND2_X2 U471 ( .A1(n391), .A2(n736), .ZN(n655) );
  NOR2_X2 U472 ( .A1(n655), .A2(n650), .ZN(n652) );
  NOR2_X1 U473 ( .A1(n650), .A2(n498), .ZN(n377) );
  NAND2_X1 U474 ( .A1(n655), .A2(n384), .ZN(n380) );
  INV_X1 U475 ( .A(KEYINPUT79), .ZN(n385) );
  NAND2_X1 U476 ( .A1(n563), .A2(n512), .ZN(n386) );
  NAND2_X1 U477 ( .A1(n387), .A2(n601), .ZN(n603) );
  XNOR2_X1 U478 ( .A(n389), .B(n388), .ZN(n387) );
  INV_X1 U479 ( .A(KEYINPUT44), .ZN(n388) );
  NAND2_X1 U480 ( .A1(n390), .A2(n579), .ZN(n389) );
  NOR2_X1 U481 ( .A1(n737), .A2(n578), .ZN(n390) );
  NAND2_X1 U482 ( .A1(n738), .A2(n397), .ZN(n552) );
  XNOR2_X1 U483 ( .A(n397), .B(G137), .ZN(G39) );
  XNOR2_X1 U484 ( .A(n545), .B(n398), .ZN(n397) );
  INV_X1 U485 ( .A(KEYINPUT42), .ZN(n398) );
  INV_X1 U486 ( .A(n537), .ZN(n663) );
  INV_X1 U487 ( .A(n546), .ZN(n595) );
  NAND2_X1 U488 ( .A1(n353), .A2(n548), .ZN(n400) );
  INV_X1 U489 ( .A(n522), .ZN(n401) );
  XNOR2_X1 U490 ( .A(n457), .B(n351), .ZN(n402) );
  NAND2_X1 U491 ( .A1(n608), .A2(n454), .ZN(n452) );
  XNOR2_X2 U492 ( .A(n502), .B(n501), .ZN(n536) );
  OR2_X2 U493 ( .A1(n624), .A2(n498), .ZN(n502) );
  XOR2_X1 U494 ( .A(n427), .B(n426), .Z(n410) );
  XOR2_X1 U495 ( .A(n700), .B(n699), .Z(n411) );
  INV_X1 U496 ( .A(KEYINPUT72), .ZN(n570) );
  AND2_X1 U497 ( .A1(n541), .A2(n540), .ZN(n542) );
  BUF_X1 U498 ( .A(n650), .Z(n713) );
  NOR2_X1 U499 ( .A1(n664), .A2(n663), .ZN(n539) );
  XNOR2_X1 U500 ( .A(n543), .B(KEYINPUT1), .ZN(n580) );
  XNOR2_X1 U501 ( .A(n698), .B(n411), .ZN(n701) );
  INV_X1 U502 ( .A(KEYINPUT70), .ZN(n414) );
  XNOR2_X1 U503 ( .A(n414), .B(G110), .ZN(n487) );
  XOR2_X1 U504 ( .A(G140), .B(G107), .Z(n416) );
  XNOR2_X1 U505 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U506 ( .A(n487), .B(n417), .Z(n419) );
  NAND2_X1 U507 ( .A1(G227), .A2(n479), .ZN(n418) );
  XNOR2_X1 U508 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U509 ( .A(n451), .B(n420), .ZN(n698) );
  XNOR2_X2 U510 ( .A(n421), .B(G469), .ZN(n543) );
  NAND2_X1 U511 ( .A1(n479), .A2(G234), .ZN(n423) );
  XNOR2_X1 U512 ( .A(n423), .B(n422), .ZN(n459) );
  NAND2_X1 U513 ( .A1(G221), .A2(n459), .ZN(n424) );
  XNOR2_X1 U514 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U515 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n427) );
  XNOR2_X1 U516 ( .A(n429), .B(n428), .ZN(n710) );
  NOR2_X1 U517 ( .A1(G902), .A2(n710), .ZN(n434) );
  NAND2_X1 U518 ( .A1(n604), .A2(G234), .ZN(n430) );
  XNOR2_X1 U519 ( .A(n430), .B(KEYINPUT96), .ZN(n431) );
  XNOR2_X1 U520 ( .A(KEYINPUT20), .B(n431), .ZN(n435) );
  NAND2_X1 U521 ( .A1(G217), .A2(n435), .ZN(n432) );
  AND2_X1 U522 ( .A1(n435), .A2(G221), .ZN(n436) );
  XNOR2_X1 U523 ( .A(n436), .B(KEYINPUT21), .ZN(n671) );
  AND2_X1 U524 ( .A1(n529), .A2(n671), .ZN(n581) );
  NAND2_X1 U525 ( .A1(G234), .A2(G237), .ZN(n437) );
  XNOR2_X1 U526 ( .A(n438), .B(n437), .ZN(n439) );
  NAND2_X1 U527 ( .A1(G952), .A2(n439), .ZN(n692) );
  NOR2_X1 U528 ( .A1(G953), .A2(n692), .ZN(n510) );
  NAND2_X1 U529 ( .A1(n439), .A2(G902), .ZN(n440) );
  XOR2_X1 U530 ( .A(n440), .B(KEYINPUT91), .Z(n508) );
  OR2_X1 U531 ( .A1(n479), .A2(n508), .ZN(n441) );
  XNOR2_X1 U532 ( .A(KEYINPUT108), .B(n441), .ZN(n442) );
  NOR2_X1 U533 ( .A1(G900), .A2(n442), .ZN(n443) );
  NOR2_X1 U534 ( .A1(n510), .A2(n443), .ZN(n522) );
  XOR2_X1 U535 ( .A(KEYINPUT5), .B(KEYINPUT97), .Z(n446) );
  XNOR2_X1 U536 ( .A(G113), .B(G116), .ZN(n445) );
  XNOR2_X1 U537 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U538 ( .A(n492), .B(n447), .Z(n449) );
  NOR2_X1 U539 ( .A1(G953), .A2(G237), .ZN(n474) );
  NAND2_X1 U540 ( .A1(n474), .A2(G210), .ZN(n448) );
  XNOR2_X1 U541 ( .A(n449), .B(n448), .ZN(n450) );
  INV_X1 U542 ( .A(G237), .ZN(n453) );
  NAND2_X1 U543 ( .A1(n454), .A2(n453), .ZN(n499) );
  NAND2_X1 U544 ( .A1(n499), .A2(G214), .ZN(n455) );
  XNOR2_X1 U545 ( .A(n455), .B(KEYINPUT88), .ZN(n660) );
  NAND2_X1 U546 ( .A1(n540), .A2(n660), .ZN(n457) );
  XNOR2_X1 U547 ( .A(KEYINPUT111), .B(KEYINPUT30), .ZN(n456) );
  AND2_X1 U548 ( .A1(n546), .A2(n548), .ZN(n504) );
  XOR2_X1 U549 ( .A(n458), .B(n494), .Z(n460) );
  XOR2_X1 U550 ( .A(KEYINPUT101), .B(KEYINPUT103), .Z(n462) );
  XNOR2_X1 U551 ( .A(G134), .B(KEYINPUT9), .ZN(n461) );
  XNOR2_X1 U552 ( .A(n462), .B(n461), .ZN(n465) );
  XNOR2_X1 U553 ( .A(G122), .B(KEYINPUT7), .ZN(n463) );
  XNOR2_X1 U554 ( .A(n350), .B(n463), .ZN(n464) );
  XOR2_X1 U555 ( .A(n465), .B(n464), .Z(n466) );
  NOR2_X1 U556 ( .A1(n704), .A2(G902), .ZN(n469) );
  XNOR2_X1 U557 ( .A(KEYINPUT13), .B(G475), .ZN(n477) );
  XOR2_X1 U558 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n471) );
  XNOR2_X1 U559 ( .A(G143), .B(G131), .ZN(n473) );
  NAND2_X1 U560 ( .A1(G214), .A2(n474), .ZN(n475) );
  NOR2_X1 U561 ( .A1(G902), .A2(n618), .ZN(n476) );
  NAND2_X1 U562 ( .A1(n519), .A2(n560), .ZN(n478) );
  XNOR2_X1 U563 ( .A(n478), .B(KEYINPUT107), .ZN(n584) );
  NAND2_X1 U564 ( .A1(n479), .A2(G224), .ZN(n480) );
  XNOR2_X1 U565 ( .A(n480), .B(KEYINPUT75), .ZN(n482) );
  XNOR2_X1 U566 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U567 ( .A(n484), .B(n483), .ZN(n490) );
  XNOR2_X1 U568 ( .A(KEYINPUT86), .B(KEYINPUT17), .ZN(n486) );
  XNOR2_X1 U569 ( .A(KEYINPUT18), .B(KEYINPUT84), .ZN(n485) );
  XNOR2_X1 U570 ( .A(n486), .B(n485), .ZN(n488) );
  XNOR2_X1 U571 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U572 ( .A(n490), .B(n489), .ZN(n497) );
  INV_X1 U573 ( .A(KEYINPUT16), .ZN(n493) );
  XNOR2_X1 U574 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U575 ( .A(n496), .B(n495), .ZN(n719) );
  XNOR2_X1 U576 ( .A(n497), .B(n719), .ZN(n624) );
  INV_X1 U577 ( .A(n604), .ZN(n498) );
  NAND2_X1 U578 ( .A1(n499), .A2(G210), .ZN(n500) );
  XNOR2_X1 U579 ( .A(n500), .B(KEYINPUT87), .ZN(n501) );
  INV_X1 U580 ( .A(n536), .ZN(n553) );
  AND2_X1 U581 ( .A1(n584), .A2(n536), .ZN(n503) );
  AND2_X1 U582 ( .A1(n504), .A2(n503), .ZN(n558) );
  XOR2_X1 U583 ( .A(G143), .B(n558), .Z(G45) );
  INV_X1 U584 ( .A(KEYINPUT105), .ZN(n505) );
  NAND2_X1 U585 ( .A1(n537), .A2(n671), .ZN(n513) );
  NAND2_X1 U586 ( .A1(n536), .A2(n660), .ZN(n506) );
  XNOR2_X1 U587 ( .A(G898), .B(KEYINPUT89), .ZN(n716) );
  NAND2_X1 U588 ( .A1(n716), .A2(G953), .ZN(n507) );
  XNOR2_X1 U589 ( .A(n507), .B(KEYINPUT90), .ZN(n721) );
  NOR2_X1 U590 ( .A1(n721), .A2(n508), .ZN(n509) );
  OR2_X1 U591 ( .A1(n510), .A2(n509), .ZN(n511) );
  XNOR2_X1 U592 ( .A(n511), .B(KEYINPUT92), .ZN(n512) );
  XNOR2_X1 U593 ( .A(KEYINPUT71), .B(KEYINPUT22), .ZN(n514) );
  XNOR2_X1 U594 ( .A(n515), .B(n514), .ZN(n591) );
  OR2_X1 U595 ( .A1(n587), .A2(n529), .ZN(n516) );
  NOR2_X1 U596 ( .A1(n680), .A2(n516), .ZN(n517) );
  AND2_X1 U597 ( .A1(n591), .A2(n517), .ZN(n578) );
  XOR2_X1 U598 ( .A(G110), .B(n578), .Z(G12) );
  XNOR2_X1 U599 ( .A(KEYINPUT43), .B(KEYINPUT109), .ZN(n526) );
  INV_X1 U600 ( .A(KEYINPUT6), .ZN(n518) );
  XNOR2_X1 U601 ( .A(n680), .B(n518), .ZN(n589) );
  INV_X1 U602 ( .A(n519), .ZN(n559) );
  NAND2_X1 U603 ( .A1(n560), .A2(n559), .ZN(n641) );
  INV_X1 U604 ( .A(n529), .ZN(n520) );
  NAND2_X1 U605 ( .A1(n520), .A2(n671), .ZN(n521) );
  NOR2_X1 U606 ( .A1(n522), .A2(n521), .ZN(n541) );
  NAND2_X1 U607 ( .A1(n541), .A2(n660), .ZN(n523) );
  NOR2_X1 U608 ( .A1(n641), .A2(n523), .ZN(n524) );
  NAND2_X1 U609 ( .A1(n589), .A2(n524), .ZN(n554) );
  NOR2_X1 U610 ( .A1(n587), .A2(n554), .ZN(n525) );
  XOR2_X1 U611 ( .A(n526), .B(n525), .Z(n527) );
  NOR2_X1 U612 ( .A1(n527), .A2(n536), .ZN(n574) );
  XOR2_X1 U613 ( .A(n574), .B(G140), .Z(G42) );
  INV_X1 U614 ( .A(KEYINPUT106), .ZN(n528) );
  XNOR2_X1 U615 ( .A(n529), .B(n528), .ZN(n673) );
  NAND2_X1 U616 ( .A1(n673), .A2(n587), .ZN(n530) );
  NOR2_X1 U617 ( .A1(n589), .A2(n530), .ZN(n531) );
  NAND2_X1 U618 ( .A1(n591), .A2(n531), .ZN(n533) );
  XNOR2_X1 U619 ( .A(KEYINPUT65), .B(KEYINPUT32), .ZN(n532) );
  XNOR2_X1 U620 ( .A(n533), .B(n532), .ZN(n577) );
  XNOR2_X1 U621 ( .A(G119), .B(KEYINPUT127), .ZN(n534) );
  XNOR2_X1 U622 ( .A(n577), .B(n534), .ZN(G21) );
  XNOR2_X1 U623 ( .A(KEYINPUT74), .B(KEYINPUT38), .ZN(n535) );
  XNOR2_X1 U624 ( .A(n536), .B(n535), .ZN(n547) );
  INV_X1 U625 ( .A(n547), .ZN(n661) );
  NAND2_X1 U626 ( .A1(n661), .A2(n660), .ZN(n664) );
  XNOR2_X1 U627 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n538) );
  XNOR2_X1 U628 ( .A(n539), .B(n538), .ZN(n670) );
  XNOR2_X1 U629 ( .A(KEYINPUT28), .B(n542), .ZN(n544) );
  NAND2_X1 U630 ( .A1(n544), .A2(n543), .ZN(n565) );
  NOR2_X1 U631 ( .A1(n670), .A2(n565), .ZN(n545) );
  XOR2_X1 U632 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n551) );
  XNOR2_X1 U633 ( .A(n552), .B(n551), .ZN(n557) );
  NOR2_X1 U634 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U635 ( .A(n555), .B(KEYINPUT36), .ZN(n556) );
  NAND2_X1 U636 ( .A1(n556), .A2(n587), .ZN(n648) );
  NAND2_X1 U637 ( .A1(n557), .A2(n648), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n558), .B(KEYINPUT77), .ZN(n562) );
  NOR2_X1 U639 ( .A1(n560), .A2(n559), .ZN(n636) );
  INV_X1 U640 ( .A(n636), .ZN(n644) );
  NAND2_X1 U641 ( .A1(n644), .A2(n641), .ZN(n598) );
  INV_X1 U642 ( .A(n598), .ZN(n665) );
  NAND2_X1 U643 ( .A1(n665), .A2(KEYINPUT47), .ZN(n561) );
  NAND2_X1 U644 ( .A1(n562), .A2(n561), .ZN(n569) );
  INV_X1 U645 ( .A(n563), .ZN(n564) );
  NOR2_X2 U646 ( .A1(n565), .A2(n564), .ZN(n567) );
  INV_X1 U647 ( .A(KEYINPUT47), .ZN(n566) );
  NOR2_X1 U648 ( .A1(KEYINPUT47), .A2(n665), .ZN(n568) );
  XNOR2_X1 U649 ( .A(n571), .B(n570), .ZN(n572) );
  NOR2_X1 U650 ( .A1(n575), .A2(n644), .ZN(n576) );
  XNOR2_X1 U651 ( .A(n576), .B(KEYINPUT113), .ZN(n736) );
  INV_X1 U652 ( .A(n577), .ZN(n579) );
  INV_X1 U653 ( .A(n580), .ZN(n677) );
  INV_X1 U654 ( .A(n581), .ZN(n676) );
  XNOR2_X1 U655 ( .A(n582), .B(KEYINPUT33), .ZN(n668) );
  NOR2_X1 U656 ( .A1(n668), .A2(n597), .ZN(n583) );
  XNOR2_X1 U657 ( .A(n583), .B(KEYINPUT34), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U659 ( .A(n586), .B(KEYINPUT35), .ZN(n737) );
  OR2_X1 U660 ( .A1(n673), .A2(n587), .ZN(n588) );
  NOR2_X1 U661 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U662 ( .A1(n591), .A2(n590), .ZN(n630) );
  NAND2_X1 U663 ( .A1(n680), .A2(n592), .ZN(n685) );
  OR2_X1 U664 ( .A1(n597), .A2(n685), .ZN(n594) );
  INV_X1 U665 ( .A(KEYINPUT31), .ZN(n593) );
  XNOR2_X1 U666 ( .A(n594), .B(n593), .ZN(n643) );
  OR2_X1 U667 ( .A1(n680), .A2(n595), .ZN(n596) );
  OR2_X1 U668 ( .A1(n597), .A2(n596), .ZN(n632) );
  NAND2_X1 U669 ( .A1(n643), .A2(n632), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n599), .A2(n598), .ZN(n600) );
  AND2_X1 U671 ( .A1(n630), .A2(n600), .ZN(n601) );
  INV_X1 U672 ( .A(KEYINPUT45), .ZN(n602) );
  XNOR2_X2 U673 ( .A(n603), .B(n602), .ZN(n650) );
  XNOR2_X1 U674 ( .A(n652), .B(KEYINPUT2), .ZN(n605) );
  NOR2_X4 U675 ( .A1(n606), .A2(n605), .ZN(n708) );
  NAND2_X1 U676 ( .A1(n708), .A2(G472), .ZN(n610) );
  XOR2_X1 U677 ( .A(KEYINPUT114), .B(KEYINPUT62), .Z(n607) );
  XNOR2_X1 U678 ( .A(n608), .B(n607), .ZN(n609) );
  XNOR2_X1 U679 ( .A(n610), .B(n609), .ZN(n612) );
  INV_X1 U680 ( .A(G952), .ZN(n611) );
  NOR2_X2 U681 ( .A1(n612), .A2(n712), .ZN(n614) );
  XNOR2_X1 U682 ( .A(KEYINPUT83), .B(KEYINPUT63), .ZN(n613) );
  XNOR2_X1 U683 ( .A(n614), .B(n613), .ZN(G57) );
  NAND2_X1 U684 ( .A1(n708), .A2(G475), .ZN(n620) );
  XOR2_X1 U685 ( .A(KEYINPUT85), .B(KEYINPUT121), .Z(n616) );
  XNOR2_X1 U686 ( .A(KEYINPUT59), .B(KEYINPUT66), .ZN(n615) );
  XNOR2_X1 U687 ( .A(n616), .B(n615), .ZN(n617) );
  XNOR2_X1 U688 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U689 ( .A(n620), .B(n619), .ZN(n621) );
  NOR2_X2 U690 ( .A1(n621), .A2(n712), .ZN(n622) );
  XNOR2_X1 U691 ( .A(n622), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U692 ( .A1(n708), .A2(G210), .ZN(n626) );
  XOR2_X1 U693 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n623) );
  XNOR2_X1 U694 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U695 ( .A(n626), .B(n625), .ZN(n627) );
  NOR2_X2 U696 ( .A1(n627), .A2(n712), .ZN(n629) );
  XOR2_X1 U697 ( .A(KEYINPUT81), .B(KEYINPUT56), .Z(n628) );
  XNOR2_X1 U698 ( .A(n629), .B(n628), .ZN(G51) );
  XNOR2_X1 U699 ( .A(G101), .B(n630), .ZN(G3) );
  NOR2_X1 U700 ( .A1(n641), .A2(n632), .ZN(n631) );
  XOR2_X1 U701 ( .A(G104), .B(n631), .Z(G6) );
  NOR2_X1 U702 ( .A1(n644), .A2(n632), .ZN(n634) );
  XNOR2_X1 U703 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n633) );
  XNOR2_X1 U704 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U705 ( .A(G107), .B(n635), .ZN(G9) );
  XOR2_X1 U706 ( .A(G128), .B(KEYINPUT29), .Z(n638) );
  NAND2_X1 U707 ( .A1(n567), .A2(n636), .ZN(n637) );
  XNOR2_X1 U708 ( .A(n638), .B(n637), .ZN(G30) );
  INV_X1 U709 ( .A(n641), .ZN(n639) );
  NAND2_X1 U710 ( .A1(n567), .A2(n639), .ZN(n640) );
  XNOR2_X1 U711 ( .A(n640), .B(G146), .ZN(G48) );
  NOR2_X1 U712 ( .A1(n641), .A2(n643), .ZN(n642) );
  XOR2_X1 U713 ( .A(G113), .B(n642), .Z(G15) );
  NOR2_X1 U714 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U715 ( .A(G116), .B(n645), .Z(G18) );
  XOR2_X1 U716 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n647) );
  XNOR2_X1 U717 ( .A(G125), .B(KEYINPUT37), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n647), .B(n646), .ZN(n649) );
  XOR2_X1 U719 ( .A(n649), .B(n648), .Z(G27) );
  INV_X1 U720 ( .A(KEYINPUT2), .ZN(n656) );
  NAND2_X1 U721 ( .A1(n713), .A2(n656), .ZN(n651) );
  XNOR2_X1 U722 ( .A(n651), .B(KEYINPUT78), .ZN(n654) );
  NAND2_X1 U723 ( .A1(n652), .A2(KEYINPUT2), .ZN(n653) );
  NAND2_X1 U724 ( .A1(n654), .A2(n653), .ZN(n658) );
  AND2_X1 U725 ( .A1(n655), .A2(n656), .ZN(n657) );
  NOR2_X1 U726 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U727 ( .A1(G953), .A2(n659), .ZN(n696) );
  NOR2_X1 U728 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U729 ( .A1(n663), .A2(n662), .ZN(n667) );
  NOR2_X1 U730 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U731 ( .A1(n667), .A2(n666), .ZN(n669) );
  NOR2_X1 U732 ( .A1(n669), .A2(n668), .ZN(n689) );
  INV_X1 U733 ( .A(n671), .ZN(n672) );
  NAND2_X1 U734 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U735 ( .A(n674), .B(KEYINPUT117), .ZN(n675) );
  XNOR2_X1 U736 ( .A(KEYINPUT49), .B(n675), .ZN(n683) );
  XOR2_X1 U737 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n679) );
  NAND2_X1 U738 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U739 ( .A(n679), .B(n678), .ZN(n681) );
  NOR2_X1 U740 ( .A1(n681), .A2(n680), .ZN(n682) );
  NAND2_X1 U741 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U742 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U743 ( .A(KEYINPUT51), .B(n686), .ZN(n687) );
  NOR2_X1 U744 ( .A1(n670), .A2(n687), .ZN(n688) );
  NOR2_X1 U745 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U746 ( .A(n690), .B(KEYINPUT52), .ZN(n691) );
  NOR2_X1 U747 ( .A1(n692), .A2(n691), .ZN(n694) );
  NOR2_X1 U748 ( .A1(n670), .A2(n668), .ZN(n693) );
  NOR2_X1 U749 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U750 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U751 ( .A(KEYINPUT53), .B(n697), .Z(G75) );
  NAND2_X1 U752 ( .A1(n708), .A2(G469), .ZN(n702) );
  XOR2_X1 U753 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n700) );
  XNOR2_X1 U754 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n699) );
  XNOR2_X1 U755 ( .A(n702), .B(n701), .ZN(n703) );
  NOR2_X1 U756 ( .A1(n712), .A2(n703), .ZN(G54) );
  NAND2_X1 U757 ( .A1(n708), .A2(G478), .ZN(n706) );
  XNOR2_X1 U758 ( .A(n704), .B(KEYINPUT122), .ZN(n705) );
  XNOR2_X1 U759 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U760 ( .A1(n712), .A2(n707), .ZN(G63) );
  NAND2_X1 U761 ( .A1(n708), .A2(G217), .ZN(n709) );
  XNOR2_X1 U762 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U763 ( .A1(n712), .A2(n711), .ZN(G66) );
  NOR2_X1 U764 ( .A1(n713), .A2(G953), .ZN(n718) );
  NAND2_X1 U765 ( .A1(G953), .A2(G224), .ZN(n714) );
  XOR2_X1 U766 ( .A(KEYINPUT61), .B(n714), .Z(n715) );
  NOR2_X1 U767 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U768 ( .A1(n718), .A2(n717), .ZN(n724) );
  XNOR2_X1 U769 ( .A(n719), .B(G110), .ZN(n720) );
  XNOR2_X1 U770 ( .A(n720), .B(KEYINPUT123), .ZN(n722) );
  NAND2_X1 U771 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U772 ( .A(n724), .B(n723), .ZN(n725) );
  XNOR2_X1 U773 ( .A(KEYINPUT124), .B(n725), .ZN(G69) );
  INV_X1 U774 ( .A(n730), .ZN(n727) );
  XOR2_X1 U775 ( .A(n727), .B(n655), .Z(n728) );
  NOR2_X1 U776 ( .A1(G953), .A2(n728), .ZN(n729) );
  XNOR2_X1 U777 ( .A(KEYINPUT125), .B(n729), .ZN(n734) );
  XOR2_X1 U778 ( .A(G227), .B(n730), .Z(n731) );
  NAND2_X1 U779 ( .A1(n731), .A2(G900), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n732), .A2(G953), .ZN(n733) );
  NAND2_X1 U781 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U782 ( .A(KEYINPUT126), .B(n735), .ZN(G72) );
  XNOR2_X1 U783 ( .A(G134), .B(n736), .ZN(G36) );
  XOR2_X1 U784 ( .A(G122), .B(n737), .Z(G24) );
  XNOR2_X1 U785 ( .A(n738), .B(G131), .ZN(G33) );
endmodule

