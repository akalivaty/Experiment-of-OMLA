//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n203));
  NOR2_X1   g002(.A1(G29gat), .A2(G36gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT14), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT90), .ZN(new_n206));
  INV_X1    g005(.A(G29gat), .ZN(new_n207));
  INV_X1    g006(.A(G36gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NOR3_X1   g008(.A1(new_n203), .A2(new_n205), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n202), .A2(KEYINPUT15), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(KEYINPUT17), .ZN(new_n213));
  INV_X1    g012(.A(G8gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(G15gat), .B(G22gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT16), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(G1gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT91), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n214), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n217), .B1(G1gat), .B2(new_n215), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n219), .B(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n213), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G229gat), .A2(G233gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n212), .A2(new_n221), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT18), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n223), .A2(KEYINPUT18), .A3(new_n224), .A4(new_n225), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n212), .B(new_n221), .ZN(new_n230));
  XOR2_X1   g029(.A(new_n224), .B(KEYINPUT13), .Z(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n228), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(KEYINPUT88), .B(KEYINPUT11), .Z(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(KEYINPUT89), .ZN(new_n235));
  XOR2_X1   g034(.A(G113gat), .B(G141gat), .Z(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(G169gat), .B(G197gat), .Z(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT12), .Z(new_n240));
  XOR2_X1   g039(.A(new_n233), .B(new_n240), .Z(new_n241));
  XOR2_X1   g040(.A(G8gat), .B(G36gat), .Z(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT75), .ZN(new_n243));
  XNOR2_X1  g042(.A(G64gat), .B(G92gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT25), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n248));
  NAND2_X1  g047(.A1(G183gat), .A2(G190gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT64), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n251), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT64), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n250), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(G169gat), .A2(G176gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT23), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT23), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n259), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(G169gat), .A2(G176gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n247), .B1(new_n255), .B2(new_n262), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n264));
  OR2_X1    g063(.A1(new_n253), .A2(KEYINPUT66), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n253), .A2(KEYINPUT66), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(new_n250), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n264), .A2(KEYINPUT25), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G169gat), .ZN(new_n270));
  INV_X1    g069(.A(G176gat), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n271), .A3(KEYINPUT26), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT26), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n261), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n249), .B(new_n272), .C1(new_n274), .C2(new_n256), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G183gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT27), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT27), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G183gat), .ZN(new_n280));
  INV_X1    g079(.A(G190gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT28), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT27), .B(G183gat), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT28), .B1(new_n285), .B2(new_n281), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n276), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT67), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n282), .A2(new_n283), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n285), .A2(KEYINPUT28), .A3(new_n281), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n275), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT67), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n269), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT74), .B(KEYINPUT29), .ZN(new_n295));
  NAND2_X1  g094(.A1(G226gat), .A2(G233gat), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(G197gat), .B(G204gat), .ZN(new_n299));
  INV_X1    g098(.A(G218gat), .ZN(new_n300));
  OR2_X1    g099(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n299), .B1(new_n303), .B2(KEYINPUT22), .ZN(new_n304));
  XNOR2_X1  g103(.A(G211gat), .B(G218gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n299), .B(new_n305), .C1(new_n303), .C2(KEYINPUT22), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n292), .B1(new_n263), .B2(new_n268), .ZN(new_n311));
  INV_X1    g110(.A(new_n296), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n298), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n269), .A2(new_n287), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n312), .A2(KEYINPUT29), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n269), .A2(new_n289), .A3(new_n293), .A4(new_n312), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n310), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n246), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n317), .A2(new_n318), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n309), .ZN(new_n322));
  AOI22_X1  g121(.A1(new_n294), .A2(new_n297), .B1(new_n312), .B2(new_n311), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n310), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n322), .A2(new_n324), .A3(new_n245), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n320), .A2(new_n325), .A3(KEYINPUT30), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n314), .A2(new_n319), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT30), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(new_n328), .A3(new_n245), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G134gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n331), .A2(G127gat), .ZN(new_n332));
  INV_X1    g131(.A(G127gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G134gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G113gat), .B(G120gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n335), .B1(new_n336), .B2(KEYINPUT1), .ZN(new_n337));
  INV_X1    g136(.A(G120gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(G113gat), .ZN(new_n339));
  INV_X1    g138(.A(G113gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G120gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G127gat), .B(G134gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT1), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n337), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G155gat), .ZN(new_n347));
  INV_X1    g146(.A(G162gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G155gat), .A2(G162gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(G141gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(G148gat), .ZN(new_n353));
  INV_X1    g152(.A(G148gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(G141gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT2), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n351), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT77), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n357), .A2(new_n347), .A3(new_n348), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n354), .A2(G141gat), .ZN(new_n362));
  AOI22_X1  g161(.A1(new_n361), .A2(new_n350), .B1(new_n362), .B2(KEYINPUT76), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n353), .A2(new_n355), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n360), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n361), .A2(new_n350), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n352), .A2(KEYINPUT76), .A3(G148gat), .ZN(new_n368));
  AND4_X1   g167(.A1(new_n360), .A2(new_n367), .A3(new_n365), .A4(new_n368), .ZN(new_n369));
  OAI211_X1 g168(.A(new_n346), .B(new_n359), .C1(new_n366), .C2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT4), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT80), .ZN(new_n372));
  INV_X1    g171(.A(new_n365), .ZN(new_n373));
  NOR3_X1   g172(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n350), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n368), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT77), .B1(new_n373), .B2(new_n376), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n367), .A2(new_n365), .A3(new_n360), .A4(new_n368), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n358), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n379), .A2(new_n380), .A3(new_n346), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n371), .A2(new_n372), .A3(new_n381), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n379), .A2(KEYINPUT80), .A3(new_n380), .A4(new_n346), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(G225gat), .A2(G233gat), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n346), .B1(new_n379), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n359), .B1(new_n366), .B2(new_n369), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT3), .ZN(new_n390));
  AOI211_X1 g189(.A(KEYINPUT5), .B(new_n386), .C1(new_n388), .C2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n371), .A2(new_n381), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n388), .A2(new_n390), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n393), .A3(new_n385), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT5), .ZN(new_n395));
  INV_X1    g194(.A(new_n346), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n389), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n370), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n395), .B1(new_n398), .B2(new_n386), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n384), .A2(new_n391), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  XOR2_X1   g199(.A(KEYINPUT78), .B(KEYINPUT0), .Z(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT79), .ZN(new_n402));
  XNOR2_X1  g201(.A(G1gat), .B(G29gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n402), .B(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G57gat), .B(G85gat), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT84), .B1(new_n400), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT6), .B1(new_n400), .B2(new_n406), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n394), .A2(new_n399), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n386), .B1(new_n388), .B2(new_n390), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n410), .A2(new_n382), .A3(new_n395), .A4(new_n383), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n406), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT84), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n407), .A2(new_n408), .A3(new_n414), .A4(KEYINPUT86), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(KEYINPUT6), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n409), .A2(new_n411), .ZN(new_n418));
  INV_X1    g217(.A(new_n406), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n413), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI211_X1 g219(.A(KEYINPUT84), .B(new_n406), .C1(new_n409), .C2(new_n411), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT86), .B1(new_n422), .B2(new_n408), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n330), .B1(new_n417), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT87), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT87), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n426), .B(new_n330), .C1(new_n417), .C2(new_n423), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n269), .A2(new_n289), .A3(new_n346), .A4(new_n293), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT68), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI211_X1 g229(.A(new_n288), .B(new_n275), .C1(new_n290), .C2(new_n291), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n290), .A2(new_n291), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT67), .B1(new_n432), .B2(new_n276), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n434), .A2(KEYINPUT68), .A3(new_n346), .A4(new_n269), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n294), .A2(new_n396), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n430), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(G227gat), .A2(G233gat), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(KEYINPUT32), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT70), .ZN(new_n444));
  XOR2_X1   g243(.A(G15gat), .B(G43gat), .Z(new_n445));
  XNOR2_X1  g244(.A(new_n445), .B(KEYINPUT69), .ZN(new_n446));
  XNOR2_X1  g245(.A(G71gat), .B(G99gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n442), .A2(new_n443), .A3(new_n444), .A4(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT33), .B1(new_n437), .B2(new_n439), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT32), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(new_n437), .B2(new_n439), .ZN(new_n452));
  INV_X1    g251(.A(new_n448), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n450), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n448), .A2(KEYINPUT33), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n440), .A2(KEYINPUT32), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT70), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n449), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n437), .A2(new_n439), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT34), .B1(new_n439), .B2(KEYINPUT71), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT35), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n461), .B(new_n449), .C1(new_n454), .C2(new_n457), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT31), .B(G50gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(G228gat), .A2(G233gat), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT29), .ZN(new_n468));
  INV_X1    g267(.A(new_n308), .ZN(new_n469));
  AND2_X1   g268(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n470));
  NOR2_X1   g269(.A1(KEYINPUT73), .A2(G211gat), .ZN(new_n471));
  OAI21_X1  g270(.A(G218gat), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT22), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n305), .B1(new_n474), .B2(new_n299), .ZN(new_n475));
  OAI211_X1 g274(.A(KEYINPUT82), .B(new_n468), .C1(new_n469), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n387), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT82), .B1(new_n309), .B2(new_n468), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n389), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n379), .A2(new_n387), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n295), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(new_n310), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n467), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n309), .B1(new_n480), .B2(new_n295), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n309), .A2(new_n295), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n379), .B1(new_n485), .B2(new_n387), .ZN(new_n486));
  INV_X1    g285(.A(new_n467), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n466), .B1(new_n483), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G78gat), .B(G106gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(G22gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n485), .A2(new_n387), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(new_n389), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n482), .A2(new_n493), .A3(new_n467), .ZN(new_n494));
  INV_X1    g293(.A(new_n466), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n468), .B1(new_n469), .B2(new_n475), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT82), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n498), .A2(new_n387), .A3(new_n476), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n484), .B1(new_n499), .B2(new_n389), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n494), .B(new_n495), .C1(new_n500), .C2(new_n467), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n489), .A2(new_n491), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n491), .B1(new_n489), .B2(new_n501), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n463), .A2(new_n464), .A3(new_n465), .A4(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n425), .A2(new_n427), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n330), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n418), .A2(new_n419), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT6), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n409), .A2(new_n411), .A3(new_n406), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT81), .ZN(new_n513));
  AOI22_X1  g312(.A1(new_n512), .A2(new_n513), .B1(KEYINPUT6), .B2(new_n412), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n509), .A2(KEYINPUT81), .A3(new_n510), .A4(new_n511), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n508), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n516), .A2(new_n463), .A3(new_n465), .A4(new_n504), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT35), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n507), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n382), .A2(new_n383), .A3(new_n393), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n386), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n521), .B(KEYINPUT39), .C1(new_n386), .C2(new_n398), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT39), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n520), .A2(new_n523), .A3(new_n386), .ZN(new_n524));
  AND3_X1   g323(.A1(new_n524), .A2(KEYINPUT83), .A3(new_n406), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT83), .B1(new_n524), .B2(new_n406), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n522), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT40), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT85), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n526), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n524), .A2(KEYINPUT83), .A3(new_n406), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT85), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n532), .A2(new_n533), .A3(KEYINPUT40), .A4(new_n522), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n527), .A2(new_n528), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n330), .A2(new_n420), .A3(new_n421), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n529), .A2(new_n534), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n407), .A2(new_n408), .A3(new_n414), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT86), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT38), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT37), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n245), .B1(new_n327), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n322), .A2(new_n324), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT37), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n541), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n246), .B1(new_n544), .B2(KEYINPUT37), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n321), .A2(new_n310), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n323), .A2(new_n309), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT37), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n541), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n325), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n540), .A2(new_n553), .A3(new_n416), .A4(new_n415), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n537), .A2(new_n504), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT72), .ZN(new_n556));
  INV_X1    g355(.A(new_n465), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n442), .A2(new_n443), .A3(new_n448), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n444), .B1(new_n452), .B2(new_n455), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n461), .B1(new_n560), .B2(new_n449), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n556), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT36), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n511), .A2(new_n510), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n513), .B1(new_n565), .B2(new_n412), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n566), .A2(new_n515), .A3(new_n416), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n330), .ZN(new_n568));
  INV_X1    g367(.A(new_n504), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n463), .A2(new_n465), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n571), .A2(new_n556), .A3(KEYINPUT36), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n555), .A2(new_n564), .A3(new_n570), .A4(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n241), .B1(new_n519), .B2(new_n573), .ZN(new_n574));
  AND2_X1   g373(.A1(G71gat), .A2(G78gat), .ZN(new_n575));
  NOR2_X1   g374(.A1(G71gat), .A2(G78gat), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(G57gat), .B(G64gat), .Z(new_n578));
  INV_X1    g377(.A(KEYINPUT92), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n578), .B1(KEYINPUT9), .B2(new_n575), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT94), .ZN(new_n583));
  INV_X1    g382(.A(G85gat), .ZN(new_n584));
  INV_X1    g383(.A(G92gat), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(KEYINPUT94), .A2(G85gat), .A3(G92gat), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n586), .A2(KEYINPUT7), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G99gat), .B(G106gat), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT7), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n583), .B(new_n590), .C1(new_n584), .C2(new_n585), .ZN(new_n591));
  NAND2_X1  g390(.A1(G99gat), .A2(G106gat), .ZN(new_n592));
  AOI22_X1  g391(.A1(KEYINPUT8), .A2(new_n592), .B1(new_n584), .B2(new_n585), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n588), .A2(new_n589), .A3(new_n591), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT95), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n582), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n588), .A2(new_n591), .A3(new_n593), .ZN(new_n597));
  INV_X1    g396(.A(new_n589), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(new_n594), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n596), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G230gat), .A2(G233gat), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n603), .B(KEYINPUT96), .Z(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  OR2_X1    g405(.A1(new_n606), .A2(KEYINPUT98), .ZN(new_n607));
  XNOR2_X1  g406(.A(G120gat), .B(G148gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(G176gat), .B(G204gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  NAND2_X1  g409(.A1(new_n606), .A2(KEYINPUT98), .ZN(new_n611));
  AND3_X1   g410(.A1(new_n607), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT10), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n602), .A2(new_n613), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n601), .A2(KEYINPUT10), .A3(new_n582), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n605), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(KEYINPUT97), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n616), .A2(KEYINPUT97), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n612), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT99), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n612), .A2(KEYINPUT99), .A3(new_n617), .A4(new_n618), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT100), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n616), .A2(new_n624), .ZN(new_n625));
  OAI211_X1 g424(.A(KEYINPUT100), .B(new_n605), .C1(new_n614), .C2(new_n615), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n627), .A2(new_n607), .A3(new_n611), .ZN(new_n628));
  INV_X1    g427(.A(new_n610), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n623), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n213), .A2(new_n600), .ZN(new_n632));
  AND2_X1   g431(.A1(G232gat), .A2(G233gat), .ZN(new_n633));
  AOI22_X1  g432(.A1(new_n212), .A2(new_n601), .B1(KEYINPUT41), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(G190gat), .B(G218gat), .Z(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n633), .A2(KEYINPUT41), .ZN(new_n638));
  XNOR2_X1  g437(.A(G134gat), .B(G162gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n635), .A2(new_n636), .ZN(new_n642));
  OR3_X1    g441(.A1(new_n637), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n641), .B1(new_n642), .B2(new_n637), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n582), .A2(KEYINPUT21), .ZN(new_n646));
  XOR2_X1   g445(.A(G127gat), .B(G155gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n221), .B1(KEYINPUT21), .B2(new_n582), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(G231gat), .A2(G233gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT93), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G183gat), .B(G211gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n650), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n645), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n631), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n574), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n660), .A2(new_n567), .ZN(new_n661));
  XOR2_X1   g460(.A(KEYINPUT101), .B(G1gat), .Z(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1324gat));
  INV_X1    g462(.A(new_n660), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n508), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT16), .B(G8gat), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n667), .A2(KEYINPUT102), .A3(KEYINPUT42), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n214), .B1(new_n664), .B2(new_n508), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670));
  OAI22_X1  g469(.A1(new_n669), .A2(new_n670), .B1(new_n665), .B2(new_n666), .ZN(new_n671));
  AOI21_X1  g470(.A(KEYINPUT102), .B1(new_n667), .B2(KEYINPUT42), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n668), .B1(new_n671), .B2(new_n672), .ZN(G1325gat));
  NOR3_X1   g472(.A1(new_n660), .A2(G15gat), .A3(new_n571), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT36), .B1(new_n571), .B2(new_n556), .ZN(new_n675));
  AOI211_X1 g474(.A(KEYINPUT72), .B(new_n563), .C1(new_n463), .C2(new_n465), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n664), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n674), .B1(G15gat), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT103), .ZN(G1326gat));
  NOR2_X1   g480(.A1(new_n660), .A2(new_n504), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT43), .B(G22gat), .Z(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1327gat));
  AOI21_X1  g483(.A(new_n645), .B1(new_n519), .B2(new_n573), .ZN(new_n685));
  NOR3_X1   g484(.A1(new_n631), .A2(new_n241), .A3(new_n657), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n687), .A2(G29gat), .A3(new_n567), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n688), .B(KEYINPUT45), .Z(new_n689));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n690), .B1(new_n685), .B2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n645), .ZN(new_n693));
  AND4_X1   g492(.A1(new_n570), .A2(new_n555), .A3(new_n564), .A4(new_n572), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n505), .B1(new_n424), .B2(KEYINPUT87), .ZN(new_n695));
  AOI22_X1  g494(.A1(new_n695), .A2(new_n427), .B1(KEYINPUT35), .B2(new_n517), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n693), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n697), .A2(KEYINPUT104), .A3(KEYINPUT44), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n568), .B2(new_n569), .ZN(new_n701));
  AOI211_X1 g500(.A(KEYINPUT105), .B(new_n504), .C1(new_n567), .C2(new_n330), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n677), .A2(new_n703), .A3(new_n555), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n519), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n519), .A2(new_n704), .A3(KEYINPUT106), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n707), .A2(new_n691), .A3(new_n693), .A4(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n699), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n710), .A2(new_n686), .ZN(new_n711));
  INV_X1    g510(.A(new_n567), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n689), .B1(new_n713), .B2(new_n207), .ZN(G1328gat));
  NOR2_X1   g513(.A1(new_n631), .A2(new_n657), .ZN(new_n715));
  AOI211_X1 g514(.A(G36gat), .B(new_n645), .C1(KEYINPUT107), .C2(KEYINPUT46), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n574), .A2(new_n508), .A3(new_n715), .A4(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n717), .B(new_n718), .Z(new_n719));
  NAND2_X1  g518(.A1(new_n711), .A2(new_n508), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n719), .B1(new_n720), .B2(G36gat), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT108), .ZN(G1329gat));
  NOR3_X1   g521(.A1(new_n687), .A2(G43gat), .A3(new_n571), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n711), .A2(new_n678), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n723), .B1(new_n724), .B2(G43gat), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g525(.A(G50gat), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n727), .B1(new_n711), .B2(new_n569), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n569), .A2(new_n727), .ZN(new_n729));
  OAI21_X1  g528(.A(KEYINPUT48), .B1(new_n687), .B2(new_n729), .ZN(new_n730));
  OR2_X1    g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n731), .A2(KEYINPUT110), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n731), .A2(KEYINPUT110), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n687), .A2(new_n729), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT109), .Z(new_n735));
  NOR2_X1   g534(.A1(new_n728), .A2(new_n735), .ZN(new_n736));
  OAI22_X1  g535(.A1(new_n732), .A2(new_n733), .B1(KEYINPUT48), .B2(new_n736), .ZN(G1331gat));
  AND2_X1   g536(.A1(new_n707), .A2(new_n708), .ZN(new_n738));
  INV_X1    g537(.A(new_n241), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(new_n658), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(new_n631), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT111), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n712), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g545(.A1(new_n743), .A2(new_n330), .ZN(new_n747));
  NOR2_X1   g546(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n748));
  AND2_X1   g547(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(new_n747), .B2(new_n748), .ZN(G1333gat));
  OAI21_X1  g550(.A(G71gat), .B1(new_n743), .B2(new_n677), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n571), .A2(G71gat), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n752), .B1(new_n743), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g553(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n754), .B(new_n755), .ZN(G1334gat));
  NOR2_X1   g555(.A1(new_n743), .A2(new_n504), .ZN(new_n757));
  XOR2_X1   g556(.A(KEYINPUT113), .B(G78gat), .Z(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1335gat));
  OAI21_X1  g558(.A(KEYINPUT114), .B1(new_n739), .B2(new_n657), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT114), .ZN(new_n761));
  INV_X1    g560(.A(new_n657), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n241), .A2(new_n761), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n631), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n765), .B1(new_n699), .B2(new_n709), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G85gat), .B1(new_n767), .B2(new_n567), .ZN(new_n768));
  AOI22_X1  g567(.A1(new_n621), .A2(new_n622), .B1(new_n629), .B2(new_n628), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n645), .B1(new_n760), .B2(new_n763), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n705), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n705), .A2(KEYINPUT51), .A3(new_n770), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n769), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n775), .A2(new_n584), .A3(new_n712), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n768), .A2(new_n776), .ZN(G1336gat));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n330), .A2(G92gat), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n705), .A2(KEYINPUT51), .A3(new_n770), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT51), .B1(new_n705), .B2(new_n770), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n631), .B(new_n779), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  AOI211_X1 g581(.A(new_n330), .B(new_n765), .C1(new_n699), .C2(new_n709), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n778), .B(new_n782), .C1(new_n783), .C2(new_n585), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(KEYINPUT115), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n773), .A2(new_n774), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n786), .A2(new_n787), .A3(new_n631), .A4(new_n779), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n785), .B(new_n788), .C1(new_n783), .C2(new_n585), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT116), .B1(new_n789), .B2(KEYINPUT52), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n585), .B1(new_n766), .B2(new_n508), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n785), .A2(new_n788), .ZN(new_n792));
  OAI211_X1 g591(.A(KEYINPUT116), .B(KEYINPUT52), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n784), .B1(new_n790), .B2(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT117), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI211_X1 g596(.A(KEYINPUT117), .B(new_n784), .C1(new_n790), .C2(new_n794), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(G1337gat));
  OAI21_X1  g598(.A(G99gat), .B1(new_n767), .B2(new_n677), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n571), .A2(G99gat), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n775), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(G1338gat));
  OAI21_X1  g602(.A(G106gat), .B1(new_n767), .B2(new_n504), .ZN(new_n804));
  INV_X1    g603(.A(G106gat), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n775), .A2(new_n805), .A3(new_n569), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(new_n806), .B2(KEYINPUT118), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n807), .B(new_n809), .ZN(G1339gat));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n614), .A2(new_n615), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n811), .B1(new_n812), .B2(new_n604), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n618), .A2(new_n617), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n625), .A2(new_n811), .A3(new_n626), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(new_n629), .A3(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n623), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n814), .A2(KEYINPUT55), .A3(new_n629), .A4(new_n815), .ZN(new_n821));
  OR2_X1    g620(.A1(new_n233), .A2(new_n240), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n224), .B1(new_n223), .B2(new_n225), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n230), .A2(new_n231), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n239), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(new_n645), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n819), .A2(new_n820), .A3(new_n821), .A4(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n827), .A2(new_n623), .A3(new_n821), .A4(new_n818), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT119), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT120), .ZN(new_n832));
  INV_X1    g631(.A(new_n826), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n631), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(KEYINPUT120), .B1(new_n769), .B2(new_n826), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n739), .A2(new_n623), .A3(new_n821), .A4(new_n818), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n645), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n657), .B1(new_n831), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n740), .A2(new_n769), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n842), .A2(new_n571), .A3(new_n569), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(new_n712), .A3(new_n330), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n844), .A2(new_n340), .A3(new_n241), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n712), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT121), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n843), .A2(new_n848), .A3(new_n712), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n850), .A2(new_n330), .A3(new_n739), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n845), .B1(new_n851), .B2(new_n340), .ZN(G1340gat));
  NAND2_X1  g651(.A1(new_n631), .A2(new_n338), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT122), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n850), .A2(new_n330), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(G120gat), .B1(new_n844), .B2(new_n769), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1341gat));
  NAND4_X1  g656(.A1(new_n850), .A2(new_n333), .A3(new_n330), .A4(new_n657), .ZN(new_n858));
  OAI21_X1  g657(.A(G127gat), .B1(new_n844), .B2(new_n762), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1342gat));
  NOR2_X1   g659(.A1(new_n645), .A2(new_n508), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(G134gat), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n847), .A2(new_n849), .A3(new_n863), .ZN(new_n864));
  OR2_X1    g663(.A1(new_n864), .A2(KEYINPUT56), .ZN(new_n865));
  OAI21_X1  g664(.A(G134gat), .B1(new_n846), .B2(new_n862), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(KEYINPUT56), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(G1343gat));
  NOR3_X1   g667(.A1(new_n678), .A2(new_n567), .A3(new_n508), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n569), .B(new_n869), .C1(new_n839), .C2(new_n841), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(G141gat), .B1(new_n871), .B2(new_n739), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n569), .B1(new_n839), .B2(new_n841), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n869), .B1(new_n873), .B2(KEYINPUT57), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT123), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n631), .A2(new_n833), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n693), .B1(new_n876), .B2(new_n836), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n831), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n875), .B1(new_n879), .B2(new_n762), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n828), .A2(new_n830), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n875), .B(new_n762), .C1(new_n881), .C2(new_n877), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n840), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n569), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n874), .B1(KEYINPUT57), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n241), .A2(new_n352), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n872), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n888));
  OR3_X1    g687(.A1(new_n887), .A2(new_n888), .A3(KEYINPUT58), .ZN(new_n889));
  OAI21_X1  g688(.A(KEYINPUT58), .B1(new_n887), .B2(new_n888), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(G1344gat));
  INV_X1    g690(.A(KEYINPUT125), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n873), .A2(KEYINPUT57), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n657), .B1(new_n878), .B2(new_n829), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n894), .B(new_n569), .C1(new_n895), .C2(new_n841), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n893), .A2(new_n631), .A3(new_n869), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(G148gat), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n884), .A2(KEYINPUT57), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n839), .A2(new_n841), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(new_n894), .A3(new_n569), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n899), .A2(new_n631), .A3(new_n869), .A4(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n354), .A2(KEYINPUT59), .ZN(new_n903));
  AOI22_X1  g702(.A1(new_n898), .A2(KEYINPUT59), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n870), .A2(G148gat), .A3(new_n769), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n892), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n905), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n902), .A2(new_n903), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n909), .B1(new_n897), .B2(G148gat), .ZN(new_n910));
  OAI211_X1 g709(.A(KEYINPUT125), .B(new_n907), .C1(new_n908), .C2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n906), .A2(new_n911), .ZN(G1345gat));
  NAND3_X1  g711(.A1(new_n871), .A2(new_n347), .A3(new_n657), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n885), .A2(new_n657), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n347), .ZN(G1346gat));
  AND2_X1   g714(.A1(new_n885), .A2(new_n693), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n862), .A2(G162gat), .A3(new_n567), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n677), .ZN(new_n918));
  OAI22_X1  g717(.A1(new_n916), .A2(new_n348), .B1(new_n873), .B2(new_n918), .ZN(G1347gat));
  NOR2_X1   g718(.A1(new_n712), .A2(new_n330), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n843), .A2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n739), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT126), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n923), .A2(new_n924), .A3(G169gat), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n924), .B1(new_n923), .B2(G169gat), .ZN(new_n927));
  OAI22_X1  g726(.A1(new_n926), .A2(new_n927), .B1(G169gat), .B2(new_n923), .ZN(G1348gat));
  NOR2_X1   g727(.A1(new_n921), .A2(new_n769), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(new_n271), .ZN(G1349gat));
  OR3_X1    g729(.A1(new_n921), .A2(new_n285), .A3(new_n762), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n277), .B1(new_n921), .B2(new_n762), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n932), .B1(new_n931), .B2(new_n933), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(G1350gat));
  OAI22_X1  g735(.A1(new_n921), .A2(new_n645), .B1(KEYINPUT61), .B2(G190gat), .ZN(new_n937));
  NAND2_X1  g736(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n937), .B(new_n938), .ZN(G1351gat));
  INV_X1    g738(.A(new_n920), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n678), .A2(new_n504), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n900), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(G197gat), .B1(new_n943), .B2(new_n739), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n678), .A2(new_n940), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n893), .A2(new_n896), .A3(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n739), .A2(G197gat), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(G1352gat));
  OR3_X1    g748(.A1(new_n942), .A2(G204gat), .A3(new_n769), .ZN(new_n950));
  XOR2_X1   g749(.A(new_n950), .B(KEYINPUT62), .Z(new_n951));
  OAI21_X1  g750(.A(G204gat), .B1(new_n946), .B2(new_n769), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1353gat));
  NAND4_X1  g752(.A1(new_n943), .A2(new_n301), .A3(new_n302), .A4(new_n657), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n893), .A2(new_n657), .A3(new_n896), .A4(new_n945), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n955), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n956));
  AOI21_X1  g755(.A(KEYINPUT63), .B1(new_n955), .B2(G211gat), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT127), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI211_X1 g759(.A(KEYINPUT127), .B(new_n954), .C1(new_n956), .C2(new_n957), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1354gat));
  OAI21_X1  g761(.A(G218gat), .B1(new_n946), .B2(new_n645), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n943), .A2(new_n300), .A3(new_n693), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1355gat));
endmodule


