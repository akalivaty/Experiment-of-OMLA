//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n567,
    new_n568, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G259));
  XOR2_X1   g019(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(KEYINPUT69), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT69), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n461), .A2(new_n463), .A3(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n467), .A2(KEYINPUT3), .A3(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n470), .A2(G137), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n464), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT70), .ZN(new_n473));
  XNOR2_X1  g048(.A(new_n472), .B(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n462), .A2(G2104), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n475), .A2(new_n476), .A3(G125), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n480));
  AOI22_X1  g055(.A1(new_n479), .A2(G2105), .B1(G101), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n474), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  AND2_X1   g058(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n484));
  NOR2_X1   g059(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n466), .B1(KEYINPUT69), .B2(new_n462), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n486), .A2(KEYINPUT3), .B1(new_n487), .B2(new_n461), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(new_n470), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G136), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G124), .ZN(new_n494));
  OR2_X1    g069(.A1(G100), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n491), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G162));
  AND2_X1   g073(.A1(new_n470), .A2(G138), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n464), .A2(new_n469), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  OAI211_X1 g077(.A(G138), .B(new_n470), .C1(new_n502), .C2(KEYINPUT71), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n502), .A2(KEYINPUT71), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n475), .A2(new_n476), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n464), .A2(new_n469), .A3(G126), .A4(G2105), .ZN(new_n509));
  OR2_X1    g084(.A1(G102), .A2(G2105), .ZN(new_n510));
  OAI211_X1 g085(.A(new_n510), .B(G2104), .C1(G114), .C2(new_n470), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n508), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n500), .A2(KEYINPUT4), .B1(new_n506), .B2(new_n505), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n509), .A2(new_n511), .ZN(new_n516));
  OAI21_X1  g091(.A(KEYINPUT72), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(G164));
  OAI21_X1  g094(.A(KEYINPUT5), .B1(KEYINPUT73), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n520), .B1(KEYINPUT74), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT74), .ZN(new_n523));
  NAND4_X1  g098(.A1(new_n523), .A2(KEYINPUT73), .A3(KEYINPUT5), .A4(G543), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n525), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n526));
  INV_X1    g101(.A(G651), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n531), .B1(new_n522), .B2(new_n524), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n521), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n532), .A2(G88), .B1(new_n533), .B2(G50), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n528), .A2(new_n534), .ZN(G303));
  INV_X1    g110(.A(G303), .ZN(G166));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  INV_X1    g113(.A(new_n531), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n525), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G89), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(KEYINPUT75), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n544), .B(new_n538), .C1(new_n540), .C2(new_n541), .ZN(new_n545));
  AND2_X1   g120(.A1(G63), .A2(G651), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n533), .A2(G51), .B1(new_n525), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n543), .A2(new_n545), .A3(new_n547), .ZN(G286));
  INV_X1    g123(.A(G286), .ZN(G168));
  AOI22_X1  g124(.A1(new_n525), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n527), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n532), .A2(G90), .B1(new_n533), .B2(G52), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  AOI22_X1  g129(.A1(new_n532), .A2(G81), .B1(new_n533), .B2(G43), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  AND2_X1   g132(.A1(new_n522), .A2(new_n524), .ZN(new_n558));
  INV_X1    g133(.A(G56), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n527), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI211_X1 g137(.A(KEYINPUT76), .B(new_n557), .C1(new_n558), .C2(new_n559), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n556), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(G153));
  NAND4_X1  g140(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g141(.A1(G1), .A2(G3), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g143(.A1(G319), .A2(G483), .A3(G661), .A4(new_n568), .ZN(G188));
  NAND2_X1  g144(.A1(new_n533), .A2(G53), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT9), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n572), .B2(KEYINPUT77), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n522), .B2(new_n524), .ZN(new_n577));
  AND2_X1   g152(.A1(G78), .A2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n532), .A2(G91), .ZN(new_n580));
  NAND2_X1  g155(.A1(KEYINPUT78), .A2(KEYINPUT9), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n533), .A2(G53), .A3(new_n573), .A4(new_n581), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n575), .A2(new_n579), .A3(new_n580), .A4(new_n582), .ZN(G299));
  NAND2_X1  g158(.A1(new_n532), .A2(G87), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n525), .B2(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n533), .A2(G49), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G288));
  AND2_X1   g162(.A1(new_n525), .A2(G61), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT79), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n532), .A2(G86), .B1(new_n533), .B2(G48), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(new_n532), .A2(G85), .B1(new_n533), .B2(G47), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n525), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n527), .B2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n597), .B(KEYINPUT80), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT10), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n532), .A2(new_n600), .A3(G92), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n600), .B1(new_n532), .B2(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n599), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT81), .B1(new_n540), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n606), .A2(new_n601), .A3(KEYINPUT10), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G66), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n558), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n610), .A2(G651), .B1(G54), .B2(new_n533), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n604), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n598), .B1(G868), .B2(new_n613), .ZN(G284));
  OAI21_X1  g189(.A(new_n598), .B1(G868), .B2(new_n613), .ZN(G321));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(G299), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G168), .B2(new_n616), .ZN(G297));
  OAI21_X1  g193(.A(new_n617), .B1(G168), .B2(new_n616), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n562), .A2(new_n563), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(new_n555), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(new_n616), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n612), .A2(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(new_n616), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g202(.A1(new_n506), .A2(new_n480), .ZN(new_n628));
  XOR2_X1   g203(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(KEYINPUT83), .B(KEYINPUT13), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(G2100), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT84), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n490), .A2(G135), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n493), .A2(G123), .ZN(new_n637));
  OR2_X1    g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n638), .B(G2104), .C1(G111), .C2(new_n470), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(G2096), .ZN(new_n642));
  AOI22_X1  g217(.A1(new_n633), .A2(new_n632), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n635), .B(new_n643), .C1(new_n642), .C2(new_n641), .ZN(G156));
  INV_X1    g219(.A(G14), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n649), .A2(KEYINPUT14), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n651), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2443), .B(G2446), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1341), .B(G1348), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT85), .ZN(new_n660));
  AOI211_X1 g235(.A(new_n645), .B(new_n660), .C1(new_n658), .C2(new_n656), .ZN(G401));
  INV_X1    g236(.A(KEYINPUT18), .ZN(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(KEYINPUT17), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(new_n633), .ZN(new_n669));
  XOR2_X1   g244(.A(G2072), .B(G2078), .Z(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n665), .B2(KEYINPUT18), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(new_n642), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n669), .B(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(new_n678), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT20), .Z(new_n682));
  AOI211_X1 g257(.A(new_n680), .B(new_n682), .C1(new_n675), .C2(new_n679), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT86), .ZN(new_n684));
  XOR2_X1   g259(.A(G1981), .B(G1986), .Z(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n684), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(G229));
  MUX2_X1   g266(.A(G6), .B(G305), .S(G16), .Z(new_n692));
  XOR2_X1   g267(.A(KEYINPUT32), .B(G1981), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n694), .A2(KEYINPUT90), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(KEYINPUT90), .ZN(new_n696));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G22), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G166), .B2(new_n697), .ZN(new_n699));
  INV_X1    g274(.A(G1971), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n697), .A2(G23), .ZN(new_n702));
  INV_X1    g277(.A(G288), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n697), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT33), .B(G1976), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n695), .A2(new_n696), .A3(new_n701), .A4(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT89), .B(KEYINPUT34), .Z(new_n708));
  OR2_X1    g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT88), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n697), .B1(G290), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n711), .B2(G290), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n697), .A2(G24), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT87), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n716), .A2(G1986), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n490), .A2(G131), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n493), .A2(G119), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n470), .A2(G107), .ZN(new_n720));
  OAI21_X1  g295(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n718), .B(new_n719), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  MUX2_X1   g297(.A(G25), .B(new_n722), .S(G29), .Z(new_n723));
  XOR2_X1   g298(.A(KEYINPUT35), .B(G1991), .Z(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n723), .B(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G1986), .B2(new_n716), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n709), .A2(new_n710), .A3(new_n717), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT36), .ZN(new_n729));
  INV_X1    g304(.A(G29), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n730), .A2(G26), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT93), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT28), .ZN(new_n733));
  OR2_X1    g308(.A1(G104), .A2(G2105), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n734), .B(G2104), .C1(G116), .C2(new_n470), .ZN(new_n735));
  INV_X1    g310(.A(G140), .ZN(new_n736));
  INV_X1    g311(.A(G128), .ZN(new_n737));
  OAI221_X1 g312(.A(new_n735), .B1(new_n489), .B2(new_n736), .C1(new_n737), .C2(new_n492), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n738), .A2(KEYINPUT92), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(KEYINPUT92), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n733), .B1(new_n741), .B2(G29), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT94), .B(G2067), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n742), .B(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G34), .ZN(new_n745));
  AOI21_X1  g320(.A(G29), .B1(new_n745), .B2(KEYINPUT24), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(KEYINPUT24), .B2(new_n745), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n482), .B2(new_n730), .ZN(new_n748));
  INV_X1    g323(.A(G2084), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(KEYINPUT96), .ZN(new_n751));
  NOR2_X1   g326(.A1(G4), .A2(G16), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(new_n613), .B2(G16), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT91), .B(G1348), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n697), .A2(G20), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT98), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT23), .ZN(new_n758));
  INV_X1    g333(.A(G299), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n759), .B2(new_n697), .ZN(new_n760));
  INV_X1    g335(.A(G1956), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n750), .A2(KEYINPUT96), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR4_X1   g339(.A1(new_n744), .A2(new_n751), .A3(new_n755), .A4(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n730), .A2(G35), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G162), .B2(new_n730), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT29), .Z(new_n768));
  INV_X1    g343(.A(G2090), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(G168), .A2(G16), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G16), .B2(G21), .ZN(new_n772));
  INV_X1    g347(.A(G1966), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G16), .A2(G19), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n564), .B2(G16), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(G1341), .Z(new_n777));
  NAND3_X1  g352(.A1(new_n770), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g353(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT25), .ZN(new_n780));
  AOI22_X1  g355(.A1(new_n506), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(new_n470), .ZN(new_n782));
  AOI211_X1 g357(.A(new_n780), .B(new_n782), .C1(G139), .C2(new_n490), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G29), .ZN(new_n784));
  OR2_X1    g359(.A1(G29), .A2(G33), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT95), .B(G2072), .ZN(new_n786));
  AND3_X1   g361(.A1(new_n784), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n786), .B1(new_n784), .B2(new_n785), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT30), .B(G28), .ZN(new_n789));
  OR2_X1    g364(.A1(KEYINPUT31), .A2(G11), .ZN(new_n790));
  NAND2_X1  g365(.A1(KEYINPUT31), .A2(G11), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n789), .A2(new_n730), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n640), .B2(new_n730), .ZN(new_n793));
  NOR3_X1   g368(.A1(new_n787), .A2(new_n788), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G5), .A2(G16), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G171), .B2(G16), .ZN(new_n796));
  INV_X1    g371(.A(G1961), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n748), .A2(new_n749), .ZN(new_n799));
  NAND3_X1  g374(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT26), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  AOI22_X1  g378(.A1(G105), .A2(new_n480), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(G141), .ZN(new_n805));
  INV_X1    g380(.A(G129), .ZN(new_n806));
  OAI221_X1 g381(.A(new_n804), .B1(new_n489), .B2(new_n805), .C1(new_n806), .C2(new_n492), .ZN(new_n807));
  MUX2_X1   g382(.A(G32), .B(new_n807), .S(G29), .Z(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT27), .B(G1996), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n794), .A2(new_n798), .A3(new_n799), .A4(new_n810), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n768), .A2(new_n769), .B1(new_n773), .B2(new_n772), .ZN(new_n812));
  NOR3_X1   g387(.A1(new_n778), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n730), .A2(G27), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(G164), .B2(new_n730), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT97), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G2078), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n729), .A2(new_n765), .A3(new_n813), .A4(new_n817), .ZN(G150));
  INV_X1    g393(.A(G150), .ZN(G311));
  AOI22_X1  g394(.A1(new_n532), .A2(G93), .B1(new_n533), .B2(G55), .ZN(new_n820));
  NAND2_X1  g395(.A1(G80), .A2(G543), .ZN(new_n821));
  INV_X1    g396(.A(G67), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n558), .B2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT99), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n525), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n826));
  OAI21_X1  g401(.A(G651), .B1(new_n826), .B2(KEYINPUT99), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n820), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT100), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g405(.A(KEYINPUT100), .B(new_n820), .C1(new_n825), .C2(new_n827), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n830), .A2(new_n623), .A3(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n825), .A2(new_n827), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n564), .A2(new_n833), .A3(KEYINPUT100), .A4(new_n820), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT38), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n613), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n840));
  NOR3_X1   g415(.A1(new_n839), .A2(new_n840), .A3(G860), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n828), .A2(G860), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT37), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n841), .A2(new_n843), .ZN(G145));
  NOR2_X1   g419(.A1(new_n515), .A2(new_n516), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n741), .B(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n807), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n783), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n722), .B(KEYINPUT101), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n493), .A2(G130), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n470), .A2(G118), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(G142), .B2(new_n490), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n849), .B(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n630), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n848), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n497), .B(new_n640), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n482), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n848), .A2(new_n856), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n857), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n856), .A2(KEYINPUT102), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n859), .B1(new_n848), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n848), .B2(new_n862), .ZN(new_n864));
  INV_X1    g439(.A(G37), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n861), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g442(.A1(new_n828), .A2(new_n616), .ZN(new_n868));
  XOR2_X1   g443(.A(G305), .B(G290), .Z(new_n869));
  XNOR2_X1  g444(.A(G303), .B(new_n703), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n869), .B(new_n870), .Z(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n872), .A2(KEYINPUT105), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT42), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n612), .A2(new_n759), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n604), .A2(G299), .A3(new_n607), .A4(new_n611), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT103), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n612), .A2(KEYINPUT103), .A3(new_n759), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(new_n876), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT41), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(KEYINPUT104), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n881), .A2(new_n885), .A3(new_n882), .ZN(new_n886));
  AND2_X1   g461(.A1(new_n876), .A2(KEYINPUT41), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n875), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n884), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n835), .B(new_n625), .ZN(new_n890));
  MUX2_X1   g465(.A(new_n877), .B(new_n889), .S(new_n890), .Z(new_n891));
  XOR2_X1   g466(.A(new_n874), .B(new_n891), .Z(new_n892));
  OAI21_X1  g467(.A(new_n868), .B1(new_n892), .B2(new_n616), .ZN(G295));
  OAI21_X1  g468(.A(new_n868), .B1(new_n892), .B2(new_n616), .ZN(G331));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n551), .A2(KEYINPUT106), .A3(new_n552), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT106), .B1(new_n551), .B2(new_n552), .ZN(new_n899));
  OAI21_X1  g474(.A(G168), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n901), .A2(G286), .A3(new_n897), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n835), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n832), .A2(new_n900), .A3(new_n902), .A4(new_n834), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(new_n877), .A3(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT107), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n905), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n889), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n909), .A3(new_n872), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n910), .A2(new_n865), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n907), .A2(new_n909), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(new_n871), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n896), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n879), .A2(new_n887), .A3(new_n880), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n877), .A2(new_n882), .ZN(new_n916));
  AOI22_X1  g491(.A1(new_n904), .A2(new_n905), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n906), .B1(new_n917), .B2(new_n918), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n871), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n910), .A2(new_n865), .A3(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n922), .A2(KEYINPUT43), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n895), .B1(new_n914), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n895), .B1(new_n922), .B2(KEYINPUT43), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n913), .A2(new_n896), .A3(new_n865), .A4(new_n910), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n925), .A2(KEYINPUT109), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(KEYINPUT109), .B1(new_n925), .B2(new_n926), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n924), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT110), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n924), .B(KEYINPUT110), .C1(new_n927), .C2(new_n928), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(G397));
  AOI21_X1  g508(.A(KEYINPUT70), .B1(new_n488), .B2(new_n471), .ZN(new_n934));
  AND4_X1   g509(.A1(KEYINPUT70), .A2(new_n464), .A3(new_n469), .A4(new_n471), .ZN(new_n935));
  OAI211_X1 g510(.A(G40), .B(new_n481), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n474), .A2(KEYINPUT111), .A3(G40), .A4(new_n481), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G1384), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(new_n515), .B2(new_n516), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n940), .A2(new_n945), .ZN(new_n946));
  OR3_X1    g521(.A1(new_n946), .A2(G1986), .A3(G290), .ZN(new_n947));
  INV_X1    g522(.A(new_n946), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n948), .A2(G1986), .A3(G290), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g525(.A(new_n950), .B(KEYINPUT112), .Z(new_n951));
  NAND2_X1  g526(.A1(new_n741), .A2(G2067), .ZN(new_n952));
  INV_X1    g527(.A(G2067), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n739), .A2(new_n953), .A3(new_n740), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n807), .B(G1996), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n722), .B(new_n724), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n948), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n951), .A2(new_n960), .ZN(new_n961));
  OAI211_X1 g536(.A(KEYINPUT45), .B(new_n941), .C1(new_n515), .C2(new_n516), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n938), .A2(new_n939), .A3(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n513), .B1(new_n508), .B2(new_n512), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT72), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n941), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n943), .ZN(new_n968));
  AOI21_X1  g543(.A(G1971), .B1(new_n964), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n970), .B1(new_n518), .B2(new_n941), .ZN(new_n971));
  OAI211_X1 g546(.A(new_n970), .B(new_n941), .C1(new_n515), .C2(new_n516), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n938), .A2(new_n939), .A3(new_n972), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n971), .A2(new_n973), .A3(G2090), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT113), .B1(new_n969), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT45), .B1(new_n518), .B2(new_n941), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n700), .B1(new_n976), .B2(new_n963), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n938), .A2(new_n939), .A3(new_n972), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n967), .A2(KEYINPUT50), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n977), .B(new_n978), .C1(new_n981), .C2(G2090), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n975), .A2(G8), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G8), .ZN(new_n984));
  NOR2_X1   g559(.A1(G166), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g560(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n986));
  OR2_X1    g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n985), .B1(KEYINPUT114), .B2(KEYINPUT55), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n983), .A2(new_n990), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n975), .A2(G8), .A3(new_n982), .A4(new_n989), .ZN(new_n992));
  INV_X1    g567(.A(new_n942), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n938), .A2(new_n939), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(G8), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n703), .A2(G1976), .ZN(new_n997));
  INV_X1    g572(.A(G1976), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT52), .B1(G288), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n996), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(G305), .A2(G1981), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT49), .ZN(new_n1002));
  INV_X1    g577(.A(G1981), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n1003), .B1(new_n591), .B2(new_n592), .ZN(new_n1004));
  OR3_X1    g579(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1002), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n996), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n994), .A2(G8), .A3(new_n997), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT52), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n1000), .A2(new_n1007), .A3(new_n1009), .ZN(new_n1010));
  AOI211_X1 g585(.A(new_n943), .B(G1384), .C1(new_n514), .C2(new_n517), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n938), .A2(new_n944), .A3(new_n939), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n773), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(new_n981), .B2(G2084), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(G8), .A3(G168), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT63), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n991), .A2(new_n992), .A3(new_n1010), .A4(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n992), .A2(new_n1010), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n942), .A2(KEYINPUT50), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n938), .A2(new_n1020), .A3(new_n939), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n518), .A2(new_n970), .A3(new_n941), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n769), .A3(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n977), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n984), .B1(new_n1025), .B2(KEYINPUT115), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1024), .A2(new_n977), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n989), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n1019), .A2(new_n1029), .A3(new_n1015), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1018), .B1(new_n1030), .B2(KEYINPUT63), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1010), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1032), .A2(new_n992), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1007), .A2(new_n998), .A3(new_n703), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(G1981), .B2(G305), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1033), .B1(new_n996), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1031), .A2(new_n1036), .ZN(new_n1037));
  XOR2_X1   g612(.A(G299), .B(KEYINPUT57), .Z(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(G1956), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1040));
  XNOR2_X1  g615(.A(KEYINPUT56), .B(G2072), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NOR3_X1   g617(.A1(new_n976), .A2(new_n963), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1039), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1348), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n971), .B2(new_n973), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n940), .A2(new_n953), .A3(new_n993), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n613), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1044), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n964), .A2(new_n968), .A3(new_n1041), .ZN(new_n1051));
  AOI211_X1 g626(.A(KEYINPUT50), .B(G1384), .C1(new_n514), .C2(new_n517), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n761), .B1(new_n1052), .B2(new_n1021), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1053), .A3(new_n1038), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1050), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1038), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT61), .B1(new_n1056), .B2(KEYINPUT118), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1044), .A2(new_n1054), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1044), .A2(KEYINPUT118), .A3(KEYINPUT61), .A4(new_n1054), .ZN(new_n1060));
  AND2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G1996), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n964), .A2(new_n968), .A3(new_n1062), .ZN(new_n1063));
  XOR2_X1   g638(.A(KEYINPUT58), .B(G1341), .Z(new_n1064));
  NAND2_X1  g639(.A1(new_n994), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n994), .A2(KEYINPUT116), .A3(new_n1064), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1063), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n564), .ZN(new_n1070));
  NOR2_X1   g645(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1071));
  AND2_X1   g646(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1069), .A2(new_n564), .A3(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1046), .A2(new_n1047), .A3(KEYINPUT60), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n612), .A2(KEYINPUT119), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n612), .A2(KEYINPUT119), .ZN(new_n1078));
  OR3_X1    g653(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT60), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1080), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1073), .A2(new_n1075), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1055), .B1(new_n1061), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n1019), .B2(new_n1029), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1012), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n518), .A2(KEYINPUT45), .A3(new_n941), .ZN(new_n1087));
  AOI21_X1  g662(.A(G1966), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n971), .A2(new_n973), .A3(G2084), .ZN(new_n1089));
  OAI21_X1  g664(.A(G8), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n1091));
  NAND2_X1  g666(.A1(G286), .A2(G8), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1092), .B(KEYINPUT120), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1090), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1093), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT51), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1093), .B1(new_n1014), .B2(G8), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1095), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(G2078), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1086), .A2(new_n1087), .A3(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n797), .B1(new_n971), .B2(new_n973), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n976), .A2(new_n963), .A3(G2078), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1102), .B(new_n1103), .C1(new_n1104), .C2(KEYINPUT53), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(G171), .ZN(new_n1106));
  INV_X1    g681(.A(G2078), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n964), .A2(new_n968), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n1100), .ZN(new_n1109));
  INV_X1    g684(.A(new_n936), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n944), .A2(new_n1110), .A3(new_n962), .A4(new_n1101), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1109), .A2(G301), .A3(new_n1103), .A4(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT54), .B1(new_n1106), .B2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1099), .A2(new_n1113), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1052), .A2(new_n1021), .A3(G2090), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT115), .B1(new_n969), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1116), .A2(G8), .A3(new_n1028), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n990), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1118), .A2(KEYINPUT121), .A3(new_n992), .A4(new_n1010), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1103), .B(new_n1111), .C1(new_n1104), .C2(KEYINPUT53), .ZN(new_n1120));
  AOI21_X1  g695(.A(G301), .B1(new_n1120), .B2(KEYINPUT122), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1109), .A2(new_n1122), .A3(new_n1103), .A4(new_n1111), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  OR2_X1    g699(.A1(new_n1105), .A2(G171), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1124), .A2(KEYINPUT54), .A3(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1085), .A2(new_n1114), .A3(new_n1119), .A4(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1083), .B1(new_n1127), .B2(KEYINPUT123), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT54), .B1(new_n1105), .B2(G171), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1129), .B1(new_n1123), .B2(new_n1121), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1130), .A2(new_n1099), .A3(new_n1113), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1131), .A2(new_n1132), .A3(new_n1085), .A4(new_n1119), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1037), .B1(new_n1128), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1106), .B1(new_n1099), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1136), .A2(new_n1085), .A3(new_n1119), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT124), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1136), .A2(new_n1085), .A3(new_n1139), .A4(new_n1119), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1099), .A2(new_n1135), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1138), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n961), .B1(new_n1134), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n948), .B1(new_n955), .B2(new_n807), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT125), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n948), .A2(new_n1062), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT46), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT47), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n722), .A2(new_n725), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n957), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n946), .B1(new_n1151), .B2(new_n954), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n947), .B(KEYINPUT48), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1152), .B1(new_n960), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1149), .A2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT126), .B1(new_n1143), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1127), .A2(KEYINPUT123), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1083), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1157), .A2(new_n1133), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1037), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(new_n1142), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n961), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1155), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1156), .A2(new_n1166), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g742(.A1(G227), .A2(new_n458), .ZN(new_n1169));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n1170));
  NOR2_X1   g744(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  AND2_X1   g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1172));
  NOR4_X1   g746(.A1(G401), .A2(G229), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  NAND2_X1  g747(.A1(new_n866), .A2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g748(.A1(new_n914), .A2(new_n923), .ZN(new_n1175));
  NOR2_X1   g749(.A1(new_n1174), .A2(new_n1175), .ZN(G308));
  INV_X1    g750(.A(G308), .ZN(G225));
endmodule


