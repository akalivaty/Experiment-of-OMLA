

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(G164), .A2(G1384), .ZN(n794) );
  NOR2_X1 U556 ( .A1(n530), .A2(n529), .ZN(G164) );
  XNOR2_X2 U557 ( .A(KEYINPUT1), .B(n546), .ZN(n602) );
  XNOR2_X1 U558 ( .A(KEYINPUT97), .B(KEYINPUT31), .ZN(n727) );
  AND2_X1 U559 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U560 ( .A1(G2104), .A2(n525), .ZN(n887) );
  NOR2_X1 U561 ( .A1(G651), .A2(G543), .ZN(n647) );
  NOR2_X1 U562 ( .A1(n539), .A2(n538), .ZN(G160) );
  NAND2_X2 U563 ( .A1(n794), .A2(n690), .ZN(n730) );
  INV_X1 U564 ( .A(KEYINPUT29), .ZN(n712) );
  XNOR2_X1 U565 ( .A(n712), .B(KEYINPUT94), .ZN(n713) );
  XNOR2_X1 U566 ( .A(n714), .B(n713), .ZN(n718) );
  XNOR2_X1 U567 ( .A(n728), .B(n727), .ZN(n745) );
  INV_X1 U568 ( .A(n990), .ZN(n754) );
  INV_X1 U569 ( .A(KEYINPUT74), .ZN(n593) );
  XNOR2_X1 U570 ( .A(n593), .B(KEYINPUT13), .ZN(n594) );
  XNOR2_X1 U571 ( .A(n595), .B(n594), .ZN(n596) );
  NOR2_X1 U572 ( .A1(n644), .A2(n544), .ZN(n651) );
  AND2_X1 U573 ( .A1(G2105), .A2(G2104), .ZN(n889) );
  NAND2_X1 U574 ( .A1(G114), .A2(n889), .ZN(n521) );
  INV_X1 U575 ( .A(G2105), .ZN(n525) );
  NAND2_X1 U576 ( .A1(G126), .A2(n887), .ZN(n520) );
  NAND2_X1 U577 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U578 ( .A(KEYINPUT88), .B(n522), .ZN(n530) );
  NOR2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  XOR2_X1 U580 ( .A(KEYINPUT17), .B(n523), .Z(n524) );
  XNOR2_X1 U581 ( .A(KEYINPUT66), .B(n524), .ZN(n623) );
  NAND2_X1 U582 ( .A1(G138), .A2(n623), .ZN(n527) );
  AND2_X2 U583 ( .A1(n525), .A2(G2104), .ZN(n895) );
  NAND2_X1 U584 ( .A1(n895), .A2(G102), .ZN(n526) );
  NAND2_X1 U585 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U586 ( .A(n528), .B(KEYINPUT89), .Z(n529) );
  NAND2_X1 U587 ( .A1(G113), .A2(n889), .ZN(n532) );
  NAND2_X1 U588 ( .A1(G137), .A2(n623), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n532), .A2(n531), .ZN(n539) );
  INV_X1 U590 ( .A(KEYINPUT65), .ZN(n537) );
  NAND2_X1 U591 ( .A1(n895), .A2(G101), .ZN(n533) );
  XOR2_X1 U592 ( .A(KEYINPUT23), .B(n533), .Z(n535) );
  NAND2_X1 U593 ( .A1(n887), .A2(G125), .ZN(n534) );
  NAND2_X1 U594 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U595 ( .A(n537), .B(n536), .ZN(n538) );
  NAND2_X1 U596 ( .A1(G90), .A2(n647), .ZN(n542) );
  XNOR2_X1 U597 ( .A(G543), .B(KEYINPUT0), .ZN(n540) );
  XNOR2_X1 U598 ( .A(n540), .B(KEYINPUT67), .ZN(n644) );
  XOR2_X1 U599 ( .A(KEYINPUT68), .B(G651), .Z(n544) );
  NAND2_X1 U600 ( .A1(G77), .A2(n651), .ZN(n541) );
  NAND2_X1 U601 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U602 ( .A(KEYINPUT9), .B(n543), .ZN(n550) );
  NOR2_X1 U603 ( .A1(G543), .A2(n544), .ZN(n545) );
  XNOR2_X1 U604 ( .A(n545), .B(KEYINPUT69), .ZN(n546) );
  NAND2_X1 U605 ( .A1(n602), .A2(G64), .ZN(n548) );
  NOR2_X2 U606 ( .A1(G651), .A2(n644), .ZN(n648) );
  NAND2_X1 U607 ( .A1(n648), .A2(G52), .ZN(n547) );
  AND2_X1 U608 ( .A1(n548), .A2(n547), .ZN(n549) );
  NAND2_X1 U609 ( .A1(n550), .A2(n549), .ZN(G301) );
  INV_X1 U610 ( .A(G301), .ZN(G171) );
  NAND2_X1 U611 ( .A1(n648), .A2(G47), .ZN(n552) );
  NAND2_X1 U612 ( .A1(G60), .A2(n602), .ZN(n551) );
  NAND2_X1 U613 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U614 ( .A1(G85), .A2(n647), .ZN(n554) );
  NAND2_X1 U615 ( .A1(G72), .A2(n651), .ZN(n553) );
  NAND2_X1 U616 ( .A1(n554), .A2(n553), .ZN(n555) );
  OR2_X1 U617 ( .A1(n556), .A2(n555), .ZN(G290) );
  AND2_X1 U618 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U619 ( .A(G132), .ZN(G219) );
  INV_X1 U620 ( .A(G82), .ZN(G220) );
  INV_X1 U621 ( .A(G57), .ZN(G237) );
  INV_X1 U622 ( .A(G120), .ZN(G236) );
  NAND2_X1 U623 ( .A1(G88), .A2(n647), .ZN(n558) );
  NAND2_X1 U624 ( .A1(G75), .A2(n651), .ZN(n557) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U626 ( .A1(n648), .A2(G50), .ZN(n560) );
  NAND2_X1 U627 ( .A1(G62), .A2(n602), .ZN(n559) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U629 ( .A1(n562), .A2(n561), .ZN(G166) );
  NAND2_X1 U630 ( .A1(n648), .A2(G53), .ZN(n563) );
  XOR2_X1 U631 ( .A(KEYINPUT71), .B(n563), .Z(n565) );
  NAND2_X1 U632 ( .A1(G65), .A2(n602), .ZN(n564) );
  NAND2_X1 U633 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U634 ( .A(KEYINPUT72), .B(n566), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n647), .A2(G91), .ZN(n567) );
  XOR2_X1 U636 ( .A(KEYINPUT70), .B(n567), .Z(n568) );
  NOR2_X1 U637 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U638 ( .A1(G78), .A2(n651), .ZN(n570) );
  NAND2_X1 U639 ( .A1(n571), .A2(n570), .ZN(G299) );
  NAND2_X1 U640 ( .A1(n647), .A2(G89), .ZN(n572) );
  XNOR2_X1 U641 ( .A(KEYINPUT4), .B(n572), .ZN(n575) );
  NAND2_X1 U642 ( .A1(G76), .A2(n651), .ZN(n573) );
  XOR2_X1 U643 ( .A(KEYINPUT77), .B(n573), .Z(n574) );
  NAND2_X1 U644 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U645 ( .A(n576), .B(KEYINPUT5), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n648), .A2(G51), .ZN(n577) );
  XNOR2_X1 U647 ( .A(n577), .B(KEYINPUT78), .ZN(n579) );
  NAND2_X1 U648 ( .A1(G63), .A2(n602), .ZN(n578) );
  NAND2_X1 U649 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U650 ( .A(KEYINPUT6), .B(n580), .Z(n581) );
  NAND2_X1 U651 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U652 ( .A(n583), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U653 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U654 ( .A1(G7), .A2(G661), .ZN(n584) );
  XNOR2_X1 U655 ( .A(n584), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U656 ( .A(G223), .ZN(n833) );
  NAND2_X1 U657 ( .A1(n833), .A2(G567), .ZN(n585) );
  XNOR2_X1 U658 ( .A(n585), .B(KEYINPUT11), .ZN(n586) );
  XNOR2_X1 U659 ( .A(KEYINPUT73), .B(n586), .ZN(G234) );
  NAND2_X1 U660 ( .A1(G56), .A2(n602), .ZN(n587) );
  XNOR2_X1 U661 ( .A(n587), .B(KEYINPUT14), .ZN(n589) );
  NAND2_X1 U662 ( .A1(G43), .A2(n648), .ZN(n588) );
  NAND2_X1 U663 ( .A1(n589), .A2(n588), .ZN(n597) );
  NAND2_X1 U664 ( .A1(n647), .A2(G81), .ZN(n590) );
  XNOR2_X1 U665 ( .A(n590), .B(KEYINPUT12), .ZN(n592) );
  NAND2_X1 U666 ( .A1(G68), .A2(n651), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n592), .A2(n591), .ZN(n595) );
  NOR2_X1 U668 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U669 ( .A(KEYINPUT75), .B(n598), .ZN(n984) );
  INV_X1 U670 ( .A(n984), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n599), .A2(G860), .ZN(G153) );
  NAND2_X1 U672 ( .A1(G868), .A2(G301), .ZN(n610) );
  NAND2_X1 U673 ( .A1(n648), .A2(G54), .ZN(n601) );
  NAND2_X1 U674 ( .A1(G79), .A2(n651), .ZN(n600) );
  NAND2_X1 U675 ( .A1(n601), .A2(n600), .ZN(n607) );
  NAND2_X1 U676 ( .A1(n647), .A2(G92), .ZN(n604) );
  NAND2_X1 U677 ( .A1(G66), .A2(n602), .ZN(n603) );
  NAND2_X1 U678 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U679 ( .A(KEYINPUT76), .B(n605), .ZN(n606) );
  NOR2_X1 U680 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U681 ( .A(n608), .B(KEYINPUT15), .ZN(n696) );
  INV_X1 U682 ( .A(G868), .ZN(n669) );
  NAND2_X1 U683 ( .A1(n696), .A2(n669), .ZN(n609) );
  NAND2_X1 U684 ( .A1(n610), .A2(n609), .ZN(G284) );
  NOR2_X1 U685 ( .A1(G868), .A2(G299), .ZN(n611) );
  XOR2_X1 U686 ( .A(KEYINPUT79), .B(n611), .Z(n613) );
  NOR2_X1 U687 ( .A1(G286), .A2(n669), .ZN(n612) );
  NOR2_X1 U688 ( .A1(n613), .A2(n612), .ZN(G297) );
  INV_X1 U689 ( .A(G559), .ZN(n616) );
  NOR2_X1 U690 ( .A1(G860), .A2(n616), .ZN(n614) );
  NOR2_X1 U691 ( .A1(n696), .A2(n614), .ZN(n615) );
  XOR2_X1 U692 ( .A(KEYINPUT16), .B(n615), .Z(G148) );
  INV_X1 U693 ( .A(n696), .ZN(n976) );
  NAND2_X1 U694 ( .A1(n616), .A2(n976), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n617), .A2(G868), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n984), .A2(n669), .ZN(n618) );
  NAND2_X1 U697 ( .A1(n619), .A2(n618), .ZN(G282) );
  NAND2_X1 U698 ( .A1(n887), .A2(G123), .ZN(n620) );
  XNOR2_X1 U699 ( .A(n620), .B(KEYINPUT18), .ZN(n622) );
  NAND2_X1 U700 ( .A1(G99), .A2(n895), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n622), .A2(n621), .ZN(n627) );
  NAND2_X1 U702 ( .A1(G111), .A2(n889), .ZN(n625) );
  BUF_X1 U703 ( .A(n623), .Z(n893) );
  NAND2_X1 U704 ( .A1(G135), .A2(n893), .ZN(n624) );
  NAND2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U706 ( .A1(n627), .A2(n626), .ZN(n932) );
  XNOR2_X1 U707 ( .A(G2096), .B(n932), .ZN(n629) );
  INV_X1 U708 ( .A(G2100), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(G156) );
  NAND2_X1 U710 ( .A1(G559), .A2(n976), .ZN(n630) );
  XNOR2_X1 U711 ( .A(n630), .B(KEYINPUT80), .ZN(n667) );
  XNOR2_X1 U712 ( .A(n667), .B(n984), .ZN(n631) );
  NOR2_X1 U713 ( .A1(n631), .A2(G860), .ZN(n639) );
  NAND2_X1 U714 ( .A1(G93), .A2(n647), .ZN(n633) );
  NAND2_X1 U715 ( .A1(G80), .A2(n651), .ZN(n632) );
  NAND2_X1 U716 ( .A1(n633), .A2(n632), .ZN(n638) );
  NAND2_X1 U717 ( .A1(n648), .A2(G55), .ZN(n635) );
  NAND2_X1 U718 ( .A1(G67), .A2(n602), .ZN(n634) );
  NAND2_X1 U719 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U720 ( .A(KEYINPUT81), .B(n636), .Z(n637) );
  OR2_X1 U721 ( .A1(n638), .A2(n637), .ZN(n670) );
  XOR2_X1 U722 ( .A(n639), .B(n670), .Z(G145) );
  NAND2_X1 U723 ( .A1(G49), .A2(n648), .ZN(n641) );
  NAND2_X1 U724 ( .A1(G74), .A2(G651), .ZN(n640) );
  NAND2_X1 U725 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U726 ( .A(KEYINPUT82), .B(n642), .ZN(n643) );
  NOR2_X1 U727 ( .A1(n602), .A2(n643), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n644), .A2(G87), .ZN(n645) );
  NAND2_X1 U729 ( .A1(n646), .A2(n645), .ZN(G288) );
  NAND2_X1 U730 ( .A1(G86), .A2(n647), .ZN(n650) );
  NAND2_X1 U731 ( .A1(G48), .A2(n648), .ZN(n649) );
  NAND2_X1 U732 ( .A1(n650), .A2(n649), .ZN(n655) );
  NAND2_X1 U733 ( .A1(n651), .A2(G73), .ZN(n652) );
  XNOR2_X1 U734 ( .A(n652), .B(KEYINPUT2), .ZN(n653) );
  XNOR2_X1 U735 ( .A(n653), .B(KEYINPUT83), .ZN(n654) );
  NOR2_X1 U736 ( .A1(n655), .A2(n654), .ZN(n657) );
  NAND2_X1 U737 ( .A1(G61), .A2(n602), .ZN(n656) );
  NAND2_X1 U738 ( .A1(n657), .A2(n656), .ZN(G305) );
  XOR2_X1 U739 ( .A(KEYINPUT84), .B(KEYINPUT86), .Z(n659) );
  XNOR2_X1 U740 ( .A(KEYINPUT85), .B(KEYINPUT19), .ZN(n658) );
  XNOR2_X1 U741 ( .A(n659), .B(n658), .ZN(n662) );
  XNOR2_X1 U742 ( .A(G166), .B(G290), .ZN(n660) );
  XNOR2_X1 U743 ( .A(n660), .B(G288), .ZN(n661) );
  XNOR2_X1 U744 ( .A(n662), .B(n661), .ZN(n664) );
  XOR2_X1 U745 ( .A(G305), .B(n670), .Z(n663) );
  XNOR2_X1 U746 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U747 ( .A(n665), .B(n984), .ZN(n666) );
  XNOR2_X1 U748 ( .A(n666), .B(G299), .ZN(n906) );
  XOR2_X1 U749 ( .A(n906), .B(n667), .Z(n668) );
  NOR2_X1 U750 ( .A1(n669), .A2(n668), .ZN(n672) );
  NOR2_X1 U751 ( .A1(G868), .A2(n670), .ZN(n671) );
  NOR2_X1 U752 ( .A1(n672), .A2(n671), .ZN(G295) );
  NAND2_X1 U753 ( .A1(G2084), .A2(G2078), .ZN(n673) );
  XOR2_X1 U754 ( .A(KEYINPUT20), .B(n673), .Z(n674) );
  NAND2_X1 U755 ( .A1(G2090), .A2(n674), .ZN(n675) );
  XNOR2_X1 U756 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U757 ( .A1(n676), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U759 ( .A1(G236), .A2(G237), .ZN(n677) );
  NAND2_X1 U760 ( .A1(G69), .A2(n677), .ZN(n678) );
  XNOR2_X1 U761 ( .A(KEYINPUT87), .B(n678), .ZN(n679) );
  NAND2_X1 U762 ( .A1(n679), .A2(G108), .ZN(n839) );
  NAND2_X1 U763 ( .A1(n839), .A2(G567), .ZN(n684) );
  NOR2_X1 U764 ( .A1(G220), .A2(G219), .ZN(n680) );
  XOR2_X1 U765 ( .A(KEYINPUT22), .B(n680), .Z(n681) );
  NOR2_X1 U766 ( .A1(G218), .A2(n681), .ZN(n682) );
  NAND2_X1 U767 ( .A1(G96), .A2(n682), .ZN(n840) );
  NAND2_X1 U768 ( .A1(n840), .A2(G2106), .ZN(n683) );
  NAND2_X1 U769 ( .A1(n684), .A2(n683), .ZN(n841) );
  NAND2_X1 U770 ( .A1(G483), .A2(G661), .ZN(n685) );
  NOR2_X1 U771 ( .A1(n841), .A2(n685), .ZN(n838) );
  NAND2_X1 U772 ( .A1(n838), .A2(G36), .ZN(G176) );
  INV_X1 U773 ( .A(G166), .ZN(G303) );
  NAND2_X1 U774 ( .A1(G160), .A2(G40), .ZN(n793) );
  INV_X1 U775 ( .A(n793), .ZN(n690) );
  INV_X1 U776 ( .A(G1996), .ZN(n860) );
  NOR2_X1 U777 ( .A1(n730), .A2(n860), .ZN(n686) );
  XNOR2_X1 U778 ( .A(n686), .B(KEYINPUT26), .ZN(n688) );
  AND2_X1 U779 ( .A1(n730), .A2(G1341), .ZN(n687) );
  OR2_X1 U780 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U781 ( .A1(n689), .A2(n984), .ZN(n694) );
  NAND2_X1 U782 ( .A1(G1348), .A2(n730), .ZN(n692) );
  AND2_X1 U783 ( .A1(n690), .A2(n794), .ZN(n699) );
  NAND2_X1 U784 ( .A1(n699), .A2(G2067), .ZN(n691) );
  NAND2_X1 U785 ( .A1(n692), .A2(n691), .ZN(n695) );
  NOR2_X1 U786 ( .A1(n696), .A2(n695), .ZN(n693) );
  NOR2_X1 U787 ( .A1(n694), .A2(n693), .ZN(n698) );
  AND2_X1 U788 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U789 ( .A1(n698), .A2(n697), .ZN(n705) );
  NAND2_X1 U790 ( .A1(n699), .A2(G2072), .ZN(n700) );
  XOR2_X1 U791 ( .A(n700), .B(KEYINPUT27), .Z(n707) );
  NAND2_X1 U792 ( .A1(G1956), .A2(n730), .ZN(n706) );
  INV_X1 U793 ( .A(G299), .ZN(n701) );
  AND2_X1 U794 ( .A1(n706), .A2(n701), .ZN(n702) );
  AND2_X1 U795 ( .A1(n707), .A2(n702), .ZN(n703) );
  XOR2_X1 U796 ( .A(n703), .B(KEYINPUT93), .Z(n704) );
  NOR2_X1 U797 ( .A1(n705), .A2(n704), .ZN(n711) );
  NAND2_X1 U798 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U799 ( .A1(G299), .A2(n708), .ZN(n709) );
  XOR2_X1 U800 ( .A(KEYINPUT28), .B(n709), .Z(n710) );
  NOR2_X1 U801 ( .A1(n711), .A2(n710), .ZN(n714) );
  XNOR2_X1 U802 ( .A(G2078), .B(KEYINPUT25), .ZN(n964) );
  NOR2_X1 U803 ( .A1(n730), .A2(n964), .ZN(n716) );
  AND2_X1 U804 ( .A1(n730), .A2(G1961), .ZN(n715) );
  NOR2_X1 U805 ( .A1(n716), .A2(n715), .ZN(n720) );
  AND2_X1 U806 ( .A1(G171), .A2(n720), .ZN(n717) );
  NOR2_X1 U807 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U808 ( .A(n719), .B(KEYINPUT95), .ZN(n744) );
  NOR2_X1 U809 ( .A1(G171), .A2(n720), .ZN(n726) );
  NAND2_X1 U810 ( .A1(G8), .A2(n730), .ZN(n808) );
  NOR2_X1 U811 ( .A1(G1966), .A2(n808), .ZN(n747) );
  NOR2_X1 U812 ( .A1(G2084), .A2(n730), .ZN(n743) );
  NOR2_X1 U813 ( .A1(n747), .A2(n743), .ZN(n721) );
  XNOR2_X1 U814 ( .A(n721), .B(KEYINPUT96), .ZN(n722) );
  NAND2_X1 U815 ( .A1(n722), .A2(G8), .ZN(n723) );
  XNOR2_X1 U816 ( .A(KEYINPUT30), .B(n723), .ZN(n724) );
  NOR2_X1 U817 ( .A1(G168), .A2(n724), .ZN(n725) );
  NOR2_X1 U818 ( .A1(n726), .A2(n725), .ZN(n728) );
  INV_X1 U819 ( .A(G8), .ZN(n735) );
  NOR2_X1 U820 ( .A1(G1971), .A2(n808), .ZN(n729) );
  XNOR2_X1 U821 ( .A(n729), .B(KEYINPUT98), .ZN(n732) );
  NOR2_X1 U822 ( .A1(n730), .A2(G2090), .ZN(n731) );
  NOR2_X1 U823 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U824 ( .A1(n733), .A2(G303), .ZN(n734) );
  OR2_X1 U825 ( .A1(n735), .A2(n734), .ZN(n737) );
  AND2_X1 U826 ( .A1(n745), .A2(n737), .ZN(n736) );
  NAND2_X1 U827 ( .A1(n744), .A2(n736), .ZN(n740) );
  INV_X1 U828 ( .A(n737), .ZN(n738) );
  OR2_X1 U829 ( .A1(n738), .A2(G286), .ZN(n739) );
  NAND2_X1 U830 ( .A1(n740), .A2(n739), .ZN(n742) );
  XOR2_X1 U831 ( .A(KEYINPUT32), .B(KEYINPUT99), .Z(n741) );
  XNOR2_X1 U832 ( .A(n742), .B(n741), .ZN(n751) );
  NAND2_X1 U833 ( .A1(G8), .A2(n743), .ZN(n749) );
  AND2_X1 U834 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U836 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n751), .A2(n750), .ZN(n800) );
  NOR2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n759) );
  NOR2_X1 U839 ( .A1(G1971), .A2(G303), .ZN(n752) );
  NOR2_X1 U840 ( .A1(n759), .A2(n752), .ZN(n753) );
  NAND2_X1 U841 ( .A1(n800), .A2(n753), .ZN(n756) );
  NAND2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n990) );
  NOR2_X1 U843 ( .A1(n808), .A2(n754), .ZN(n755) );
  XNOR2_X1 U844 ( .A(KEYINPUT64), .B(n757), .ZN(n758) );
  NOR2_X1 U845 ( .A1(n758), .A2(KEYINPUT33), .ZN(n799) );
  XNOR2_X1 U846 ( .A(G1981), .B(G305), .ZN(n980) );
  INV_X1 U847 ( .A(n980), .ZN(n764) );
  INV_X1 U848 ( .A(KEYINPUT33), .ZN(n761) );
  INV_X1 U849 ( .A(n759), .ZN(n989) );
  OR2_X1 U850 ( .A1(n808), .A2(n989), .ZN(n760) );
  NOR2_X1 U851 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U852 ( .A(n762), .B(KEYINPUT100), .Z(n763) );
  NAND2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n797) );
  XOR2_X1 U854 ( .A(G1986), .B(G290), .Z(n988) );
  XNOR2_X1 U855 ( .A(G2067), .B(KEYINPUT37), .ZN(n765) );
  XOR2_X1 U856 ( .A(n765), .B(KEYINPUT90), .Z(n824) );
  NAND2_X1 U857 ( .A1(n895), .A2(G104), .ZN(n767) );
  NAND2_X1 U858 ( .A1(G140), .A2(n893), .ZN(n766) );
  NAND2_X1 U859 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U860 ( .A(KEYINPUT34), .B(n768), .ZN(n774) );
  NAND2_X1 U861 ( .A1(n889), .A2(G116), .ZN(n769) );
  XOR2_X1 U862 ( .A(KEYINPUT91), .B(n769), .Z(n771) );
  NAND2_X1 U863 ( .A1(n887), .A2(G128), .ZN(n770) );
  NAND2_X1 U864 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U865 ( .A(KEYINPUT35), .B(n772), .Z(n773) );
  NOR2_X1 U866 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U867 ( .A(KEYINPUT36), .B(n775), .Z(n903) );
  NAND2_X1 U868 ( .A1(n824), .A2(n903), .ZN(n822) );
  INV_X1 U869 ( .A(n822), .ZN(n792) );
  NAND2_X1 U870 ( .A1(G129), .A2(n887), .ZN(n777) );
  NAND2_X1 U871 ( .A1(G141), .A2(n893), .ZN(n776) );
  NAND2_X1 U872 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U873 ( .A1(n895), .A2(G105), .ZN(n778) );
  XOR2_X1 U874 ( .A(KEYINPUT38), .B(n778), .Z(n779) );
  NOR2_X1 U875 ( .A1(n780), .A2(n779), .ZN(n782) );
  NAND2_X1 U876 ( .A1(n889), .A2(G117), .ZN(n781) );
  NAND2_X1 U877 ( .A1(n782), .A2(n781), .ZN(n873) );
  NAND2_X1 U878 ( .A1(n873), .A2(G1996), .ZN(n790) );
  NAND2_X1 U879 ( .A1(G119), .A2(n887), .ZN(n784) );
  NAND2_X1 U880 ( .A1(G131), .A2(n893), .ZN(n783) );
  NAND2_X1 U881 ( .A1(n784), .A2(n783), .ZN(n788) );
  NAND2_X1 U882 ( .A1(G107), .A2(n889), .ZN(n786) );
  NAND2_X1 U883 ( .A1(G95), .A2(n895), .ZN(n785) );
  NAND2_X1 U884 ( .A1(n786), .A2(n785), .ZN(n787) );
  OR2_X1 U885 ( .A1(n788), .A2(n787), .ZN(n869) );
  NAND2_X1 U886 ( .A1(G1991), .A2(n869), .ZN(n789) );
  NAND2_X1 U887 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U888 ( .A(n791), .B(KEYINPUT92), .ZN(n818) );
  NOR2_X1 U889 ( .A1(n792), .A2(n818), .ZN(n939) );
  NAND2_X1 U890 ( .A1(n988), .A2(n939), .ZN(n795) );
  NOR2_X1 U891 ( .A1(n794), .A2(n793), .ZN(n827) );
  NAND2_X1 U892 ( .A1(n795), .A2(n827), .ZN(n812) );
  INV_X1 U893 ( .A(n812), .ZN(n796) );
  OR2_X1 U894 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U895 ( .A1(n799), .A2(n798), .ZN(n814) );
  INV_X1 U896 ( .A(n800), .ZN(n803) );
  NAND2_X1 U897 ( .A1(G166), .A2(G8), .ZN(n801) );
  NOR2_X1 U898 ( .A1(G2090), .A2(n801), .ZN(n802) );
  NOR2_X1 U899 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U900 ( .A(n804), .B(KEYINPUT101), .ZN(n805) );
  NAND2_X1 U901 ( .A1(n805), .A2(n808), .ZN(n810) );
  NOR2_X1 U902 ( .A1(G1981), .A2(G305), .ZN(n806) );
  XOR2_X1 U903 ( .A(n806), .B(KEYINPUT24), .Z(n807) );
  OR2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n809) );
  NAND2_X1 U905 ( .A1(n810), .A2(n809), .ZN(n811) );
  AND2_X1 U906 ( .A1(n812), .A2(n811), .ZN(n813) );
  NOR2_X1 U907 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U908 ( .A(n815), .B(KEYINPUT102), .ZN(n830) );
  NOR2_X1 U909 ( .A1(G1996), .A2(n873), .ZN(n930) );
  NOR2_X1 U910 ( .A1(G1986), .A2(G290), .ZN(n816) );
  NOR2_X1 U911 ( .A1(G1991), .A2(n869), .ZN(n933) );
  NOR2_X1 U912 ( .A1(n816), .A2(n933), .ZN(n817) );
  NOR2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U914 ( .A1(n930), .A2(n819), .ZN(n820) );
  XOR2_X1 U915 ( .A(n820), .B(KEYINPUT103), .Z(n821) );
  XNOR2_X1 U916 ( .A(KEYINPUT39), .B(n821), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n826) );
  NOR2_X1 U918 ( .A1(n903), .A2(n824), .ZN(n825) );
  XOR2_X1 U919 ( .A(KEYINPUT104), .B(n825), .Z(n941) );
  NAND2_X1 U920 ( .A1(n826), .A2(n941), .ZN(n828) );
  NAND2_X1 U921 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U922 ( .A1(n830), .A2(n829), .ZN(n832) );
  XOR2_X1 U923 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n831) );
  XNOR2_X1 U924 ( .A(n832), .B(n831), .ZN(G329) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n833), .ZN(G217) );
  NAND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n835) );
  INV_X1 U927 ( .A(G661), .ZN(n834) );
  NOR2_X1 U928 ( .A1(n835), .A2(n834), .ZN(n836) );
  XNOR2_X1 U929 ( .A(n836), .B(KEYINPUT109), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U931 ( .A1(n838), .A2(n837), .ZN(G188) );
  XOR2_X1 U932 ( .A(G108), .B(KEYINPUT118), .Z(G238) );
  INV_X1 U934 ( .A(G96), .ZN(G221) );
  NOR2_X1 U935 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  INV_X1 U937 ( .A(n841), .ZN(G319) );
  XOR2_X1 U938 ( .A(G2096), .B(G2678), .Z(n843) );
  XNOR2_X1 U939 ( .A(G2072), .B(KEYINPUT43), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U941 ( .A(n844), .B(KEYINPUT42), .Z(n846) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2090), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U944 ( .A(KEYINPUT110), .B(G2100), .Z(n848) );
  XNOR2_X1 U945 ( .A(G2084), .B(G2078), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(G227) );
  XOR2_X1 U948 ( .A(G1981), .B(G1961), .Z(n852) );
  XNOR2_X1 U949 ( .A(G1991), .B(G1966), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n856) );
  XOR2_X1 U951 ( .A(G1976), .B(G1971), .Z(n854) );
  XNOR2_X1 U952 ( .A(G1986), .B(G1956), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U954 ( .A(n856), .B(n855), .Z(n858) );
  XNOR2_X1 U955 ( .A(G2474), .B(KEYINPUT111), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U957 ( .A(KEYINPUT41), .B(n859), .ZN(n861) );
  XNOR2_X1 U958 ( .A(n861), .B(n860), .ZN(G229) );
  NAND2_X1 U959 ( .A1(n887), .A2(G124), .ZN(n862) );
  XNOR2_X1 U960 ( .A(n862), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U961 ( .A1(G100), .A2(n895), .ZN(n863) );
  NAND2_X1 U962 ( .A1(n864), .A2(n863), .ZN(n868) );
  NAND2_X1 U963 ( .A1(G112), .A2(n889), .ZN(n866) );
  NAND2_X1 U964 ( .A1(G136), .A2(n893), .ZN(n865) );
  NAND2_X1 U965 ( .A1(n866), .A2(n865), .ZN(n867) );
  NOR2_X1 U966 ( .A1(n868), .A2(n867), .ZN(G162) );
  XNOR2_X1 U967 ( .A(KEYINPUT115), .B(KEYINPUT46), .ZN(n871) );
  XNOR2_X1 U968 ( .A(n869), .B(KEYINPUT48), .ZN(n870) );
  XNOR2_X1 U969 ( .A(n871), .B(n870), .ZN(n872) );
  XNOR2_X1 U970 ( .A(n932), .B(n872), .ZN(n875) );
  XNOR2_X1 U971 ( .A(n873), .B(G164), .ZN(n874) );
  XNOR2_X1 U972 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U973 ( .A(n876), .B(G162), .Z(n886) );
  NAND2_X1 U974 ( .A1(G115), .A2(n889), .ZN(n878) );
  NAND2_X1 U975 ( .A1(G127), .A2(n887), .ZN(n877) );
  NAND2_X1 U976 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U977 ( .A(n879), .B(KEYINPUT47), .ZN(n881) );
  NAND2_X1 U978 ( .A1(G139), .A2(n893), .ZN(n880) );
  NAND2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n884) );
  NAND2_X1 U980 ( .A1(n895), .A2(G103), .ZN(n882) );
  XOR2_X1 U981 ( .A(KEYINPUT116), .B(n882), .Z(n883) );
  NOR2_X1 U982 ( .A1(n884), .A2(n883), .ZN(n943) );
  XNOR2_X1 U983 ( .A(G160), .B(n943), .ZN(n885) );
  XNOR2_X1 U984 ( .A(n886), .B(n885), .ZN(n902) );
  NAND2_X1 U985 ( .A1(n887), .A2(G130), .ZN(n888) );
  XNOR2_X1 U986 ( .A(n888), .B(KEYINPUT112), .ZN(n891) );
  NAND2_X1 U987 ( .A1(G118), .A2(n889), .ZN(n890) );
  NAND2_X1 U988 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U989 ( .A(KEYINPUT113), .B(n892), .Z(n900) );
  NAND2_X1 U990 ( .A1(G142), .A2(n893), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n894), .B(KEYINPUT114), .ZN(n897) );
  NAND2_X1 U992 ( .A1(G106), .A2(n895), .ZN(n896) );
  NAND2_X1 U993 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U994 ( .A(n898), .B(KEYINPUT45), .Z(n899) );
  NOR2_X1 U995 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U996 ( .A(n902), .B(n901), .Z(n904) );
  XNOR2_X1 U997 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U998 ( .A1(G37), .A2(n905), .ZN(G395) );
  XNOR2_X1 U999 ( .A(n976), .B(G286), .ZN(n907) );
  XNOR2_X1 U1000 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1001 ( .A(n908), .B(G171), .ZN(n909) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n909), .ZN(G397) );
  XOR2_X1 U1003 ( .A(G2451), .B(KEYINPUT108), .Z(n911) );
  XNOR2_X1 U1004 ( .A(G2443), .B(G2446), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(n911), .B(n910), .ZN(n915) );
  XOR2_X1 U1006 ( .A(G2435), .B(G2438), .Z(n913) );
  XNOR2_X1 U1007 ( .A(G2454), .B(G2430), .ZN(n912) );
  XNOR2_X1 U1008 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1009 ( .A(n915), .B(n914), .Z(n917) );
  XNOR2_X1 U1010 ( .A(G2427), .B(KEYINPUT106), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(n917), .B(n916), .ZN(n920) );
  XOR2_X1 U1012 ( .A(G1341), .B(G1348), .Z(n918) );
  XNOR2_X1 U1013 ( .A(KEYINPUT107), .B(n918), .ZN(n919) );
  XOR2_X1 U1014 ( .A(n920), .B(n919), .Z(n921) );
  NAND2_X1 U1015 ( .A1(G14), .A2(n921), .ZN(n928) );
  NAND2_X1 U1016 ( .A1(G319), .A2(n928), .ZN(n925) );
  NOR2_X1 U1017 ( .A1(G227), .A2(G229), .ZN(n922) );
  XOR2_X1 U1018 ( .A(KEYINPUT49), .B(n922), .Z(n923) );
  XNOR2_X1 U1019 ( .A(n923), .B(KEYINPUT117), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(n925), .A2(n924), .ZN(n927) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n926) );
  NAND2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(G225) );
  INV_X1 U1023 ( .A(G225), .ZN(G308) );
  INV_X1 U1024 ( .A(G69), .ZN(G235) );
  INV_X1 U1025 ( .A(n928), .ZN(G401) );
  XOR2_X1 U1026 ( .A(G2090), .B(G162), .Z(n929) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1028 ( .A(KEYINPUT51), .B(n931), .Z(n935) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n937) );
  XOR2_X1 U1031 ( .A(G160), .B(G2084), .Z(n936) );
  NOR2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1034 ( .A(KEYINPUT119), .B(n940), .ZN(n942) );
  NAND2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n948) );
  XOR2_X1 U1036 ( .A(G2072), .B(n943), .Z(n945) );
  XOR2_X1 U1037 ( .A(G164), .B(G2078), .Z(n944) );
  NOR2_X1 U1038 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1039 ( .A(KEYINPUT50), .B(n946), .Z(n947) );
  NOR2_X1 U1040 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1041 ( .A(KEYINPUT52), .B(n949), .ZN(n951) );
  INV_X1 U1042 ( .A(KEYINPUT55), .ZN(n950) );
  NAND2_X1 U1043 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1044 ( .A1(n952), .A2(G29), .ZN(n1030) );
  XNOR2_X1 U1045 ( .A(G29), .B(KEYINPUT123), .ZN(n974) );
  XOR2_X1 U1046 ( .A(G2090), .B(G35), .Z(n956) );
  XNOR2_X1 U1047 ( .A(KEYINPUT54), .B(KEYINPUT121), .ZN(n953) );
  XNOR2_X1 U1048 ( .A(n953), .B(G34), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(n954), .B(G2084), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n970) );
  XNOR2_X1 U1051 ( .A(G1996), .B(G32), .ZN(n958) );
  XNOR2_X1 U1052 ( .A(G33), .B(G2072), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n963) );
  XOR2_X1 U1054 ( .A(G1991), .B(G25), .Z(n959) );
  NAND2_X1 U1055 ( .A1(n959), .A2(G28), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(G26), .B(G2067), .ZN(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n966) );
  XOR2_X1 U1059 ( .A(G27), .B(n964), .Z(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(KEYINPUT120), .B(n967), .ZN(n968) );
  XNOR2_X1 U1062 ( .A(KEYINPUT53), .B(n968), .ZN(n969) );
  NOR2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(KEYINPUT55), .B(n971), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(n972), .B(KEYINPUT122), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1067 ( .A1(n975), .A2(G11), .ZN(n1028) );
  XNOR2_X1 U1068 ( .A(G16), .B(KEYINPUT56), .ZN(n1000) );
  XNOR2_X1 U1069 ( .A(n976), .B(G1348), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(G171), .B(G1961), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n983) );
  XOR2_X1 U1072 ( .A(G1966), .B(G168), .Z(n979) );
  NOR2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(n981), .B(KEYINPUT57), .ZN(n982) );
  NOR2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n998) );
  XNOR2_X1 U1076 ( .A(n984), .B(G1341), .ZN(n996) );
  XNOR2_X1 U1077 ( .A(G299), .B(G1956), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(G303), .B(G1971), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n993) );
  NAND2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(KEYINPUT124), .B(n991), .ZN(n992) );
  NOR2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(KEYINPUT125), .B(n994), .ZN(n995) );
  NOR2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1026) );
  INV_X1 U1088 ( .A(G16), .ZN(n1024) );
  XNOR2_X1 U1089 ( .A(G1961), .B(G5), .ZN(n1001) );
  XNOR2_X1 U1090 ( .A(n1001), .B(KEYINPUT126), .ZN(n1008) );
  XNOR2_X1 U1091 ( .A(G1971), .B(G22), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(G23), .B(G1976), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  XOR2_X1 U1094 ( .A(G1986), .B(G24), .Z(n1004) );
  NAND2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(KEYINPUT58), .B(n1006), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1019) );
  XNOR2_X1 U1098 ( .A(KEYINPUT59), .B(KEYINPUT127), .ZN(n1009) );
  XNOR2_X1 U1099 ( .A(n1009), .B(G4), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(G1348), .B(n1010), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(G1981), .B(G6), .ZN(n1011) );
  NOR2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(G1341), .B(G19), .ZN(n1014) );
  XNOR2_X1 U1104 ( .A(G1956), .B(G20), .ZN(n1013) );
  NOR2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1106 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XOR2_X1 U1107 ( .A(KEYINPUT60), .B(n1017), .Z(n1018) );
  NAND2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1021) );
  XNOR2_X1 U1109 ( .A(G21), .B(G1966), .ZN(n1020) );
  NOR2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1111 ( .A(KEYINPUT61), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

