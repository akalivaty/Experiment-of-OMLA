//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n788, new_n789, new_n790, new_n791, new_n793,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1024, new_n1025, new_n1026,
    new_n1027;
  INV_X1    g000(.A(KEYINPUT39), .ZN(new_n202));
  NAND2_X1  g001(.A1(G225gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  AND2_X1   g003(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n206));
  OAI21_X1  g005(.A(G155gat), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT2), .ZN(new_n208));
  INV_X1    g007(.A(G141gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n209), .A2(KEYINPUT78), .A3(G148gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT78), .ZN(new_n211));
  INV_X1    g010(.A(G148gat), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n211), .B1(G141gat), .B2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(G141gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n210), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AND2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n208), .A2(new_n215), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT77), .B1(G155gat), .B2(G162gat), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NOR3_X1   g021(.A1(KEYINPUT77), .A2(G155gat), .A3(G162gat), .ZN(new_n223));
  NOR3_X1   g022(.A1(new_n222), .A2(new_n223), .A3(new_n216), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT2), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n209), .A2(G148gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(new_n214), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n220), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT80), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n220), .A2(KEYINPUT80), .A3(new_n228), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(KEYINPUT3), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT81), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n231), .A2(KEYINPUT81), .A3(KEYINPUT3), .A4(new_n232), .ZN(new_n236));
  INV_X1    g035(.A(G127gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n237), .A2(G134gat), .ZN(new_n238));
  INV_X1    g037(.A(G134gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n239), .A2(G127gat), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT67), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(G127gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n237), .A2(G134gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n241), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G113gat), .ZN(new_n247));
  INV_X1    g046(.A(G120gat), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT1), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(new_n247), .B2(new_n248), .ZN(new_n250));
  AND3_X1   g049(.A1(new_n249), .A2(new_n242), .A3(new_n243), .ZN(new_n251));
  XNOR2_X1  g050(.A(KEYINPUT68), .B(G113gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(G120gat), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n246), .A2(new_n250), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  XOR2_X1   g054(.A(KEYINPUT82), .B(KEYINPUT3), .Z(new_n256));
  NAND3_X1  g055(.A1(new_n220), .A2(new_n228), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n235), .A2(new_n236), .A3(new_n259), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n244), .B1(new_n242), .B2(new_n243), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n250), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n238), .A2(new_n240), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n253), .A2(new_n249), .A3(new_n264), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n220), .A2(new_n228), .A3(new_n263), .A4(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(KEYINPUT4), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n202), .B(new_n204), .C1(new_n260), .C2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G1gat), .B(G29gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT0), .ZN(new_n274));
  XNOR2_X1  g073(.A(G57gat), .B(G85gat), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n274), .B(new_n275), .Z(new_n276));
  AOI21_X1  g075(.A(new_n258), .B1(new_n233), .B2(new_n234), .ZN(new_n277));
  AOI22_X1  g076(.A1(new_n277), .A2(new_n236), .B1(new_n269), .B2(new_n270), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n278), .A2(new_n203), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n231), .A2(new_n232), .A3(new_n255), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(new_n266), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT39), .B1(new_n281), .B2(new_n204), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n272), .B(new_n276), .C1(new_n279), .C2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT40), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT88), .ZN(new_n286));
  OR2_X1    g085(.A1(new_n283), .A2(new_n284), .ZN(new_n287));
  XOR2_X1   g086(.A(G211gat), .B(G218gat), .Z(new_n288));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n289));
  XOR2_X1   g088(.A(G197gat), .B(G204gat), .Z(new_n290));
  AOI21_X1  g089(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  OR2_X1    g091(.A1(G197gat), .A2(G204gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(G197gat), .A2(G204gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n291), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n295), .A2(KEYINPUT74), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n288), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n288), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G226gat), .A2(G233gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n302), .B(KEYINPUT75), .ZN(new_n303));
  INV_X1    g102(.A(G169gat), .ZN(new_n304));
  INV_X1    g103(.A(G176gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(new_n305), .A3(KEYINPUT23), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT23), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(G169gat), .B2(G176gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n306), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT25), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n315));
  INV_X1    g114(.A(G183gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT65), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT65), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G183gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n314), .B(new_n315), .C1(new_n320), .C2(G190gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n312), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G190gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n316), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n315), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT64), .ZN(new_n326));
  NAND2_X1  g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT24), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n326), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n310), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n322), .B1(new_n332), .B2(KEYINPUT25), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT27), .ZN(new_n334));
  AOI21_X1  g133(.A(G190gat), .B1(new_n334), .B2(G183gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n316), .A2(KEYINPUT27), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(KEYINPUT28), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT27), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT66), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n317), .A2(new_n319), .A3(KEYINPUT66), .A4(KEYINPUT27), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(new_n342), .A3(new_n335), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT28), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n338), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n309), .ZN(new_n346));
  NOR2_X1   g145(.A1(G169gat), .A2(G176gat), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n346), .A2(new_n347), .A3(KEYINPUT26), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(KEYINPUT26), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n327), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n333), .B1(new_n345), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT29), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n303), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n342), .A2(new_n335), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT65), .B(G183gat), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT66), .B1(new_n357), .B2(KEYINPUT27), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n344), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n337), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n351), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n302), .B1(new_n361), .B2(new_n333), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n301), .B1(new_n355), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n288), .ZN(new_n364));
  AOI211_X1 g163(.A(new_n289), .B(new_n291), .C1(new_n293), .C2(new_n294), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT74), .B1(new_n295), .B2(new_n296), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n299), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n303), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT29), .B1(new_n361), .B2(new_n333), .ZN(new_n370));
  INV_X1    g169(.A(new_n302), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n368), .B(new_n369), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(G64gat), .B(G92gat), .Z(new_n373));
  XNOR2_X1  g172(.A(G8gat), .B(G36gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n363), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n375), .B(KEYINPUT76), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n378), .B1(new_n363), .B2(new_n372), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT30), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT30), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n204), .A2(KEYINPUT5), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n278), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT83), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n385), .B1(new_n266), .B2(KEYINPUT4), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n209), .A2(G148gat), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(new_n226), .B2(new_n211), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n218), .B1(new_n388), .B2(new_n210), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n389), .A2(new_n208), .B1(new_n227), .B2(new_n224), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n390), .A2(new_n254), .A3(KEYINPUT83), .A4(new_n268), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n386), .A2(new_n270), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n203), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT5), .B1(new_n260), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT84), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n395), .B1(new_n281), .B2(new_n204), .ZN(new_n396));
  AOI211_X1 g195(.A(KEYINPUT84), .B(new_n203), .C1(new_n280), .C2(new_n266), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n384), .B1(new_n394), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n276), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n380), .A2(new_n382), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT88), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n283), .A2(new_n402), .A3(new_n284), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n286), .A2(new_n287), .A3(new_n401), .A4(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT89), .B(KEYINPUT37), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n363), .A2(new_n372), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n368), .B1(new_n355), .B2(new_n362), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n301), .B(new_n369), .C1(new_n370), .C2(new_n371), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n407), .A2(new_n408), .A3(KEYINPUT37), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n378), .A2(KEYINPUT38), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n406), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n376), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n363), .A2(new_n372), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT37), .ZN(new_n414));
  INV_X1    g213(.A(new_n375), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n415), .A3(new_n406), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n412), .B1(KEYINPUT38), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n399), .A2(new_n400), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT6), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n276), .B(new_n384), .C1(new_n394), .C2(new_n398), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n399), .A2(KEYINPUT6), .A3(new_n400), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n417), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n257), .A2(new_n354), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(new_n301), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT85), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT29), .B1(new_n367), .B2(new_n299), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n231), .B(new_n232), .C1(new_n428), .C2(KEYINPUT3), .ZN(new_n429));
  INV_X1    g228(.A(G228gat), .ZN(new_n430));
  INV_X1    g229(.A(G233gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n424), .A2(new_n301), .A3(KEYINPUT85), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n427), .A2(new_n429), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(G22gat), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n354), .B1(new_n298), .B2(new_n300), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n390), .B1(new_n436), .B2(new_n256), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n368), .B1(new_n354), .B2(new_n257), .ZN(new_n438));
  OAI22_X1  g237(.A1(new_n437), .A2(new_n438), .B1(new_n430), .B2(new_n431), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n434), .A2(new_n435), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT86), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(G78gat), .B(G106gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT31), .B(G50gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n434), .A2(new_n439), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(G22gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n440), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n448), .A2(KEYINPUT86), .A3(new_n440), .A4(new_n445), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n404), .A2(new_n423), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n352), .B1(new_n359), .B2(new_n337), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n308), .A2(new_n309), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n324), .B(new_n315), .C1(new_n313), .C2(new_n326), .ZN(new_n456));
  INV_X1    g255(.A(new_n331), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n455), .B(new_n306), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  AOI22_X1  g257(.A1(new_n458), .A2(new_n311), .B1(new_n321), .B2(new_n312), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n254), .B1(new_n454), .B2(new_n459), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n255), .B(new_n333), .C1(new_n345), .C2(new_n352), .ZN(new_n461));
  NAND2_X1  g260(.A1(G227gat), .A2(G233gat), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(new_n461), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT33), .ZN(new_n465));
  XOR2_X1   g264(.A(G15gat), .B(G43gat), .Z(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(KEYINPUT70), .ZN(new_n467));
  XNOR2_X1  g266(.A(G71gat), .B(G99gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n467), .B(new_n468), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n464), .B(KEYINPUT32), .C1(new_n465), .C2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n469), .B1(new_n464), .B2(KEYINPUT32), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n464), .A2(KEYINPUT69), .A3(new_n465), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT69), .B1(new_n464), .B2(new_n465), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT72), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n463), .B1(new_n460), .B2(new_n461), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n479), .A2(KEYINPUT71), .A3(KEYINPUT34), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT34), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT71), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n481), .B1(new_n478), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n477), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n475), .A2(new_n476), .A3(new_n484), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(KEYINPUT36), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT73), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n484), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n480), .A2(KEYINPUT73), .A3(new_n483), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(new_n475), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT36), .ZN(new_n493));
  INV_X1    g292(.A(new_n474), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n494), .A2(new_n472), .A3(new_n471), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n495), .A2(new_n484), .A3(new_n489), .A4(new_n470), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n492), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n488), .A2(new_n497), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n450), .A2(KEYINPUT87), .A3(new_n451), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT87), .B1(new_n450), .B2(new_n451), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n380), .A2(new_n382), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n502), .B1(new_n421), .B2(new_n422), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n498), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT35), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n452), .A2(new_n486), .A3(new_n487), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n505), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(new_n502), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n420), .A2(new_n419), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT5), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n391), .A2(new_n270), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n204), .B1(new_n511), .B2(new_n386), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n235), .A2(new_n236), .A3(new_n259), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n510), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n220), .A2(KEYINPUT80), .A3(new_n228), .ZN(new_n515));
  AOI21_X1  g314(.A(KEYINPUT80), .B1(new_n220), .B2(new_n228), .ZN(new_n516));
  NOR3_X1   g315(.A1(new_n515), .A2(new_n516), .A3(new_n254), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n204), .B1(new_n517), .B2(new_n267), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT84), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n281), .A2(new_n395), .A3(new_n204), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n514), .A2(new_n521), .B1(new_n278), .B2(new_n383), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n522), .A2(new_n276), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n509), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n422), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n508), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n492), .A2(new_n496), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n527), .A2(new_n505), .A3(new_n452), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  OAI22_X1  g328(.A1(new_n453), .A2(new_n504), .B1(new_n507), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT96), .ZN(new_n531));
  INV_X1    g330(.A(G50gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(G43gat), .ZN(new_n533));
  INV_X1    g332(.A(G43gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(G50gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n533), .A2(new_n535), .A3(KEYINPUT15), .ZN(new_n536));
  NOR2_X1   g335(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n537));
  INV_X1    g336(.A(G36gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT90), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n537), .A2(KEYINPUT90), .A3(new_n538), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  AND2_X1   g343(.A1(KEYINPUT91), .A2(G29gat), .ZN(new_n545));
  NOR2_X1   g344(.A1(KEYINPUT91), .A2(G29gat), .ZN(new_n546));
  OAI21_X1  g345(.A(G36gat), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n536), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n539), .A2(new_n543), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n549), .A2(new_n547), .A3(new_n536), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT93), .ZN(new_n551));
  AND2_X1   g350(.A1(KEYINPUT92), .A2(G43gat), .ZN(new_n552));
  NOR2_X1   g351(.A1(KEYINPUT92), .A2(G43gat), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n551), .B(new_n532), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT15), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT92), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(new_n534), .ZN(new_n557));
  NAND2_X1  g356(.A1(KEYINPUT92), .A2(G43gat), .ZN(new_n558));
  AOI21_X1  g357(.A(G50gat), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n535), .A2(KEYINPUT93), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n554), .B(new_n555), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n550), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT94), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT94), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n550), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n548), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT95), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n435), .A2(G15gat), .ZN(new_n568));
  INV_X1    g367(.A(G15gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(G22gat), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n567), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n568), .A2(new_n570), .A3(new_n567), .ZN(new_n573));
  INV_X1    g372(.A(G1gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(KEYINPUT16), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n568), .A2(new_n570), .A3(new_n567), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n576), .B1(new_n577), .B2(new_n571), .ZN(new_n578));
  INV_X1    g377(.A(G8gat), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n575), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n579), .B1(new_n575), .B2(new_n578), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n531), .B1(new_n566), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n548), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n550), .A2(new_n561), .A3(new_n564), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n564), .B1(new_n550), .B2(new_n561), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n575), .A2(new_n578), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(G8gat), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n575), .A2(new_n578), .A3(new_n579), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n587), .A2(new_n591), .A3(KEYINPUT96), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n583), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G229gat), .A2(G233gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT17), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n587), .A2(new_n595), .ZN(new_n596));
  OAI211_X1 g395(.A(KEYINPUT17), .B(new_n584), .C1(new_n585), .C2(new_n586), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n596), .A2(new_n582), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n593), .A2(new_n594), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT18), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n593), .A2(KEYINPUT18), .A3(new_n594), .A4(new_n598), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n566), .A2(new_n582), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n593), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n594), .B(KEYINPUT13), .Z(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n601), .A2(new_n602), .A3(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G113gat), .B(G141gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(G197gat), .ZN(new_n609));
  XOR2_X1   g408(.A(KEYINPUT11), .B(G169gat), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT97), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n601), .A2(new_n606), .A3(new_n612), .A4(new_n602), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n607), .A2(KEYINPUT97), .A3(new_n613), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n530), .A2(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n622), .A2(KEYINPUT41), .ZN(new_n623));
  XNOR2_X1  g422(.A(G134gat), .B(G162gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G85gat), .A2(G92gat), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT7), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G99gat), .A2(G106gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT8), .ZN(new_n631));
  OR2_X1    g430(.A1(G85gat), .A2(G92gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(KEYINPUT101), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT101), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n631), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n629), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(G99gat), .B(G106gat), .Z(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(KEYINPUT103), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n627), .B(KEYINPUT7), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n631), .A2(new_n635), .A3(new_n632), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n635), .B1(new_n631), .B2(new_n632), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT103), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n644), .A2(new_n645), .A3(new_n638), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT102), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n637), .B2(new_n639), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n639), .B(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(KEYINPUT102), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n640), .B(new_n646), .C1(new_n648), .C2(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n651), .A2(new_n566), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(KEYINPUT41), .B2(new_n622), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n596), .A2(new_n597), .A3(new_n651), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(G190gat), .B(G218gat), .Z(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n655), .A2(new_n656), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n626), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n659), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n661), .A2(new_n625), .A3(new_n657), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AND2_X1   g463(.A1(G71gat), .A2(G78gat), .ZN(new_n665));
  NOR2_X1   g464(.A1(G71gat), .A2(G78gat), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g466(.A(G57gat), .B(G64gat), .Z(new_n668));
  INV_X1    g467(.A(KEYINPUT98), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n668), .B1(KEYINPUT9), .B2(new_n665), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n672), .A2(KEYINPUT21), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n591), .B1(KEYINPUT21), .B2(new_n672), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n675), .B(new_n676), .Z(new_n677));
  XNOR2_X1  g476(.A(G127gat), .B(G155gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT20), .ZN(new_n679));
  NAND2_X1  g478(.A1(G231gat), .A2(G233gat), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(KEYINPUT99), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n679), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(G183gat), .B(G211gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n677), .B(new_n684), .Z(new_n685));
  INV_X1    g484(.A(new_n672), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n651), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n644), .A2(new_n638), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n672), .A2(new_n649), .A3(new_n688), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(G230gat), .A2(G233gat), .ZN(new_n691));
  OR3_X1    g490(.A1(new_n690), .A2(KEYINPUT104), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT10), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n687), .A2(new_n693), .A3(new_n689), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n672), .A2(KEYINPUT10), .ZN(new_n695));
  OR2_X1    g494(.A1(new_n651), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n691), .ZN(new_n698));
  XNOR2_X1  g497(.A(G120gat), .B(G148gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(G176gat), .B(G204gat), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n699), .B(new_n700), .Z(new_n701));
  OAI21_X1  g500(.A(KEYINPUT104), .B1(new_n690), .B2(new_n691), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n692), .A2(new_n698), .A3(new_n701), .A4(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n701), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n690), .A2(new_n691), .ZN(new_n705));
  INV_X1    g504(.A(new_n691), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n706), .B1(new_n694), .B2(new_n696), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n704), .B1(new_n705), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n664), .A2(new_n685), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n621), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(new_n524), .B2(new_n525), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n421), .A2(KEYINPUT105), .A3(new_n422), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(new_n574), .ZN(G1324gat));
  INV_X1    g517(.A(KEYINPUT106), .ZN(new_n719));
  OAI21_X1  g518(.A(G8gat), .B1(new_n711), .B2(new_n508), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT16), .B(G8gat), .Z(new_n721));
  NAND4_X1  g520(.A1(new_n621), .A2(new_n502), .A3(new_n710), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(KEYINPUT42), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT42), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n719), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n725), .B1(new_n720), .B2(new_n722), .ZN(new_n728));
  INV_X1    g527(.A(new_n726), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n728), .A2(new_n729), .A3(KEYINPUT106), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n727), .A2(new_n730), .ZN(G1325gat));
  OAI21_X1  g530(.A(G15gat), .B1(new_n711), .B2(new_n498), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n527), .A2(new_n569), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n711), .B2(new_n733), .ZN(G1326gat));
  NOR2_X1   g533(.A1(new_n711), .A2(new_n501), .ZN(new_n735));
  XOR2_X1   g534(.A(KEYINPUT43), .B(G22gat), .Z(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1327gat));
  NAND2_X1  g536(.A1(new_n530), .A2(new_n620), .ZN(new_n738));
  INV_X1    g537(.A(new_n709), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n685), .A2(new_n739), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n738), .A2(new_n663), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n545), .A2(new_n546), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n741), .A2(new_n742), .A3(new_n715), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT45), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n530), .A2(KEYINPUT107), .A3(new_n664), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n530), .A2(KEYINPUT107), .A3(KEYINPUT44), .A4(new_n664), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n740), .A2(new_n619), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(new_n716), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n744), .B1(new_n742), .B2(new_n752), .ZN(G1328gat));
  NAND3_X1  g552(.A1(new_n741), .A2(new_n538), .A3(new_n502), .ZN(new_n754));
  XOR2_X1   g553(.A(new_n754), .B(KEYINPUT46), .Z(new_n755));
  OAI21_X1  g554(.A(G36gat), .B1(new_n751), .B2(new_n508), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(G1329gat));
  INV_X1    g556(.A(new_n498), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n747), .A2(new_n758), .A3(new_n748), .A4(new_n750), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n557), .A2(new_n558), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n762));
  INV_X1    g561(.A(new_n527), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n763), .A2(new_n760), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n762), .B1(new_n741), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(G1330gat));
  OAI21_X1  g567(.A(G50gat), .B1(new_n751), .B2(new_n452), .ZN(new_n769));
  INV_X1    g568(.A(new_n501), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n741), .A2(new_n532), .A3(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT48), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n749), .A2(new_n770), .A3(new_n750), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n771), .B1(new_n775), .B2(G50gat), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n774), .B1(KEYINPUT48), .B2(new_n776), .ZN(G1331gat));
  NOR2_X1   g576(.A1(new_n664), .A2(new_n685), .ZN(new_n778));
  AND4_X1   g577(.A1(new_n530), .A2(new_n619), .A3(new_n709), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n715), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g580(.A(new_n502), .B(KEYINPUT109), .Z(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n785));
  XOR2_X1   g584(.A(KEYINPUT49), .B(G64gat), .Z(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n784), .B2(new_n786), .ZN(G1333gat));
  NAND2_X1  g586(.A1(new_n779), .A2(new_n758), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n763), .A2(G71gat), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n788), .A2(G71gat), .B1(new_n779), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g589(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n790), .B(new_n791), .ZN(G1334gat));
  NAND2_X1  g591(.A1(new_n779), .A2(new_n770), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(G78gat), .ZN(G1335gat));
  INV_X1    g593(.A(new_n685), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n620), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n530), .A2(new_n664), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT51), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n530), .A2(KEYINPUT51), .A3(new_n664), .A4(new_n796), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n716), .A2(G85gat), .A3(new_n739), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n620), .A2(new_n795), .A3(new_n739), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n749), .A2(new_n715), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT111), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G85gat), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n805), .A2(new_n806), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n803), .B1(new_n808), .B2(new_n809), .ZN(G1336gat));
  NAND3_X1  g609(.A1(new_n749), .A2(new_n783), .A3(new_n804), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(new_n812), .A3(G92gat), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n782), .A2(G92gat), .A3(new_n739), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n801), .A2(new_n814), .B1(KEYINPUT112), .B2(KEYINPUT52), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n749), .A2(new_n502), .A3(new_n804), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n801), .A2(new_n814), .ZN(new_n818));
  AOI22_X1  g617(.A1(new_n817), .A2(G92gat), .B1(new_n818), .B2(KEYINPUT112), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n816), .B1(new_n819), .B2(new_n812), .ZN(G1337gat));
  NAND3_X1  g619(.A1(new_n749), .A2(new_n758), .A3(new_n804), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(G99gat), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n763), .A2(new_n739), .A3(G99gat), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n801), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(G1338gat));
  INV_X1    g624(.A(new_n452), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n749), .A2(new_n826), .A3(new_n804), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(G106gat), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n739), .A2(new_n452), .A3(G106gat), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n801), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n828), .A2(new_n829), .A3(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n747), .A2(new_n770), .A3(new_n748), .A4(new_n804), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(G106gat), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n831), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n833), .B1(new_n836), .B2(KEYINPUT53), .ZN(new_n837));
  AOI22_X1  g636(.A1(new_n834), .A2(G106gat), .B1(new_n801), .B2(new_n830), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n838), .A2(KEYINPUT113), .A3(new_n829), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n832), .B1(new_n837), .B2(new_n839), .ZN(G1339gat));
  NAND3_X1  g639(.A1(new_n778), .A2(new_n619), .A3(new_n739), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n604), .A2(new_n605), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n594), .B1(new_n593), .B2(new_n598), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n611), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n616), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n709), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n694), .A2(new_n706), .A3(new_n696), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n694), .A2(KEYINPUT114), .A3(new_n706), .A4(new_n696), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n850), .A2(new_n698), .A3(KEYINPUT54), .A4(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n701), .B1(new_n707), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT55), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n852), .A2(KEYINPUT55), .A3(new_n854), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n703), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n847), .B1(new_n859), .B2(new_n619), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n663), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n662), .A3(new_n660), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n842), .B1(new_n865), .B2(new_n685), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n770), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n716), .A2(new_n783), .A3(new_n763), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G113gat), .B1(new_n869), .B2(new_n619), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n863), .B1(new_n860), .B2(new_n663), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n841), .B1(new_n871), .B2(new_n795), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n506), .A3(new_n715), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n873), .A2(new_n874), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n782), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n619), .A2(new_n252), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n870), .B1(new_n877), .B2(new_n878), .ZN(G1340gat));
  NOR3_X1   g678(.A1(new_n869), .A2(new_n248), .A3(new_n739), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n877), .A2(new_n739), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n881), .B2(new_n248), .ZN(G1341gat));
  OAI21_X1  g681(.A(G127gat), .B1(new_n869), .B2(new_n685), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n795), .A2(new_n237), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n877), .B2(new_n884), .ZN(G1342gat));
  NOR3_X1   g684(.A1(new_n663), .A2(G134gat), .A3(new_n502), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n886), .B1(new_n875), .B2(new_n876), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n872), .A2(new_n868), .A3(new_n501), .A4(new_n664), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(G134gat), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT117), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n888), .A2(KEYINPUT117), .A3(G134gat), .ZN(new_n892));
  AOI22_X1  g691(.A1(new_n887), .A2(KEYINPUT56), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT56), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n894), .B(new_n886), .C1(new_n875), .C2(new_n876), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n895), .A2(KEYINPUT116), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n895), .A2(KEYINPUT116), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n893), .B1(new_n896), .B2(new_n897), .ZN(G1343gat));
  INV_X1    g697(.A(KEYINPUT57), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n857), .A2(KEYINPUT118), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n858), .A2(new_n703), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT55), .B1(new_n852), .B2(new_n854), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n900), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n847), .B1(new_n905), .B2(new_n619), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n863), .B1(new_n906), .B2(new_n663), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n841), .B1(new_n907), .B2(new_n795), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n899), .B1(new_n908), .B2(new_n770), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n872), .A2(new_n899), .A3(new_n826), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n715), .A2(new_n498), .A3(new_n782), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n209), .B1(new_n914), .B2(new_n620), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n758), .A2(new_n452), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n872), .A2(new_n715), .A3(new_n782), .A4(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n619), .A2(G141gat), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT120), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT119), .B1(new_n917), .B2(new_n919), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n922));
  AND3_X1   g721(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT58), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n922), .B1(new_n921), .B2(KEYINPUT58), .ZN(new_n924));
  OAI22_X1  g723(.A1(new_n915), .A2(new_n920), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n902), .A2(new_n903), .ZN(new_n926));
  AOI211_X1 g725(.A(KEYINPUT118), .B(KEYINPUT55), .C1(new_n852), .C2(new_n854), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n858), .A2(new_n703), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AOI22_X1  g728(.A1(new_n929), .A2(new_n620), .B1(new_n709), .B2(new_n846), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n864), .B1(new_n930), .B2(new_n664), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n842), .B1(new_n931), .B2(new_n685), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT57), .B1(new_n932), .B2(new_n501), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n901), .A2(new_n618), .A3(new_n617), .A4(new_n857), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n664), .B1(new_n934), .B2(new_n847), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n685), .B1(new_n935), .B2(new_n863), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n452), .B1(new_n936), .B2(new_n841), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n911), .B1(new_n937), .B2(new_n899), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n933), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(G141gat), .B1(new_n939), .B2(new_n619), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n921), .A2(KEYINPUT58), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT121), .ZN(new_n942));
  INV_X1    g741(.A(new_n920), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT58), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n940), .A2(new_n942), .A3(new_n943), .A4(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n925), .A2(new_n945), .ZN(G1344gat));
  AOI211_X1 g745(.A(KEYINPUT59), .B(new_n212), .C1(new_n914), .C2(new_n709), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT59), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n907), .A2(new_n795), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n841), .B(KEYINPUT122), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n899), .B(new_n770), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(KEYINPUT57), .B1(new_n866), .B2(new_n452), .ZN(new_n952));
  NAND4_X1  g751(.A1(new_n951), .A2(new_n709), .A3(new_n912), .A4(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n948), .B1(new_n953), .B2(G148gat), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n709), .A2(new_n212), .ZN(new_n955));
  OAI22_X1  g754(.A1(new_n947), .A2(new_n954), .B1(new_n917), .B2(new_n955), .ZN(G1345gat));
  INV_X1    g755(.A(G155gat), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n685), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(KEYINPUT123), .ZN(new_n959));
  AND3_X1   g758(.A1(new_n872), .A2(new_n715), .A3(new_n916), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n960), .A2(new_n795), .A3(new_n782), .ZN(new_n961));
  AOI22_X1  g760(.A1(new_n914), .A2(new_n959), .B1(new_n961), .B2(new_n957), .ZN(G1346gat));
  NOR2_X1   g761(.A1(new_n205), .A2(new_n206), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n960), .A2(new_n963), .A3(new_n508), .A4(new_n664), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n939), .A2(new_n663), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(new_n963), .ZN(G1347gat));
  NAND2_X1  g765(.A1(new_n716), .A2(new_n502), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n967), .A2(new_n763), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n867), .A2(new_n968), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n969), .A2(new_n304), .A3(new_n619), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT124), .ZN(new_n971));
  NOR3_X1   g770(.A1(new_n866), .A2(new_n971), .A3(new_n715), .ZN(new_n972));
  INV_X1    g771(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT124), .B1(new_n872), .B2(new_n716), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n783), .A2(new_n506), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n976), .A2(new_n620), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n970), .B1(new_n978), .B2(new_n304), .ZN(G1348gat));
  OAI21_X1  g778(.A(G176gat), .B1(new_n969), .B2(new_n739), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n976), .A2(new_n977), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n709), .A2(new_n305), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(G1349gat));
  NAND3_X1  g782(.A1(new_n867), .A2(new_n795), .A3(new_n968), .ZN(new_n984));
  AOI22_X1  g783(.A1(new_n984), .A2(new_n320), .B1(KEYINPUT125), .B2(KEYINPUT60), .ZN(new_n985));
  OR2_X1    g784(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n334), .A2(G183gat), .ZN(new_n987));
  AND3_X1   g786(.A1(new_n795), .A2(new_n987), .A3(new_n336), .ZN(new_n988));
  OAI211_X1 g787(.A(new_n977), .B(new_n988), .C1(new_n972), .C2(new_n974), .ZN(new_n989));
  AND3_X1   g788(.A1(new_n985), .A2(new_n986), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n986), .B1(new_n985), .B2(new_n989), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n990), .A2(new_n991), .ZN(G1350gat));
  NAND2_X1  g791(.A1(new_n664), .A2(new_n323), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n867), .A2(new_n664), .A3(new_n968), .ZN(new_n994));
  NOR2_X1   g793(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n323), .B1(KEYINPUT126), .B2(KEYINPUT61), .ZN(new_n996));
  AND3_X1   g795(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n995), .B1(new_n994), .B2(new_n996), .ZN(new_n998));
  OAI22_X1  g797(.A1(new_n981), .A2(new_n993), .B1(new_n997), .B2(new_n998), .ZN(G1351gat));
  NAND2_X1  g798(.A1(new_n916), .A2(new_n783), .ZN(new_n1000));
  AOI21_X1  g799(.A(new_n1000), .B1(new_n973), .B2(new_n975), .ZN(new_n1001));
  AOI21_X1  g800(.A(G197gat), .B1(new_n1001), .B2(new_n620), .ZN(new_n1002));
  AND2_X1   g801(.A1(new_n951), .A2(new_n952), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n967), .A2(new_n758), .ZN(new_n1004));
  AND2_X1   g803(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AND2_X1   g804(.A1(new_n620), .A2(G197gat), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n1002), .B1(new_n1005), .B2(new_n1006), .ZN(G1352gat));
  NAND4_X1  g806(.A1(new_n951), .A2(new_n709), .A3(new_n952), .A4(new_n1004), .ZN(new_n1008));
  INV_X1    g807(.A(new_n1000), .ZN(new_n1009));
  NOR2_X1   g808(.A1(new_n739), .A2(G204gat), .ZN(new_n1010));
  OAI211_X1 g809(.A(new_n1009), .B(new_n1010), .C1(new_n972), .C2(new_n974), .ZN(new_n1011));
  AOI22_X1  g810(.A1(G204gat), .A2(new_n1008), .B1(new_n1011), .B2(KEYINPUT62), .ZN(new_n1012));
  NOR2_X1   g811(.A1(new_n1011), .A2(KEYINPUT62), .ZN(new_n1013));
  INV_X1    g812(.A(KEYINPUT127), .ZN(new_n1014));
  NOR2_X1   g813(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NOR3_X1   g814(.A1(new_n1011), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n1016));
  OAI21_X1  g815(.A(new_n1012), .B1(new_n1015), .B2(new_n1016), .ZN(G1353gat));
  NAND4_X1  g816(.A1(new_n951), .A2(new_n795), .A3(new_n952), .A4(new_n1004), .ZN(new_n1018));
  AND3_X1   g817(.A1(new_n1018), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1019));
  AOI21_X1  g818(.A(KEYINPUT63), .B1(new_n1018), .B2(G211gat), .ZN(new_n1020));
  INV_X1    g819(.A(new_n1001), .ZN(new_n1021));
  OR2_X1    g820(.A1(new_n685), .A2(G211gat), .ZN(new_n1022));
  OAI22_X1  g821(.A1(new_n1019), .A2(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(G1354gat));
  NAND3_X1  g822(.A1(new_n1003), .A2(new_n664), .A3(new_n1004), .ZN(new_n1024));
  NAND2_X1  g823(.A1(new_n1024), .A2(G218gat), .ZN(new_n1025));
  INV_X1    g824(.A(G218gat), .ZN(new_n1026));
  NAND3_X1  g825(.A1(new_n1001), .A2(new_n1026), .A3(new_n664), .ZN(new_n1027));
  NAND2_X1  g826(.A1(new_n1025), .A2(new_n1027), .ZN(G1355gat));
endmodule


