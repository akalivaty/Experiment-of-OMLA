//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n812, new_n813, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920;
  XOR2_X1   g000(.A(G57gat), .B(G64gat), .Z(new_n202));
  AND2_X1   g001(.A1(G71gat), .A2(G78gat), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(KEYINPUT9), .B2(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(KEYINPUT9), .ZN(new_n205));
  NOR2_X1   g004(.A1(G71gat), .A2(G78gat), .ZN(new_n206));
  OAI22_X1  g005(.A1(new_n205), .A2(KEYINPUT93), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n204), .B(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT94), .B(KEYINPUT21), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G231gat), .A2(G233gat), .ZN(new_n211));
  XOR2_X1   g010(.A(new_n210), .B(new_n211), .Z(new_n212));
  XNOR2_X1  g011(.A(new_n212), .B(G127gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(G15gat), .B(G22gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT16), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n214), .B1(new_n215), .B2(G1gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(G1gat), .B2(new_n214), .ZN(new_n217));
  INV_X1    g016(.A(G8gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT21), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n219), .B1(new_n208), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n213), .B(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G183gat), .B(G211gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(KEYINPUT95), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n225));
  INV_X1    g024(.A(G155gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n224), .B(new_n227), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n222), .A2(new_n228), .ZN(new_n230));
  OR2_X1    g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G134gat), .B(G162gat), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n237));
  INV_X1    g036(.A(G29gat), .ZN(new_n238));
  INV_X1    g037(.A(G36gat), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(new_n239), .A3(KEYINPUT14), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT14), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(G29gat), .B2(G36gat), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n240), .B(new_n242), .C1(new_n238), .C2(new_n239), .ZN(new_n243));
  INV_X1    g042(.A(G43gat), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT15), .B1(new_n244), .B2(G50gat), .ZN(new_n245));
  INV_X1    g044(.A(G50gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n246), .A2(G43gat), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT15), .B1(new_n247), .B2(KEYINPUT86), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT86), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n251), .B1(new_n244), .B2(G50gat), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n250), .B1(new_n247), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  AND3_X1   g053(.A1(new_n243), .A2(KEYINPUT85), .A3(new_n248), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT85), .B1(new_n243), .B2(new_n248), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT87), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT87), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n254), .B(new_n259), .C1(new_n256), .C2(new_n255), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G85gat), .A2(G92gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT96), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(KEYINPUT96), .A2(G85gat), .A3(G92gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(KEYINPUT7), .A3(new_n265), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n262), .A2(KEYINPUT7), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n266), .A2(KEYINPUT97), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(G99gat), .A2(G106gat), .ZN(new_n269));
  INV_X1    g068(.A(G85gat), .ZN(new_n270));
  INV_X1    g069(.A(G92gat), .ZN(new_n271));
  AOI22_X1  g070(.A1(KEYINPUT8), .A2(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n272), .B1(new_n266), .B2(KEYINPUT97), .ZN(new_n273));
  XOR2_X1   g072(.A(G99gat), .B(G106gat), .Z(new_n274));
  OR3_X1    g073(.A1(new_n268), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n274), .B1(new_n268), .B2(new_n273), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n237), .B1(new_n261), .B2(new_n277), .ZN(new_n278));
  XOR2_X1   g077(.A(new_n278), .B(KEYINPUT98), .Z(new_n279));
  OAI21_X1  g078(.A(KEYINPUT88), .B1(new_n261), .B2(KEYINPUT17), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT88), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT17), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n258), .A2(new_n281), .A3(new_n282), .A4(new_n260), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  OR2_X1    g083(.A1(new_n257), .A2(new_n282), .ZN(new_n285));
  AND3_X1   g084(.A1(new_n284), .A2(new_n285), .A3(new_n277), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n279), .A2(new_n286), .ZN(new_n287));
  XOR2_X1   g086(.A(G190gat), .B(G218gat), .Z(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n287), .A2(new_n289), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n236), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n292), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(new_n235), .A3(new_n290), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G230gat), .ZN(new_n297));
  INV_X1    g096(.A(G233gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n277), .A2(new_n208), .ZN(new_n301));
  INV_X1    g100(.A(new_n208), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n302), .A2(new_n275), .A3(new_n276), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n304), .A2(KEYINPUT10), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT10), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n300), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n304), .A2(new_n299), .ZN(new_n309));
  XNOR2_X1  g108(.A(G120gat), .B(G148gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(G176gat), .B(G204gat), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n310), .B(new_n311), .Z(new_n312));
  NAND3_X1  g111(.A1(new_n308), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n312), .B1(new_n308), .B2(new_n309), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n232), .A2(new_n296), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT99), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT91), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT18), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n285), .A2(new_n219), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n323), .B1(new_n280), .B2(new_n283), .ZN(new_n324));
  NAND2_X1  g123(.A1(G229gat), .A2(G233gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n325), .B(KEYINPUT89), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n261), .A2(new_n219), .ZN(new_n327));
  NOR3_X1   g126(.A1(new_n324), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n322), .B1(new_n328), .B2(KEYINPUT90), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT90), .ZN(new_n330));
  NOR4_X1   g129(.A1(new_n324), .A2(new_n330), .A3(new_n326), .A4(new_n327), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n321), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n323), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n327), .B1(new_n284), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n326), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(new_n330), .ZN(new_n337));
  INV_X1    g136(.A(new_n331), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n337), .A2(new_n338), .A3(KEYINPUT91), .A4(new_n322), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n261), .B(new_n219), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n326), .B(KEYINPUT13), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n334), .A2(KEYINPUT18), .A3(new_n335), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n332), .A2(new_n339), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G113gat), .B(G141gat), .ZN(new_n345));
  INV_X1    g144(.A(G197gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT11), .B(G169gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n349), .B(KEYINPUT12), .Z(new_n350));
  NAND3_X1  g149(.A1(new_n337), .A2(new_n338), .A3(new_n322), .ZN(new_n351));
  INV_X1    g150(.A(new_n350), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n343), .A2(new_n352), .A3(new_n342), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT92), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n351), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT90), .B1(new_n334), .B2(new_n335), .ZN(new_n357));
  NOR3_X1   g156(.A1(new_n357), .A2(new_n331), .A3(KEYINPUT18), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT92), .B1(new_n358), .B2(new_n353), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n344), .A2(new_n350), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  XOR2_X1   g159(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n361));
  XOR2_X1   g160(.A(G127gat), .B(G134gat), .Z(new_n362));
  XNOR2_X1  g161(.A(G113gat), .B(G120gat), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n362), .B1(KEYINPUT1), .B2(new_n363), .ZN(new_n364));
  XOR2_X1   g163(.A(G113gat), .B(G120gat), .Z(new_n365));
  INV_X1    g164(.A(KEYINPUT1), .ZN(new_n366));
  XNOR2_X1  g165(.A(G127gat), .B(G134gat), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT76), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n364), .A2(new_n368), .A3(KEYINPUT76), .ZN(new_n372));
  XOR2_X1   g171(.A(G141gat), .B(G148gat), .Z(new_n373));
  INV_X1    g172(.A(G162gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n226), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G155gat), .A2(G162gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(KEYINPUT2), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n373), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G141gat), .B(G148gat), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n376), .B(new_n375), .C1(new_n380), .C2(KEYINPUT2), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n371), .A2(new_n372), .A3(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n368), .A2(new_n364), .A3(new_n379), .A4(new_n381), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G225gat), .A2(G233gat), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n361), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n382), .A2(KEYINPUT3), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT3), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n379), .A2(new_n381), .A3(new_n390), .ZN(new_n391));
  NAND4_X1  g190(.A1(new_n371), .A2(new_n389), .A3(new_n372), .A4(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n369), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n393), .A2(KEYINPUT4), .A3(new_n381), .A4(new_n379), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n384), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n392), .A2(new_n394), .A3(new_n386), .A4(new_n396), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n392), .A2(new_n386), .A3(new_n361), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n384), .A2(KEYINPUT4), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT79), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT79), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n401), .A3(KEYINPUT4), .ZN(new_n402));
  INV_X1    g201(.A(new_n395), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n400), .B(new_n402), .C1(new_n384), .C2(new_n403), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n388), .A2(new_n397), .B1(new_n398), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT6), .ZN(new_n406));
  XOR2_X1   g205(.A(G1gat), .B(G29gat), .Z(new_n407));
  XNOR2_X1  g206(.A(new_n407), .B(KEYINPUT0), .ZN(new_n408));
  XNOR2_X1  g207(.A(G57gat), .B(G85gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(new_n408), .B(new_n409), .ZN(new_n410));
  NOR3_X1   g209(.A1(new_n405), .A2(new_n406), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n388), .A2(new_n397), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n398), .A2(new_n404), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n410), .B(KEYINPUT81), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n412), .A2(new_n410), .A3(new_n413), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n406), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT83), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n411), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n417), .A2(KEYINPUT83), .A3(new_n406), .A4(new_n418), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT35), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT27), .B(G183gat), .ZN(new_n424));
  INV_X1    g223(.A(G190gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT28), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT68), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n426), .B(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(G169gat), .A2(G176gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  OR2_X1    g230(.A1(new_n431), .A2(KEYINPUT26), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(KEYINPUT26), .ZN(new_n433));
  NAND2_X1  g232(.A1(G169gat), .A2(G176gat), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(G183gat), .A2(G190gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OR2_X1    g236(.A1(new_n429), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT65), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n430), .B1(KEYINPUT23), .B2(new_n434), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT23), .ZN(new_n441));
  NOR3_X1   g240(.A1(new_n441), .A2(G169gat), .A3(G176gat), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n439), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n430), .A2(KEYINPUT23), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n441), .B1(G169gat), .B2(G176gat), .ZN(new_n445));
  OAI211_X1 g244(.A(KEYINPUT65), .B(new_n444), .C1(new_n445), .C2(new_n430), .ZN(new_n446));
  AND2_X1   g245(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT64), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n447), .A2(new_n448), .A3(G190gat), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n436), .ZN(new_n451));
  NAND3_X1  g250(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT64), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n449), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n443), .A2(new_n446), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT25), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT66), .ZN(new_n458));
  OAI211_X1 g257(.A(KEYINPUT25), .B(new_n444), .C1(new_n445), .C2(new_n430), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n436), .A2(new_n450), .B1(new_n447), .B2(G190gat), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n434), .A2(KEYINPUT23), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n442), .B1(new_n431), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n451), .A2(new_n452), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n463), .A2(KEYINPUT66), .A3(KEYINPUT25), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n457), .A2(new_n466), .A3(KEYINPUT67), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT67), .B1(new_n457), .B2(new_n466), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n438), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n369), .ZN(new_n470));
  NAND2_X1  g269(.A1(G227gat), .A2(G233gat), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n438), .B(new_n393), .C1(new_n467), .C2(new_n468), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT34), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT70), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT67), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n461), .A2(new_n465), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n444), .B1(new_n445), .B2(new_n430), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n450), .A2(new_n436), .B1(new_n452), .B2(KEYINPUT64), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n478), .A2(new_n439), .B1(new_n479), .B2(new_n449), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT25), .B1(new_n480), .B2(new_n446), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n476), .B1(new_n477), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n457), .A2(new_n466), .A3(KEYINPUT67), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n393), .B1(new_n484), .B2(new_n438), .ZN(new_n485));
  INV_X1    g284(.A(new_n472), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT34), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n487), .A2(KEYINPUT71), .A3(new_n488), .A4(new_n471), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n470), .A2(new_n488), .A3(new_n471), .A4(new_n472), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT71), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT70), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n473), .A2(new_n493), .A3(KEYINPUT34), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n475), .A2(new_n489), .A3(new_n492), .A4(new_n494), .ZN(new_n495));
  XOR2_X1   g294(.A(G71gat), .B(G99gat), .Z(new_n496));
  XNOR2_X1  g295(.A(G15gat), .B(G43gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n471), .B1(new_n470), .B2(new_n472), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT33), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n500), .A2(KEYINPUT32), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n498), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n500), .B1(new_n498), .B2(KEYINPUT69), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n503), .B1(KEYINPUT69), .B2(new_n498), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT32), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n502), .B1(new_n499), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n495), .A2(new_n506), .ZN(new_n507));
  AND3_X1   g306(.A1(new_n473), .A2(new_n493), .A3(KEYINPUT34), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n493), .B1(new_n473), .B2(KEYINPUT34), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n470), .A2(new_n472), .ZN(new_n511));
  INV_X1    g310(.A(new_n471), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n505), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n512), .B1(new_n485), .B2(new_n486), .ZN(new_n514));
  INV_X1    g313(.A(new_n501), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n513), .B1(new_n516), .B2(new_n498), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n490), .B(KEYINPUT71), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n510), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(G197gat), .B(G204gat), .ZN(new_n520));
  INV_X1    g319(.A(G211gat), .ZN(new_n521));
  INV_X1    g320(.A(G218gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n520), .B1(KEYINPUT22), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G211gat), .B(G218gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n390), .B1(new_n526), .B2(KEYINPUT29), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n382), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT29), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n391), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT80), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n391), .A2(KEYINPUT80), .A3(new_n529), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(new_n526), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n535), .A2(G228gat), .A3(G233gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(G228gat), .A2(G233gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n530), .A2(new_n526), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n528), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(KEYINPUT31), .B(G50gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n541), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n536), .A2(new_n539), .A3(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G78gat), .B(G106gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(G22gat), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n542), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n546), .B1(new_n542), .B2(new_n544), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g348(.A1(new_n423), .A2(new_n507), .A3(new_n519), .A4(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n457), .A2(new_n466), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n438), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT74), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G226gat), .A2(G233gat), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n438), .A2(new_n551), .A3(KEYINPUT74), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n556), .B1(new_n469), .B2(new_n529), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT73), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n429), .A2(new_n437), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n562), .B1(new_n482), .B2(new_n483), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n555), .B1(new_n563), .B2(KEYINPUT29), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n564), .A2(KEYINPUT73), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n526), .B1(new_n561), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(G8gat), .B(G36gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT75), .ZN(new_n568));
  XNOR2_X1  g367(.A(G64gat), .B(G92gat), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n568), .B(new_n569), .Z(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n554), .A2(new_n529), .A3(new_n555), .A4(new_n557), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n563), .A2(new_n556), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n526), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n566), .A2(new_n571), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT30), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n526), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n554), .A2(new_n557), .ZN(new_n580));
  AOI22_X1  g379(.A1(KEYINPUT73), .A2(new_n564), .B1(new_n580), .B2(new_n556), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n559), .A2(new_n560), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n570), .B1(new_n583), .B2(new_n574), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n566), .A2(KEYINPUT30), .A3(new_n571), .A4(new_n575), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n578), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n550), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n411), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n418), .A2(new_n406), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n405), .A2(new_n410), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n578), .A2(new_n584), .A3(new_n585), .A4(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n507), .A2(new_n519), .A3(new_n549), .ZN(new_n593));
  OAI21_X1  g392(.A(KEYINPUT35), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(KEYINPUT84), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT84), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n596), .B(KEYINPUT35), .C1(new_n592), .C2(new_n593), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n587), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n507), .A2(new_n519), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT72), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT36), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n600), .A2(KEYINPUT72), .A3(KEYINPUT36), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n386), .B1(new_n404), .B2(new_n392), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(KEYINPUT39), .B1(new_n385), .B2(new_n387), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n608), .B(new_n415), .C1(new_n606), .C2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT82), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT40), .ZN(new_n612));
  AND3_X1   g411(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n612), .B1(new_n610), .B2(new_n611), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n405), .A2(new_n415), .ZN(new_n615));
  NOR3_X1   g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n586), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n564), .A2(KEYINPUT73), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n618), .A2(new_n582), .A3(new_n558), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n574), .B1(new_n619), .B2(new_n526), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT37), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n571), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(new_n579), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n572), .A2(new_n573), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n621), .B1(new_n624), .B2(new_n526), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT38), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  AND3_X1   g426(.A1(new_n421), .A2(new_n576), .A3(new_n422), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT38), .ZN(new_n630));
  OAI21_X1  g429(.A(KEYINPUT37), .B1(new_n583), .B2(new_n574), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n630), .B1(new_n622), .B2(new_n631), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n617), .B(new_n549), .C1(new_n629), .C2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n549), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n592), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n605), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n360), .B1(new_n599), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n320), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n591), .B(KEYINPUT100), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n641), .B(G1gat), .Z(G1324gat));
  INV_X1    g441(.A(new_n586), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n638), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(KEYINPUT16), .B(G8gat), .Z(new_n645));
  AND2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n646), .A2(KEYINPUT42), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(KEYINPUT42), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n647), .B(new_n648), .C1(new_n218), .C2(new_n644), .ZN(G1325gat));
  XNOR2_X1  g448(.A(new_n605), .B(KEYINPUT101), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(G15gat), .B1(new_n638), .B2(new_n651), .ZN(new_n652));
  OR2_X1    g451(.A1(new_n600), .A2(G15gat), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n652), .B1(new_n638), .B2(new_n653), .ZN(G1326gat));
  NOR2_X1   g453(.A1(new_n638), .A2(new_n549), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT102), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT43), .B(G22gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(G1327gat));
  INV_X1    g457(.A(new_n316), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n232), .A2(new_n296), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n637), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n662), .A2(new_n238), .A3(new_n639), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT45), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n231), .B(KEYINPUT103), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n360), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(new_n667), .A3(new_n316), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n595), .A2(new_n597), .ZN(new_n671));
  INV_X1    g470(.A(new_n587), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AOI211_X1 g472(.A(KEYINPUT104), .B(new_n587), .C1(new_n595), .C2(new_n597), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n636), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n296), .A2(KEYINPUT44), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n296), .ZN(new_n678));
  AND4_X1   g477(.A1(new_n633), .A2(new_n635), .A3(new_n604), .A4(new_n603), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n679), .B2(new_n598), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n680), .A2(KEYINPUT44), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n669), .B1(new_n677), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(G29gat), .B1(new_n682), .B2(new_n640), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n664), .A2(new_n683), .ZN(G1328gat));
  NOR3_X1   g483(.A1(new_n661), .A2(G36gat), .A3(new_n643), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT46), .ZN(new_n686));
  OAI21_X1  g485(.A(G36gat), .B1(new_n682), .B2(new_n643), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(G1329gat));
  NOR2_X1   g487(.A1(new_n600), .A2(G43gat), .ZN(new_n689));
  AND3_X1   g488(.A1(new_n637), .A2(new_n660), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT106), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT108), .B1(new_n682), .B2(new_n605), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(G43gat), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n682), .A2(KEYINPUT108), .A3(new_n605), .ZN(new_n694));
  OAI211_X1 g493(.A(KEYINPUT47), .B(new_n691), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n675), .A2(new_n676), .B1(KEYINPUT44), .B2(new_n680), .ZN(new_n697));
  NOR3_X1   g496(.A1(new_n697), .A2(new_n651), .A3(new_n668), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n696), .B1(new_n698), .B2(new_n244), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n650), .B(new_n669), .C1(new_n677), .C2(new_n681), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n700), .A2(KEYINPUT105), .A3(G43gat), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n699), .A2(new_n701), .A3(new_n691), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT47), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n703), .B1(new_n702), .B2(new_n704), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n695), .B1(new_n705), .B2(new_n706), .ZN(G1330gat));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n682), .A2(new_n549), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n708), .B1(new_n709), .B2(new_n246), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT48), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n662), .A2(new_n246), .A3(new_n634), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(new_n709), .B2(new_n246), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n711), .B(new_n713), .ZN(G1331gat));
  INV_X1    g513(.A(new_n675), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n232), .A2(new_n360), .A3(new_n296), .A4(new_n659), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n639), .ZN(new_n718));
  XNOR2_X1  g517(.A(KEYINPUT110), .B(G57gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1332gat));
  NAND2_X1  g519(.A1(new_n717), .A2(KEYINPUT111), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(new_n715), .B2(new_n716), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n643), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n721), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n725), .A2(KEYINPUT112), .ZN(new_n726));
  NOR2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(KEYINPUT112), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n727), .B1(new_n726), .B2(new_n728), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(G1333gat));
  AND2_X1   g530(.A1(new_n721), .A2(new_n723), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n732), .A2(G71gat), .A3(new_n650), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n715), .A2(new_n600), .A3(new_n716), .ZN(new_n734));
  OR2_X1    g533(.A1(new_n734), .A2(G71gat), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n733), .A2(KEYINPUT50), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(KEYINPUT50), .B1(new_n733), .B2(new_n735), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(G1334gat));
  NAND2_X1  g537(.A1(new_n732), .A2(new_n634), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g539(.A1(new_n667), .A2(new_n232), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n659), .B(new_n741), .C1(new_n677), .C2(new_n681), .ZN(new_n742));
  OAI21_X1  g541(.A(G85gat), .B1(new_n742), .B2(new_n640), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n741), .A2(new_n678), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n715), .B2(new_n745), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n675), .A2(KEYINPUT51), .A3(new_n678), .A4(new_n741), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n639), .A2(new_n270), .A3(new_n659), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n743), .B1(new_n749), .B2(new_n750), .ZN(G1336gat));
  NOR3_X1   g550(.A1(new_n643), .A2(G92gat), .A3(new_n316), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n748), .A2(new_n752), .B1(new_n753), .B2(KEYINPUT52), .ZN(new_n754));
  OAI21_X1  g553(.A(G92gat), .B1(new_n742), .B2(new_n643), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n753), .A2(KEYINPUT52), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n756), .B(new_n757), .Z(G1337gat));
  OAI21_X1  g557(.A(G99gat), .B1(new_n742), .B2(new_n651), .ZN(new_n759));
  OR3_X1    g558(.A1(new_n600), .A2(G99gat), .A3(new_n316), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n759), .B1(new_n749), .B2(new_n760), .ZN(G1338gat));
  OAI21_X1  g560(.A(G106gat), .B1(new_n742), .B2(new_n549), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n549), .A2(new_n316), .A3(G106gat), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n356), .A2(new_n359), .ZN(new_n768));
  OAI22_X1  g567(.A1(new_n334), .A2(new_n335), .B1(new_n340), .B2(new_n341), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n349), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n768), .A2(new_n659), .A3(new_n770), .ZN(new_n771));
  OR3_X1    g570(.A1(new_n305), .A2(new_n307), .A3(new_n300), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n772), .A2(KEYINPUT54), .A3(new_n308), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT54), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n774), .B(new_n300), .C1(new_n305), .C2(new_n307), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT114), .ZN(new_n776));
  INV_X1    g575(.A(new_n312), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n776), .B1(new_n775), .B2(new_n777), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n773), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g581(.A(KEYINPUT55), .B(new_n773), .C1(new_n778), .C2(new_n779), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(new_n313), .A3(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n771), .B1(new_n360), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n296), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n296), .A2(new_n784), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n768), .A2(KEYINPUT115), .A3(new_n770), .ZN(new_n788));
  AOI21_X1  g587(.A(KEYINPUT115), .B1(new_n768), .B2(new_n770), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n665), .B1(new_n786), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n317), .A2(new_n667), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n767), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n792), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n768), .A2(new_n770), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n768), .A2(KEYINPUT115), .A3(new_n770), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AOI22_X1  g598(.A1(new_n799), .A2(new_n787), .B1(new_n785), .B2(new_n296), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n794), .B(KEYINPUT116), .C1(new_n800), .C2(new_n665), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n793), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n640), .A2(new_n586), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(new_n593), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n667), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n659), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(G120gat), .ZN(G1341gat));
  OAI21_X1  g610(.A(G127gat), .B1(new_n806), .B2(new_n666), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n231), .A2(G127gat), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n812), .B1(new_n806), .B2(new_n813), .ZN(new_n814));
  XOR2_X1   g613(.A(new_n814), .B(KEYINPUT117), .Z(G1342gat));
  OR3_X1    g614(.A1(new_n806), .A2(G134gat), .A3(new_n296), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n816), .A2(KEYINPUT56), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(KEYINPUT56), .ZN(new_n818));
  OAI21_X1  g617(.A(G134gat), .B1(new_n806), .B2(new_n296), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(G1343gat));
  INV_X1    g619(.A(KEYINPUT58), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n605), .A2(new_n803), .ZN(new_n822));
  INV_X1    g621(.A(G141gat), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n360), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n784), .A2(KEYINPUT119), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n784), .A2(KEYINPUT119), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n667), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n678), .B1(new_n829), .B2(new_n771), .ZN(new_n830));
  INV_X1    g629(.A(new_n790), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n231), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI211_X1 g631(.A(new_n826), .B(new_n549), .C1(new_n832), .C2(new_n794), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n793), .A2(new_n801), .A3(new_n634), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n826), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n833), .B1(new_n835), .B2(KEYINPUT118), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n834), .A2(new_n837), .A3(new_n826), .ZN(new_n838));
  AOI211_X1 g637(.A(new_n822), .B(new_n825), .C1(new_n836), .C2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n802), .A2(new_n634), .A3(new_n651), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n804), .ZN(new_n841));
  AOI21_X1  g640(.A(G141gat), .B1(new_n841), .B2(new_n667), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n821), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n822), .B1(new_n836), .B2(new_n838), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n824), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n841), .A2(new_n667), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n823), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n847), .A3(KEYINPUT58), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n843), .A2(new_n848), .ZN(G1344gat));
  INV_X1    g648(.A(G148gat), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n841), .A2(new_n850), .A3(new_n659), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n851), .A2(KEYINPUT120), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n851), .A2(KEYINPUT120), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n850), .A2(KEYINPUT59), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n854), .B1(new_n844), .B2(new_n659), .ZN(new_n855));
  XNOR2_X1  g654(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n832), .B1(new_n667), .B2(new_n319), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n549), .A2(KEYINPUT57), .ZN(new_n858));
  AOI22_X1  g657(.A1(KEYINPUT57), .A2(new_n834), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  XOR2_X1   g658(.A(new_n822), .B(KEYINPUT122), .Z(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n659), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n856), .B1(new_n861), .B2(G148gat), .ZN(new_n862));
  OAI22_X1  g661(.A1(new_n852), .A2(new_n853), .B1(new_n855), .B2(new_n862), .ZN(G1345gat));
  NAND3_X1  g662(.A1(new_n841), .A2(new_n226), .A3(new_n232), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n844), .A2(new_n665), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n864), .B1(new_n865), .B2(new_n226), .ZN(G1346gat));
  NAND3_X1  g665(.A1(new_n841), .A2(new_n374), .A3(new_n678), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n844), .A2(new_n678), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n867), .B1(new_n868), .B2(new_n374), .ZN(G1347gat));
  INV_X1    g668(.A(G169gat), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n643), .A2(new_n593), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n802), .A2(new_n640), .A3(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n870), .B1(new_n873), .B2(new_n667), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT124), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n874), .A2(new_n875), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n871), .B(KEYINPUT123), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n802), .A2(new_n640), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n667), .A2(new_n870), .ZN(new_n881));
  OAI22_X1  g680(.A1(new_n877), .A2(new_n878), .B1(new_n880), .B2(new_n881), .ZN(G1348gat));
  OAI21_X1  g681(.A(G176gat), .B1(new_n872), .B2(new_n316), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n316), .A2(G176gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n880), .B2(new_n884), .ZN(G1349gat));
  NAND2_X1  g684(.A1(new_n232), .A2(new_n424), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT125), .ZN(new_n888));
  OAI21_X1  g687(.A(G183gat), .B1(new_n872), .B2(new_n666), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g690(.A(G190gat), .B1(new_n872), .B2(new_n296), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT61), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n678), .A2(new_n425), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n880), .B2(new_n894), .ZN(G1351gat));
  NOR3_X1   g694(.A1(new_n650), .A2(new_n643), .A3(new_n639), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n859), .A2(new_n896), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n897), .A2(new_n346), .A3(new_n360), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n643), .A2(new_n639), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n802), .A2(new_n634), .A3(new_n651), .A4(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(G197gat), .B1(new_n901), .B2(new_n667), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n898), .A2(new_n902), .ZN(G1352gat));
  INV_X1    g702(.A(G204gat), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n659), .A2(new_n904), .ZN(new_n905));
  OR3_X1    g704(.A1(new_n900), .A2(KEYINPUT62), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT62), .B1(new_n900), .B2(new_n905), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n859), .A2(new_n659), .A3(new_n896), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n906), .B(new_n907), .C1(new_n904), .C2(new_n908), .ZN(G1353gat));
  NAND3_X1  g708(.A1(new_n901), .A2(new_n521), .A3(new_n232), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n859), .A2(new_n232), .A3(new_n896), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n911), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT63), .B1(new_n911), .B2(G211gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(G1354gat));
  NAND2_X1  g713(.A1(new_n678), .A2(G218gat), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n897), .A2(KEYINPUT127), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n897), .A2(KEYINPUT127), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n522), .B1(new_n900), .B2(new_n296), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT126), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n918), .A2(new_n920), .ZN(G1355gat));
endmodule


