

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590;

  XNOR2_X1 U324 ( .A(n369), .B(n381), .ZN(n370) );
  XNOR2_X1 U325 ( .A(KEYINPUT123), .B(KEYINPUT55), .ZN(n459) );
  XOR2_X1 U326 ( .A(n312), .B(n323), .Z(n529) );
  XNOR2_X1 U327 ( .A(n581), .B(n418), .ZN(n508) );
  INV_X1 U328 ( .A(KEYINPUT54), .ZN(n441) );
  XNOR2_X1 U329 ( .A(n417), .B(KEYINPUT64), .ZN(n418) );
  XNOR2_X1 U330 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U331 ( .A(n371), .B(n370), .ZN(n378) );
  XNOR2_X1 U332 ( .A(n460), .B(n459), .ZN(n461) );
  XOR2_X1 U333 ( .A(n334), .B(n333), .Z(n524) );
  XNOR2_X1 U334 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U335 ( .A(n466), .B(n465), .ZN(G1351GAT) );
  XOR2_X1 U336 ( .A(KEYINPUT93), .B(KEYINPUT90), .Z(n293) );
  XNOR2_X1 U337 ( .A(KEYINPUT91), .B(KEYINPUT20), .ZN(n292) );
  XNOR2_X1 U338 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U339 ( .A(G176GAT), .B(KEYINPUT94), .Z(n295) );
  XNOR2_X1 U340 ( .A(G113GAT), .B(G15GAT), .ZN(n294) );
  XNOR2_X1 U341 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U342 ( .A(n297), .B(n296), .Z(n308) );
  XOR2_X1 U343 ( .A(KEYINPUT17), .B(KEYINPUT92), .Z(n299) );
  XNOR2_X1 U344 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U346 ( .A(G169GAT), .B(n300), .Z(n429) );
  XOR2_X1 U347 ( .A(G120GAT), .B(G71GAT), .Z(n359) );
  XOR2_X1 U348 ( .A(G183GAT), .B(G99GAT), .Z(n302) );
  XNOR2_X1 U349 ( .A(G43GAT), .B(G190GAT), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U351 ( .A(n359), .B(n303), .Z(n305) );
  NAND2_X1 U352 ( .A1(G227GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n429), .B(n306), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n308), .B(n307), .ZN(n312) );
  XOR2_X1 U356 ( .A(KEYINPUT89), .B(G134GAT), .Z(n310) );
  XNOR2_X1 U357 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n309) );
  XNOR2_X1 U358 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U359 ( .A(KEYINPUT88), .B(n311), .ZN(n323) );
  INV_X1 U360 ( .A(n529), .ZN(n538) );
  XOR2_X1 U361 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n314) );
  XNOR2_X1 U362 ( .A(G141GAT), .B(KEYINPUT96), .ZN(n313) );
  XNOR2_X1 U363 ( .A(n314), .B(n313), .ZN(n450) );
  XOR2_X1 U364 ( .A(n450), .B(G57GAT), .Z(n316) );
  NAND2_X1 U365 ( .A1(G225GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n334) );
  XOR2_X1 U367 ( .A(KEYINPUT1), .B(KEYINPUT98), .Z(n318) );
  XNOR2_X1 U368 ( .A(KEYINPUT100), .B(KEYINPUT99), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U370 ( .A(KEYINPUT97), .B(KEYINPUT4), .Z(n320) );
  XNOR2_X1 U371 ( .A(KEYINPUT6), .B(KEYINPUT5), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U373 ( .A(n322), .B(n321), .Z(n332) );
  INV_X1 U374 ( .A(n323), .ZN(n330) );
  XOR2_X1 U375 ( .A(G85GAT), .B(G155GAT), .Z(n325) );
  XNOR2_X1 U376 ( .A(G120GAT), .B(G148GAT), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U378 ( .A(n326), .B(G162GAT), .Z(n328) );
  XOR2_X1 U379 ( .A(G113GAT), .B(G1GAT), .Z(n347) );
  XNOR2_X1 U380 ( .A(G29GAT), .B(n347), .ZN(n327) );
  XNOR2_X1 U381 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U382 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U383 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U384 ( .A(KEYINPUT71), .B(KEYINPUT29), .Z(n336) );
  XNOR2_X1 U385 ( .A(KEYINPUT30), .B(KEYINPUT69), .ZN(n335) );
  XNOR2_X1 U386 ( .A(n336), .B(n335), .ZN(n355) );
  XOR2_X1 U387 ( .A(G141GAT), .B(G197GAT), .Z(n338) );
  XNOR2_X1 U388 ( .A(G36GAT), .B(G50GAT), .ZN(n337) );
  XNOR2_X1 U389 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U390 ( .A(G8GAT), .B(G15GAT), .Z(n340) );
  XNOR2_X1 U391 ( .A(G169GAT), .B(G22GAT), .ZN(n339) );
  XNOR2_X1 U392 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U393 ( .A(n342), .B(n341), .Z(n353) );
  XOR2_X1 U394 ( .A(KEYINPUT70), .B(KEYINPUT72), .Z(n344) );
  XNOR2_X1 U395 ( .A(KEYINPUT68), .B(KEYINPUT73), .ZN(n343) );
  XNOR2_X1 U396 ( .A(n344), .B(n343), .ZN(n351) );
  XOR2_X1 U397 ( .A(G29GAT), .B(G43GAT), .Z(n346) );
  XNOR2_X1 U398 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n345) );
  XNOR2_X1 U399 ( .A(n346), .B(n345), .ZN(n406) );
  XOR2_X1 U400 ( .A(n406), .B(n347), .Z(n349) );
  NAND2_X1 U401 ( .A1(G229GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U402 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U403 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U404 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U405 ( .A(n355), .B(n354), .Z(n577) );
  INV_X1 U406 ( .A(n577), .ZN(n564) );
  XOR2_X1 U407 ( .A(KEYINPUT80), .B(KEYINPUT31), .Z(n357) );
  XNOR2_X1 U408 ( .A(KEYINPUT33), .B(KEYINPUT75), .ZN(n356) );
  XNOR2_X1 U409 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U410 ( .A(n359), .B(n358), .ZN(n361) );
  AND2_X1 U411 ( .A1(G230GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U412 ( .A(n361), .B(n360), .ZN(n364) );
  INV_X1 U413 ( .A(n364), .ZN(n362) );
  NAND2_X1 U414 ( .A1(n362), .A2(KEYINPUT76), .ZN(n366) );
  INV_X1 U415 ( .A(KEYINPUT76), .ZN(n363) );
  NAND2_X1 U416 ( .A1(n364), .A2(n363), .ZN(n365) );
  NAND2_X1 U417 ( .A1(n366), .A2(n365), .ZN(n371) );
  XNOR2_X1 U418 ( .A(G106GAT), .B(G78GAT), .ZN(n367) );
  XNOR2_X1 U419 ( .A(n367), .B(G148GAT), .ZN(n449) );
  XOR2_X1 U420 ( .A(n449), .B(KEYINPUT32), .Z(n369) );
  XNOR2_X1 U421 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n368) );
  XNOR2_X1 U422 ( .A(n368), .B(KEYINPUT74), .ZN(n381) );
  XOR2_X1 U423 ( .A(G64GAT), .B(KEYINPUT79), .Z(n373) );
  XNOR2_X1 U424 ( .A(G176GAT), .B(G204GAT), .ZN(n372) );
  XNOR2_X1 U425 ( .A(n373), .B(n372), .ZN(n438) );
  XOR2_X1 U426 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n375) );
  XNOR2_X1 U427 ( .A(G99GAT), .B(G92GAT), .ZN(n374) );
  XNOR2_X1 U428 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U429 ( .A(G85GAT), .B(n376), .Z(n403) );
  XNOR2_X1 U430 ( .A(n438), .B(n403), .ZN(n377) );
  XNOR2_X1 U431 ( .A(n378), .B(n377), .ZN(n581) );
  XOR2_X1 U432 ( .A(G8GAT), .B(G183GAT), .Z(n428) );
  XOR2_X1 U433 ( .A(G22GAT), .B(G155GAT), .Z(n453) );
  XOR2_X1 U434 ( .A(n428), .B(n453), .Z(n380) );
  XNOR2_X1 U435 ( .A(G211GAT), .B(G78GAT), .ZN(n379) );
  XNOR2_X1 U436 ( .A(n380), .B(n379), .ZN(n385) );
  XOR2_X1 U437 ( .A(n381), .B(KEYINPUT85), .Z(n383) );
  NAND2_X1 U438 ( .A1(G231GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U440 ( .A(n385), .B(n384), .Z(n387) );
  XNOR2_X1 U441 ( .A(G127GAT), .B(G71GAT), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n387), .B(n386), .ZN(n395) );
  XOR2_X1 U443 ( .A(KEYINPUT84), .B(G64GAT), .Z(n389) );
  XNOR2_X1 U444 ( .A(G1GAT), .B(G15GAT), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n389), .B(n388), .ZN(n393) );
  XOR2_X1 U446 ( .A(KEYINPUT86), .B(KEYINPUT12), .Z(n391) );
  XNOR2_X1 U447 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n390) );
  XNOR2_X1 U448 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U449 ( .A(n393), .B(n392), .Z(n394) );
  XNOR2_X1 U450 ( .A(n395), .B(n394), .ZN(n571) );
  INV_X1 U451 ( .A(n571), .ZN(n584) );
  XOR2_X1 U452 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n397) );
  XNOR2_X1 U453 ( .A(G134GAT), .B(G106GAT), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n410) );
  XOR2_X1 U455 ( .A(G36GAT), .B(G190GAT), .Z(n433) );
  XOR2_X1 U456 ( .A(KEYINPUT11), .B(KEYINPUT83), .Z(n399) );
  XNOR2_X1 U457 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n398) );
  XNOR2_X1 U458 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n433), .B(n400), .ZN(n402) );
  AND2_X1 U460 ( .A1(G232GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n404) );
  XNOR2_X1 U462 ( .A(n404), .B(n403), .ZN(n408) );
  XNOR2_X1 U463 ( .A(G50GAT), .B(KEYINPUT82), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n405), .B(G162GAT), .ZN(n445) );
  XOR2_X1 U465 ( .A(n406), .B(n445), .Z(n407) );
  XNOR2_X1 U466 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U467 ( .A(n410), .B(n409), .Z(n561) );
  XNOR2_X1 U468 ( .A(n561), .B(KEYINPUT36), .ZN(n588) );
  NOR2_X1 U469 ( .A1(n584), .A2(n588), .ZN(n413) );
  XOR2_X1 U470 ( .A(KEYINPUT45), .B(KEYINPUT114), .Z(n411) );
  XNOR2_X1 U471 ( .A(KEYINPUT65), .B(n411), .ZN(n412) );
  XNOR2_X1 U472 ( .A(n413), .B(n412), .ZN(n414) );
  NAND2_X1 U473 ( .A1(n581), .A2(n414), .ZN(n415) );
  XOR2_X1 U474 ( .A(KEYINPUT115), .B(n415), .Z(n416) );
  NOR2_X1 U475 ( .A1(n564), .A2(n416), .ZN(n426) );
  INV_X1 U476 ( .A(KEYINPUT41), .ZN(n417) );
  NOR2_X1 U477 ( .A1(n577), .A2(n508), .ZN(n420) );
  INV_X1 U478 ( .A(KEYINPUT46), .ZN(n419) );
  XNOR2_X1 U479 ( .A(n420), .B(n419), .ZN(n422) );
  INV_X1 U480 ( .A(n561), .ZN(n462) );
  NOR2_X1 U481 ( .A1(n462), .A2(n571), .ZN(n421) );
  NAND2_X1 U482 ( .A1(n422), .A2(n421), .ZN(n424) );
  XOR2_X1 U483 ( .A(KEYINPUT113), .B(KEYINPUT47), .Z(n423) );
  XNOR2_X1 U484 ( .A(n424), .B(n423), .ZN(n425) );
  NOR2_X1 U485 ( .A1(n426), .A2(n425), .ZN(n427) );
  XNOR2_X1 U486 ( .A(n427), .B(KEYINPUT48), .ZN(n536) );
  XOR2_X1 U487 ( .A(n428), .B(KEYINPUT101), .Z(n431) );
  XNOR2_X1 U488 ( .A(n429), .B(G92GAT), .ZN(n430) );
  XNOR2_X1 U489 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U490 ( .A(n433), .B(n432), .Z(n435) );
  NAND2_X1 U491 ( .A1(G226GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n440) );
  XOR2_X1 U493 ( .A(G211GAT), .B(KEYINPUT21), .Z(n437) );
  XNOR2_X1 U494 ( .A(G197GAT), .B(G218GAT), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n444) );
  XOR2_X1 U496 ( .A(n444), .B(n438), .Z(n439) );
  XNOR2_X1 U497 ( .A(n440), .B(n439), .ZN(n471) );
  NOR2_X1 U498 ( .A1(n536), .A2(n471), .ZN(n442) );
  NOR2_X1 U499 ( .A1(n524), .A2(n443), .ZN(n576) );
  XNOR2_X1 U500 ( .A(n445), .B(n444), .ZN(n458) );
  XOR2_X1 U501 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n447) );
  NAND2_X1 U502 ( .A1(G228GAT), .A2(G233GAT), .ZN(n446) );
  XNOR2_X1 U503 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U504 ( .A(n448), .B(KEYINPUT95), .Z(n452) );
  XNOR2_X1 U505 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U506 ( .A(n452), .B(n451), .ZN(n454) );
  XOR2_X1 U507 ( .A(n454), .B(n453), .Z(n456) );
  XNOR2_X1 U508 ( .A(G204GAT), .B(KEYINPUT23), .ZN(n455) );
  XNOR2_X1 U509 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U510 ( .A(n458), .B(n457), .ZN(n478) );
  NAND2_X1 U511 ( .A1(n576), .A2(n478), .ZN(n460) );
  NOR2_X1 U512 ( .A1(n538), .A2(n461), .ZN(n572) );
  NAND2_X1 U513 ( .A1(n572), .A2(n462), .ZN(n466) );
  XOR2_X1 U514 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n464) );
  INV_X1 U515 ( .A(G190GAT), .ZN(n463) );
  XOR2_X1 U516 ( .A(KEYINPUT103), .B(KEYINPUT34), .Z(n487) );
  NAND2_X1 U517 ( .A1(n564), .A2(n581), .ZN(n467) );
  XOR2_X1 U518 ( .A(KEYINPUT81), .B(n467), .Z(n498) );
  NAND2_X1 U519 ( .A1(n571), .A2(n561), .ZN(n468) );
  XNOR2_X1 U520 ( .A(n468), .B(KEYINPUT16), .ZN(n469) );
  XNOR2_X1 U521 ( .A(KEYINPUT87), .B(n469), .ZN(n485) );
  XOR2_X1 U522 ( .A(KEYINPUT27), .B(n471), .Z(n480) );
  NOR2_X1 U523 ( .A1(n529), .A2(n478), .ZN(n470) );
  XNOR2_X1 U524 ( .A(n470), .B(KEYINPUT26), .ZN(n575) );
  NAND2_X1 U525 ( .A1(n480), .A2(n575), .ZN(n475) );
  INV_X1 U526 ( .A(n471), .ZN(n526) );
  NAND2_X1 U527 ( .A1(n526), .A2(n529), .ZN(n472) );
  NAND2_X1 U528 ( .A1(n478), .A2(n472), .ZN(n473) );
  XOR2_X1 U529 ( .A(KEYINPUT25), .B(n473), .Z(n474) );
  NAND2_X1 U530 ( .A1(n475), .A2(n474), .ZN(n477) );
  INV_X1 U531 ( .A(n524), .ZN(n476) );
  NAND2_X1 U532 ( .A1(n477), .A2(n476), .ZN(n483) );
  XNOR2_X1 U533 ( .A(n478), .B(KEYINPUT67), .ZN(n479) );
  XNOR2_X1 U534 ( .A(n479), .B(KEYINPUT28), .ZN(n537) );
  NAND2_X1 U535 ( .A1(n524), .A2(n480), .ZN(n535) );
  NOR2_X1 U536 ( .A1(n537), .A2(n535), .ZN(n481) );
  NAND2_X1 U537 ( .A1(n538), .A2(n481), .ZN(n482) );
  NAND2_X1 U538 ( .A1(n483), .A2(n482), .ZN(n484) );
  XNOR2_X1 U539 ( .A(KEYINPUT102), .B(n484), .ZN(n495) );
  NAND2_X1 U540 ( .A1(n485), .A2(n495), .ZN(n510) );
  NOR2_X1 U541 ( .A1(n498), .A2(n510), .ZN(n493) );
  NAND2_X1 U542 ( .A1(n493), .A2(n524), .ZN(n486) );
  XNOR2_X1 U543 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U544 ( .A(G1GAT), .B(n488), .ZN(G1324GAT) );
  NAND2_X1 U545 ( .A1(n493), .A2(n526), .ZN(n489) );
  XNOR2_X1 U546 ( .A(n489), .B(KEYINPUT104), .ZN(n490) );
  XNOR2_X1 U547 ( .A(G8GAT), .B(n490), .ZN(G1325GAT) );
  XOR2_X1 U548 ( .A(G15GAT), .B(KEYINPUT35), .Z(n492) );
  NAND2_X1 U549 ( .A1(n493), .A2(n529), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n492), .B(n491), .ZN(G1326GAT) );
  NAND2_X1 U551 ( .A1(n493), .A2(n537), .ZN(n494) );
  XNOR2_X1 U552 ( .A(n494), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U553 ( .A(G29GAT), .B(KEYINPUT39), .Z(n501) );
  NAND2_X1 U554 ( .A1(n584), .A2(n495), .ZN(n496) );
  NOR2_X1 U555 ( .A1(n588), .A2(n496), .ZN(n497) );
  XNOR2_X1 U556 ( .A(KEYINPUT37), .B(n497), .ZN(n522) );
  NOR2_X1 U557 ( .A1(n498), .A2(n522), .ZN(n499) );
  XNOR2_X1 U558 ( .A(n499), .B(KEYINPUT38), .ZN(n506) );
  NAND2_X1 U559 ( .A1(n524), .A2(n506), .ZN(n500) );
  XNOR2_X1 U560 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  NAND2_X1 U561 ( .A1(n506), .A2(n526), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n502), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n504) );
  NAND2_X1 U564 ( .A1(n506), .A2(n529), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U566 ( .A(G43GAT), .B(n505), .ZN(G1330GAT) );
  NAND2_X1 U567 ( .A1(n506), .A2(n537), .ZN(n507) );
  XNOR2_X1 U568 ( .A(n507), .B(G50GAT), .ZN(G1331GAT) );
  INV_X1 U569 ( .A(n508), .ZN(n566) );
  NAND2_X1 U570 ( .A1(n566), .A2(n577), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n509), .B(KEYINPUT106), .ZN(n521) );
  NOR2_X1 U572 ( .A1(n521), .A2(n510), .ZN(n511) );
  XOR2_X1 U573 ( .A(KEYINPUT107), .B(n511), .Z(n518) );
  NAND2_X1 U574 ( .A1(n518), .A2(n524), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n512), .B(KEYINPUT42), .ZN(n513) );
  XNOR2_X1 U576 ( .A(G57GAT), .B(n513), .ZN(G1332GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n515) );
  NAND2_X1 U578 ( .A1(n518), .A2(n526), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U580 ( .A(G64GAT), .B(n516), .ZN(G1333GAT) );
  NAND2_X1 U581 ( .A1(n529), .A2(n518), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n517), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .Z(n520) );
  NAND2_X1 U584 ( .A1(n518), .A2(n537), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  NOR2_X1 U586 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(KEYINPUT110), .ZN(n531) );
  NAND2_X1 U588 ( .A1(n531), .A2(n524), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n525), .B(G85GAT), .ZN(G1336GAT) );
  XOR2_X1 U590 ( .A(G92GAT), .B(KEYINPUT111), .Z(n528) );
  NAND2_X1 U591 ( .A1(n526), .A2(n531), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(G1337GAT) );
  NAND2_X1 U593 ( .A1(n531), .A2(n529), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n533) );
  NAND2_X1 U596 ( .A1(n537), .A2(n531), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U598 ( .A(G106GAT), .B(n534), .Z(G1339GAT) );
  NOR2_X1 U599 ( .A1(n536), .A2(n535), .ZN(n551) );
  NOR2_X1 U600 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U601 ( .A1(n551), .A2(n539), .ZN(n540) );
  XNOR2_X1 U602 ( .A(KEYINPUT116), .B(n540), .ZN(n548) );
  NOR2_X1 U603 ( .A1(n548), .A2(n577), .ZN(n541) );
  XNOR2_X1 U604 ( .A(n541), .B(KEYINPUT117), .ZN(n542) );
  XNOR2_X1 U605 ( .A(G113GAT), .B(n542), .ZN(G1340GAT) );
  NOR2_X1 U606 ( .A1(n548), .A2(n508), .ZN(n544) );
  XNOR2_X1 U607 ( .A(KEYINPUT49), .B(KEYINPUT118), .ZN(n543) );
  XNOR2_X1 U608 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U609 ( .A(G120GAT), .B(n545), .ZN(G1341GAT) );
  NOR2_X1 U610 ( .A1(n584), .A2(n548), .ZN(n546) );
  XOR2_X1 U611 ( .A(KEYINPUT50), .B(n546), .Z(n547) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  XNOR2_X1 U613 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n550) );
  NOR2_X1 U614 ( .A1(n561), .A2(n548), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  NAND2_X1 U616 ( .A1(n551), .A2(n575), .ZN(n560) );
  NOR2_X1 U617 ( .A1(n577), .A2(n560), .ZN(n552) );
  XOR2_X1 U618 ( .A(G141GAT), .B(n552), .Z(G1344GAT) );
  NOR2_X1 U619 ( .A1(n560), .A2(n508), .ZN(n556) );
  XOR2_X1 U620 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n554) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(G1345GAT) );
  NOR2_X1 U624 ( .A1(n584), .A2(n560), .ZN(n558) );
  XNOR2_X1 U625 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U627 ( .A(G155GAT), .B(n559), .ZN(G1346GAT) );
  NOR2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U629 ( .A(KEYINPUT122), .B(n562), .Z(n563) );
  XNOR2_X1 U630 ( .A(G162GAT), .B(n563), .ZN(G1347GAT) );
  NAND2_X1 U631 ( .A1(n572), .A2(n564), .ZN(n565) );
  XNOR2_X1 U632 ( .A(G169GAT), .B(n565), .ZN(G1348GAT) );
  XOR2_X1 U633 ( .A(G176GAT), .B(KEYINPUT124), .Z(n568) );
  NAND2_X1 U634 ( .A1(n572), .A2(n566), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n570) );
  XNOR2_X1 U636 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n569) );
  XNOR2_X1 U637 ( .A(n570), .B(n569), .ZN(G1349GAT) );
  XOR2_X1 U638 ( .A(G183GAT), .B(KEYINPUT125), .Z(n574) );
  NAND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1350GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n587) );
  NOR2_X1 U642 ( .A1(n577), .A2(n587), .ZN(n579) );
  XNOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(n580), .ZN(G1352GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n587), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NOR2_X1 U649 ( .A1(n584), .A2(n587), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1354GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(n589), .Z(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

