

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U560 ( .A1(n634), .A2(n529), .ZN(n654) );
  OR2_X2 U561 ( .A1(G299), .A2(n751), .ZN(n525) );
  OR2_X1 U562 ( .A1(n805), .A2(n804), .ZN(n806) );
  OR2_X1 U563 ( .A1(n769), .A2(n768), .ZN(n770) );
  AND2_X2 U564 ( .A1(n539), .A2(G2104), .ZN(n899) );
  NOR2_X2 U565 ( .A1(n580), .A2(n579), .ZN(n980) );
  NOR2_X1 U566 ( .A1(G543), .A2(n529), .ZN(n526) );
  AND2_X1 U567 ( .A1(n994), .A2(n841), .ZN(n523) );
  OR2_X1 U568 ( .A1(n829), .A2(n828), .ZN(n524) );
  AND2_X1 U569 ( .A1(n752), .A2(G2072), .ZN(n746) );
  BUF_X1 U570 ( .A(n752), .Z(n762) );
  INV_X1 U571 ( .A(KEYINPUT33), .ZN(n830) );
  NOR2_X1 U572 ( .A1(n807), .A2(n806), .ZN(n822) );
  NOR2_X1 U573 ( .A1(n543), .A2(n542), .ZN(G160) );
  XOR2_X1 U574 ( .A(G543), .B(KEYINPUT0), .Z(n634) );
  NOR2_X2 U575 ( .A1(G651), .A2(n634), .ZN(n658) );
  NAND2_X1 U576 ( .A1(G53), .A2(n658), .ZN(n528) );
  INV_X1 U577 ( .A(G651), .ZN(n529) );
  XOR2_X1 U578 ( .A(KEYINPUT1), .B(n526), .Z(n661) );
  NAND2_X1 U579 ( .A1(G65), .A2(n661), .ZN(n527) );
  NAND2_X1 U580 ( .A1(n528), .A2(n527), .ZN(n533) );
  NOR2_X1 U581 ( .A1(G543), .A2(G651), .ZN(n653) );
  NAND2_X1 U582 ( .A1(G91), .A2(n653), .ZN(n531) );
  NAND2_X1 U583 ( .A1(G78), .A2(n654), .ZN(n530) );
  NAND2_X1 U584 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X1 U585 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U586 ( .A(n534), .B(KEYINPUT65), .ZN(G299) );
  NOR2_X1 U587 ( .A1(G2104), .A2(G2105), .ZN(n535) );
  XOR2_X2 U588 ( .A(KEYINPUT17), .B(n535), .Z(n898) );
  NAND2_X1 U589 ( .A1(n898), .A2(G137), .ZN(n538) );
  INV_X1 U590 ( .A(G2105), .ZN(n539) );
  NAND2_X1 U591 ( .A1(G101), .A2(n899), .ZN(n536) );
  XOR2_X1 U592 ( .A(KEYINPUT23), .B(n536), .Z(n537) );
  NAND2_X1 U593 ( .A1(n538), .A2(n537), .ZN(n543) );
  AND2_X1 U594 ( .A1(G2105), .A2(G2104), .ZN(n902) );
  NAND2_X1 U595 ( .A1(G113), .A2(n902), .ZN(n541) );
  NOR2_X2 U596 ( .A1(G2104), .A2(n539), .ZN(n903) );
  NAND2_X1 U597 ( .A1(G125), .A2(n903), .ZN(n540) );
  NAND2_X1 U598 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U599 ( .A1(n654), .A2(G76), .ZN(n544) );
  XNOR2_X1 U600 ( .A(KEYINPUT70), .B(n544), .ZN(n547) );
  NAND2_X1 U601 ( .A1(n653), .A2(G89), .ZN(n545) );
  XNOR2_X1 U602 ( .A(KEYINPUT4), .B(n545), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U604 ( .A(n548), .B(KEYINPUT5), .ZN(n553) );
  NAND2_X1 U605 ( .A1(G51), .A2(n658), .ZN(n550) );
  NAND2_X1 U606 ( .A1(G63), .A2(n661), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U608 ( .A(KEYINPUT6), .B(n551), .Z(n552) );
  NAND2_X1 U609 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U610 ( .A(n554), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U611 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U612 ( .A1(G102), .A2(n899), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G114), .A2(n902), .ZN(n556) );
  NAND2_X1 U614 ( .A1(G126), .A2(n903), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U616 ( .A1(n558), .A2(n557), .ZN(n560) );
  NAND2_X1 U617 ( .A1(G138), .A2(n898), .ZN(n559) );
  AND2_X1 U618 ( .A1(n560), .A2(n559), .ZN(G164) );
  XOR2_X1 U619 ( .A(G2443), .B(G2446), .Z(n562) );
  XNOR2_X1 U620 ( .A(G2427), .B(G2451), .ZN(n561) );
  XNOR2_X1 U621 ( .A(n562), .B(n561), .ZN(n568) );
  XOR2_X1 U622 ( .A(G2430), .B(G2454), .Z(n564) );
  INV_X1 U623 ( .A(G1341), .ZN(n935) );
  XOR2_X1 U624 ( .A(n935), .B(G1348), .Z(n563) );
  XNOR2_X1 U625 ( .A(n564), .B(n563), .ZN(n566) );
  XOR2_X1 U626 ( .A(G2435), .B(G2438), .Z(n565) );
  XNOR2_X1 U627 ( .A(n566), .B(n565), .ZN(n567) );
  XOR2_X1 U628 ( .A(n568), .B(n567), .Z(n569) );
  AND2_X1 U629 ( .A1(G14), .A2(n569), .ZN(G401) );
  AND2_X1 U630 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U631 ( .A(G132), .ZN(G219) );
  INV_X1 U632 ( .A(G82), .ZN(G220) );
  NAND2_X1 U633 ( .A1(G7), .A2(G661), .ZN(n570) );
  XOR2_X1 U634 ( .A(n570), .B(KEYINPUT10), .Z(n846) );
  NAND2_X1 U635 ( .A1(n846), .A2(G567), .ZN(n571) );
  XOR2_X1 U636 ( .A(KEYINPUT11), .B(n571), .Z(G234) );
  NAND2_X1 U637 ( .A1(n653), .A2(G81), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U639 ( .A1(G68), .A2(n654), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(KEYINPUT13), .ZN(n577) );
  NAND2_X1 U642 ( .A1(G43), .A2(n658), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n661), .A2(G56), .ZN(n578) );
  XOR2_X1 U645 ( .A(KEYINPUT14), .B(n578), .Z(n579) );
  NAND2_X1 U646 ( .A1(G860), .A2(n980), .ZN(n581) );
  XOR2_X1 U647 ( .A(KEYINPUT67), .B(n581), .Z(G153) );
  NAND2_X1 U648 ( .A1(G52), .A2(n658), .ZN(n583) );
  NAND2_X1 U649 ( .A1(G64), .A2(n661), .ZN(n582) );
  NAND2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n588) );
  NAND2_X1 U651 ( .A1(G90), .A2(n653), .ZN(n585) );
  NAND2_X1 U652 ( .A1(G77), .A2(n654), .ZN(n584) );
  NAND2_X1 U653 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U654 ( .A(KEYINPUT9), .B(n586), .Z(n587) );
  NOR2_X1 U655 ( .A1(n588), .A2(n587), .ZN(G171) );
  INV_X1 U656 ( .A(G171), .ZN(G301) );
  NAND2_X1 U657 ( .A1(G868), .A2(G301), .ZN(n603) );
  NAND2_X1 U658 ( .A1(G79), .A2(n654), .ZN(n590) );
  NAND2_X1 U659 ( .A1(G54), .A2(n658), .ZN(n589) );
  NAND2_X1 U660 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U661 ( .A(n591), .B(KEYINPUT68), .ZN(n595) );
  NAND2_X1 U662 ( .A1(G92), .A2(n653), .ZN(n593) );
  NAND2_X1 U663 ( .A1(G66), .A2(n661), .ZN(n592) );
  NAND2_X1 U664 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U665 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U666 ( .A(n596), .B(KEYINPUT15), .ZN(n597) );
  NAND2_X1 U667 ( .A1(KEYINPUT69), .A2(n597), .ZN(n601) );
  INV_X1 U668 ( .A(KEYINPUT69), .ZN(n599) );
  INV_X1 U669 ( .A(n597), .ZN(n598) );
  NAND2_X1 U670 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U671 ( .A1(n601), .A2(n600), .ZN(n667) );
  INV_X1 U672 ( .A(n667), .ZN(n985) );
  INV_X1 U673 ( .A(G868), .ZN(n610) );
  NAND2_X1 U674 ( .A1(n985), .A2(n610), .ZN(n602) );
  NAND2_X1 U675 ( .A1(n603), .A2(n602), .ZN(G284) );
  NAND2_X1 U676 ( .A1(G286), .A2(G868), .ZN(n605) );
  NAND2_X1 U677 ( .A1(G299), .A2(n610), .ZN(n604) );
  NAND2_X1 U678 ( .A1(n605), .A2(n604), .ZN(G297) );
  INV_X1 U679 ( .A(G860), .ZN(n854) );
  NAND2_X1 U680 ( .A1(n854), .A2(G559), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n606), .A2(n667), .ZN(n607) );
  XNOR2_X1 U682 ( .A(n607), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U683 ( .A1(n667), .A2(G868), .ZN(n608) );
  NOR2_X1 U684 ( .A1(G559), .A2(n608), .ZN(n609) );
  XNOR2_X1 U685 ( .A(n609), .B(KEYINPUT71), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n980), .A2(n610), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U688 ( .A(KEYINPUT72), .B(n613), .Z(G282) );
  NAND2_X1 U689 ( .A1(G111), .A2(n902), .ZN(n620) );
  NAND2_X1 U690 ( .A1(G135), .A2(n898), .ZN(n615) );
  NAND2_X1 U691 ( .A1(G99), .A2(n899), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n903), .A2(G123), .ZN(n616) );
  XOR2_X1 U694 ( .A(KEYINPUT18), .B(n616), .Z(n617) );
  NOR2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U697 ( .A(n621), .B(KEYINPUT73), .ZN(n1021) );
  XNOR2_X1 U698 ( .A(n1021), .B(G2096), .ZN(n622) );
  INV_X1 U699 ( .A(G2100), .ZN(n868) );
  NAND2_X1 U700 ( .A1(n622), .A2(n868), .ZN(G156) );
  NAND2_X1 U701 ( .A1(n654), .A2(G75), .ZN(n625) );
  NAND2_X1 U702 ( .A1(G88), .A2(n653), .ZN(n623) );
  XOR2_X1 U703 ( .A(KEYINPUT81), .B(n623), .Z(n624) );
  NAND2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U705 ( .A1(G50), .A2(n658), .ZN(n627) );
  NAND2_X1 U706 ( .A1(G62), .A2(n661), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U708 ( .A1(n629), .A2(n628), .ZN(G166) );
  NAND2_X1 U709 ( .A1(G49), .A2(n658), .ZN(n631) );
  NAND2_X1 U710 ( .A1(G74), .A2(G651), .ZN(n630) );
  NAND2_X1 U711 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U712 ( .A(KEYINPUT78), .B(n632), .ZN(n633) );
  NOR2_X1 U713 ( .A1(n661), .A2(n633), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n634), .A2(G87), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n636), .A2(n635), .ZN(G288) );
  NAND2_X1 U716 ( .A1(G86), .A2(n653), .ZN(n638) );
  NAND2_X1 U717 ( .A1(G61), .A2(n661), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U719 ( .A1(G73), .A2(n654), .ZN(n639) );
  XNOR2_X1 U720 ( .A(n639), .B(KEYINPUT2), .ZN(n640) );
  XNOR2_X1 U721 ( .A(n640), .B(KEYINPUT79), .ZN(n641) );
  NOR2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U723 ( .A(n643), .B(KEYINPUT80), .ZN(n645) );
  NAND2_X1 U724 ( .A1(G48), .A2(n658), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n645), .A2(n644), .ZN(G305) );
  NAND2_X1 U726 ( .A1(G85), .A2(n653), .ZN(n647) );
  NAND2_X1 U727 ( .A1(G72), .A2(n654), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U729 ( .A1(G47), .A2(n658), .ZN(n648) );
  XOR2_X1 U730 ( .A(KEYINPUT64), .B(n648), .Z(n649) );
  NOR2_X1 U731 ( .A1(n650), .A2(n649), .ZN(n652) );
  NAND2_X1 U732 ( .A1(n661), .A2(G60), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n652), .A2(n651), .ZN(G290) );
  NAND2_X1 U734 ( .A1(G93), .A2(n653), .ZN(n656) );
  NAND2_X1 U735 ( .A1(G80), .A2(n654), .ZN(n655) );
  NAND2_X1 U736 ( .A1(n656), .A2(n655), .ZN(n657) );
  XNOR2_X1 U737 ( .A(n657), .B(KEYINPUT75), .ZN(n660) );
  NAND2_X1 U738 ( .A1(G55), .A2(n658), .ZN(n659) );
  NAND2_X1 U739 ( .A1(n660), .A2(n659), .ZN(n664) );
  NAND2_X1 U740 ( .A1(n661), .A2(G67), .ZN(n662) );
  XOR2_X1 U741 ( .A(KEYINPUT76), .B(n662), .Z(n663) );
  NOR2_X1 U742 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U743 ( .A(KEYINPUT77), .B(n665), .Z(n853) );
  NOR2_X1 U744 ( .A1(G868), .A2(n853), .ZN(n666) );
  XNOR2_X1 U745 ( .A(n666), .B(KEYINPUT83), .ZN(n677) );
  NAND2_X1 U746 ( .A1(G559), .A2(n667), .ZN(n668) );
  XNOR2_X1 U747 ( .A(n668), .B(n980), .ZN(n855) );
  XOR2_X1 U748 ( .A(KEYINPUT82), .B(G166), .Z(n669) );
  XNOR2_X1 U749 ( .A(n669), .B(G288), .ZN(n670) );
  XNOR2_X1 U750 ( .A(KEYINPUT19), .B(n670), .ZN(n672) );
  XNOR2_X1 U751 ( .A(G305), .B(n853), .ZN(n671) );
  XNOR2_X1 U752 ( .A(n672), .B(n671), .ZN(n673) );
  XOR2_X1 U753 ( .A(n673), .B(G290), .Z(n674) );
  XNOR2_X1 U754 ( .A(G299), .B(n674), .ZN(n920) );
  XNOR2_X1 U755 ( .A(n855), .B(n920), .ZN(n675) );
  NAND2_X1 U756 ( .A1(G868), .A2(n675), .ZN(n676) );
  NAND2_X1 U757 ( .A1(n677), .A2(n676), .ZN(G295) );
  NAND2_X1 U758 ( .A1(G2084), .A2(G2078), .ZN(n678) );
  XOR2_X1 U759 ( .A(KEYINPUT20), .B(n678), .Z(n679) );
  NAND2_X1 U760 ( .A1(G2090), .A2(n679), .ZN(n680) );
  XNOR2_X1 U761 ( .A(KEYINPUT21), .B(n680), .ZN(n681) );
  NAND2_X1 U762 ( .A1(n681), .A2(G2072), .ZN(G158) );
  XOR2_X1 U763 ( .A(KEYINPUT66), .B(G57), .Z(G237) );
  XNOR2_X1 U764 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U765 ( .A1(G108), .A2(G120), .ZN(n682) );
  NOR2_X1 U766 ( .A1(G237), .A2(n682), .ZN(n683) );
  NAND2_X1 U767 ( .A1(G69), .A2(n683), .ZN(n851) );
  NAND2_X1 U768 ( .A1(n851), .A2(G567), .ZN(n688) );
  NOR2_X1 U769 ( .A1(G220), .A2(G219), .ZN(n684) );
  XOR2_X1 U770 ( .A(KEYINPUT22), .B(n684), .Z(n685) );
  NOR2_X1 U771 ( .A1(G218), .A2(n685), .ZN(n686) );
  NAND2_X1 U772 ( .A1(G96), .A2(n686), .ZN(n852) );
  NAND2_X1 U773 ( .A1(n852), .A2(G2106), .ZN(n687) );
  NAND2_X1 U774 ( .A1(n688), .A2(n687), .ZN(n931) );
  NAND2_X1 U775 ( .A1(G483), .A2(G661), .ZN(n689) );
  NOR2_X1 U776 ( .A1(n931), .A2(n689), .ZN(n850) );
  NAND2_X1 U777 ( .A1(n850), .A2(G36), .ZN(G176) );
  INV_X1 U778 ( .A(G166), .ZN(G303) );
  NAND2_X1 U779 ( .A1(G131), .A2(n898), .ZN(n691) );
  NAND2_X1 U780 ( .A1(G95), .A2(n899), .ZN(n690) );
  NAND2_X1 U781 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U782 ( .A(KEYINPUT89), .B(n692), .ZN(n697) );
  NAND2_X1 U783 ( .A1(G107), .A2(n902), .ZN(n694) );
  NAND2_X1 U784 ( .A1(G119), .A2(n903), .ZN(n693) );
  NAND2_X1 U785 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U786 ( .A(KEYINPUT88), .B(n695), .Z(n696) );
  NAND2_X1 U787 ( .A1(n697), .A2(n696), .ZN(n909) );
  NAND2_X1 U788 ( .A1(G1991), .A2(n909), .ZN(n698) );
  XOR2_X1 U789 ( .A(KEYINPUT90), .B(n698), .Z(n711) );
  NAND2_X1 U790 ( .A1(n898), .A2(G141), .ZN(n699) );
  XOR2_X1 U791 ( .A(KEYINPUT94), .B(n699), .Z(n709) );
  NAND2_X1 U792 ( .A1(G117), .A2(n902), .ZN(n700) );
  XNOR2_X1 U793 ( .A(n700), .B(KEYINPUT92), .ZN(n703) );
  NAND2_X1 U794 ( .A1(G129), .A2(n903), .ZN(n701) );
  XOR2_X1 U795 ( .A(KEYINPUT91), .B(n701), .Z(n702) );
  NAND2_X1 U796 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U797 ( .A1(n899), .A2(G105), .ZN(n704) );
  XOR2_X1 U798 ( .A(KEYINPUT38), .B(n704), .Z(n705) );
  NOR2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U800 ( .A(n707), .B(KEYINPUT93), .ZN(n708) );
  NOR2_X1 U801 ( .A1(n709), .A2(n708), .ZN(n885) );
  INV_X1 U802 ( .A(G1996), .ZN(n958) );
  NOR2_X1 U803 ( .A1(n885), .A2(n958), .ZN(n710) );
  NOR2_X1 U804 ( .A1(n711), .A2(n710), .ZN(n808) );
  XOR2_X1 U805 ( .A(G1986), .B(G290), .Z(n987) );
  NAND2_X1 U806 ( .A1(n808), .A2(n987), .ZN(n713) );
  NOR2_X1 U807 ( .A1(G164), .A2(G1384), .ZN(n712) );
  INV_X1 U808 ( .A(n712), .ZN(n728) );
  NAND2_X1 U809 ( .A1(G160), .A2(G40), .ZN(n727) );
  NOR2_X1 U810 ( .A1(n712), .A2(n727), .ZN(n819) );
  NAND2_X1 U811 ( .A1(n713), .A2(n819), .ZN(n839) );
  INV_X1 U812 ( .A(n839), .ZN(n807) );
  NAND2_X1 U813 ( .A1(n899), .A2(G104), .ZN(n714) );
  XNOR2_X1 U814 ( .A(n714), .B(KEYINPUT84), .ZN(n716) );
  NAND2_X1 U815 ( .A1(G140), .A2(n898), .ZN(n715) );
  NAND2_X1 U816 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U817 ( .A(KEYINPUT34), .B(n717), .ZN(n723) );
  NAND2_X1 U818 ( .A1(n902), .A2(G116), .ZN(n718) );
  XOR2_X1 U819 ( .A(KEYINPUT85), .B(n718), .Z(n720) );
  NAND2_X1 U820 ( .A1(n903), .A2(G128), .ZN(n719) );
  NAND2_X1 U821 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U822 ( .A(n721), .B(KEYINPUT35), .Z(n722) );
  NOR2_X1 U823 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U824 ( .A(KEYINPUT36), .B(n724), .Z(n725) );
  XOR2_X1 U825 ( .A(KEYINPUT86), .B(n725), .Z(n914) );
  XNOR2_X1 U826 ( .A(G2067), .B(KEYINPUT37), .ZN(n816) );
  OR2_X1 U827 ( .A1(n914), .A2(n816), .ZN(n726) );
  XNOR2_X1 U828 ( .A(n726), .B(KEYINPUT87), .ZN(n1019) );
  NAND2_X1 U829 ( .A1(n819), .A2(n1019), .ZN(n837) );
  INV_X1 U830 ( .A(n837), .ZN(n805) );
  NOR2_X4 U831 ( .A1(n728), .A2(n727), .ZN(n752) );
  INV_X1 U832 ( .A(n752), .ZN(n780) );
  NAND2_X1 U833 ( .A1(G8), .A2(n780), .ZN(n836) );
  NOR2_X1 U834 ( .A1(G1981), .A2(G305), .ZN(n729) );
  XNOR2_X1 U835 ( .A(n729), .B(KEYINPUT24), .ZN(n730) );
  XNOR2_X1 U836 ( .A(n730), .B(KEYINPUT95), .ZN(n731) );
  OR2_X1 U837 ( .A1(n836), .A2(n731), .ZN(n803) );
  NOR2_X1 U838 ( .A1(G1966), .A2(n836), .ZN(n795) );
  INV_X1 U839 ( .A(G2084), .ZN(n732) );
  AND2_X1 U840 ( .A1(n732), .A2(n752), .ZN(n733) );
  XNOR2_X1 U841 ( .A(KEYINPUT96), .B(n733), .ZN(n791) );
  INV_X1 U842 ( .A(n791), .ZN(n734) );
  NAND2_X1 U843 ( .A1(G8), .A2(n734), .ZN(n735) );
  NOR2_X1 U844 ( .A1(n795), .A2(n735), .ZN(n736) );
  XOR2_X1 U845 ( .A(KEYINPUT30), .B(n736), .Z(n737) );
  NOR2_X1 U846 ( .A1(G168), .A2(n737), .ZN(n738) );
  XOR2_X1 U847 ( .A(KEYINPUT102), .B(n738), .Z(n743) );
  XNOR2_X1 U848 ( .A(G2078), .B(KEYINPUT25), .ZN(n962) );
  NAND2_X1 U849 ( .A1(n762), .A2(n962), .ZN(n739) );
  XNOR2_X1 U850 ( .A(n739), .B(KEYINPUT97), .ZN(n741) );
  NOR2_X1 U851 ( .A1(n762), .A2(G1961), .ZN(n740) );
  NOR2_X1 U852 ( .A1(n741), .A2(n740), .ZN(n775) );
  NAND2_X1 U853 ( .A1(n775), .A2(G301), .ZN(n742) );
  NAND2_X1 U854 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U855 ( .A(n744), .B(KEYINPUT31), .ZN(n779) );
  XNOR2_X1 U856 ( .A(KEYINPUT98), .B(KEYINPUT27), .ZN(n745) );
  XNOR2_X1 U857 ( .A(n746), .B(n745), .ZN(n748) );
  NAND2_X1 U858 ( .A1(n780), .A2(G1956), .ZN(n747) );
  NAND2_X1 U859 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U860 ( .A(KEYINPUT99), .B(n749), .Z(n751) );
  NAND2_X1 U861 ( .A1(G299), .A2(n751), .ZN(n750) );
  XOR2_X1 U862 ( .A(KEYINPUT28), .B(n750), .Z(n773) );
  NAND2_X1 U863 ( .A1(n780), .A2(G1341), .ZN(n757) );
  INV_X1 U864 ( .A(KEYINPUT26), .ZN(n758) );
  NAND2_X1 U865 ( .A1(G1996), .A2(n752), .ZN(n753) );
  XOR2_X1 U866 ( .A(n758), .B(n753), .Z(n754) );
  NAND2_X1 U867 ( .A1(n757), .A2(n754), .ZN(n755) );
  NAND2_X1 U868 ( .A1(n755), .A2(KEYINPUT100), .ZN(n756) );
  NAND2_X1 U869 ( .A1(n756), .A2(n980), .ZN(n761) );
  NOR2_X1 U870 ( .A1(n758), .A2(n757), .ZN(n759) );
  NOR2_X1 U871 ( .A1(KEYINPUT100), .A2(n759), .ZN(n760) );
  NOR2_X1 U872 ( .A1(n761), .A2(n760), .ZN(n766) );
  NAND2_X1 U873 ( .A1(G1348), .A2(n780), .ZN(n764) );
  NAND2_X1 U874 ( .A1(G2067), .A2(n762), .ZN(n763) );
  NAND2_X1 U875 ( .A1(n764), .A2(n763), .ZN(n767) );
  NOR2_X1 U876 ( .A1(n985), .A2(n767), .ZN(n765) );
  NOR2_X1 U877 ( .A1(n766), .A2(n765), .ZN(n769) );
  AND2_X1 U878 ( .A1(n985), .A2(n767), .ZN(n768) );
  NAND2_X1 U879 ( .A1(n525), .A2(n770), .ZN(n771) );
  XNOR2_X1 U880 ( .A(n771), .B(KEYINPUT101), .ZN(n772) );
  NOR2_X1 U881 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U882 ( .A(n774), .B(KEYINPUT29), .ZN(n777) );
  OR2_X1 U883 ( .A1(G301), .A2(n775), .ZN(n776) );
  NAND2_X1 U884 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U885 ( .A1(n779), .A2(n778), .ZN(n790) );
  NAND2_X1 U886 ( .A1(n790), .A2(G286), .ZN(n786) );
  NOR2_X1 U887 ( .A1(G1971), .A2(n836), .ZN(n782) );
  NOR2_X1 U888 ( .A1(G2090), .A2(n780), .ZN(n781) );
  NOR2_X1 U889 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U890 ( .A1(n783), .A2(G303), .ZN(n784) );
  XNOR2_X1 U891 ( .A(n784), .B(KEYINPUT104), .ZN(n785) );
  NAND2_X1 U892 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U893 ( .A1(n787), .A2(G8), .ZN(n788) );
  XOR2_X1 U894 ( .A(KEYINPUT32), .B(n788), .Z(n797) );
  INV_X1 U895 ( .A(KEYINPUT103), .ZN(n789) );
  XNOR2_X1 U896 ( .A(n790), .B(n789), .ZN(n793) );
  NAND2_X1 U897 ( .A1(G8), .A2(n791), .ZN(n792) );
  NAND2_X1 U898 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U899 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X2 U900 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U901 ( .A(n798), .B(KEYINPUT105), .ZN(n825) );
  NOR2_X1 U902 ( .A1(G2090), .A2(G303), .ZN(n799) );
  NAND2_X1 U903 ( .A1(G8), .A2(n799), .ZN(n800) );
  NAND2_X1 U904 ( .A1(n825), .A2(n800), .ZN(n801) );
  NAND2_X1 U905 ( .A1(n801), .A2(n836), .ZN(n802) );
  AND2_X1 U906 ( .A1(n803), .A2(n802), .ZN(n804) );
  AND2_X1 U907 ( .A1(n958), .A2(n885), .ZN(n1008) );
  INV_X1 U908 ( .A(n808), .ZN(n1015) );
  NOR2_X1 U909 ( .A1(G1991), .A2(n909), .ZN(n1024) );
  NOR2_X1 U910 ( .A1(G1986), .A2(G290), .ZN(n809) );
  NOR2_X1 U911 ( .A1(n1024), .A2(n809), .ZN(n810) );
  XNOR2_X1 U912 ( .A(n810), .B(KEYINPUT108), .ZN(n811) );
  NOR2_X1 U913 ( .A1(n1015), .A2(n811), .ZN(n812) );
  NOR2_X1 U914 ( .A1(n1008), .A2(n812), .ZN(n813) );
  XOR2_X1 U915 ( .A(KEYINPUT39), .B(n813), .Z(n814) );
  XNOR2_X1 U916 ( .A(n814), .B(KEYINPUT109), .ZN(n815) );
  NAND2_X1 U917 ( .A1(n815), .A2(n837), .ZN(n817) );
  NAND2_X1 U918 ( .A1(n914), .A2(n816), .ZN(n1022) );
  NAND2_X1 U919 ( .A1(n817), .A2(n1022), .ZN(n818) );
  XNOR2_X1 U920 ( .A(KEYINPUT110), .B(n818), .ZN(n820) );
  AND2_X1 U921 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U922 ( .A1(n822), .A2(n821), .ZN(n844) );
  NOR2_X1 U923 ( .A1(G1976), .A2(G288), .ZN(n982) );
  NOR2_X1 U924 ( .A1(G1971), .A2(G303), .ZN(n823) );
  NOR2_X1 U925 ( .A1(n982), .A2(n823), .ZN(n824) );
  NAND2_X1 U926 ( .A1(n825), .A2(n824), .ZN(n826) );
  NAND2_X1 U927 ( .A1(G1976), .A2(G288), .ZN(n983) );
  NAND2_X1 U928 ( .A1(n826), .A2(n983), .ZN(n827) );
  XNOR2_X1 U929 ( .A(n827), .B(KEYINPUT106), .ZN(n829) );
  OR2_X1 U930 ( .A1(n836), .A2(KEYINPUT107), .ZN(n828) );
  NAND2_X1 U931 ( .A1(n524), .A2(n830), .ZN(n842) );
  XOR2_X1 U932 ( .A(G1981), .B(G305), .Z(n994) );
  INV_X1 U933 ( .A(KEYINPUT107), .ZN(n832) );
  NAND2_X1 U934 ( .A1(n982), .A2(KEYINPUT33), .ZN(n831) );
  NAND2_X1 U935 ( .A1(n832), .A2(n831), .ZN(n834) );
  NAND2_X1 U936 ( .A1(n982), .A2(KEYINPUT107), .ZN(n833) );
  NAND2_X1 U937 ( .A1(n834), .A2(n833), .ZN(n835) );
  OR2_X1 U938 ( .A1(n836), .A2(n835), .ZN(n838) );
  AND2_X1 U939 ( .A1(n838), .A2(n837), .ZN(n840) );
  AND2_X1 U940 ( .A1(n840), .A2(n839), .ZN(n841) );
  NAND2_X1 U941 ( .A1(n842), .A2(n523), .ZN(n843) );
  NAND2_X1 U942 ( .A1(n844), .A2(n843), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n845), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U944 ( .A1(G2106), .A2(n846), .ZN(G217) );
  INV_X1 U945 ( .A(n846), .ZN(G223) );
  NAND2_X1 U946 ( .A1(G15), .A2(G2), .ZN(n847) );
  XNOR2_X1 U947 ( .A(KEYINPUT111), .B(n847), .ZN(n848) );
  NAND2_X1 U948 ( .A1(n848), .A2(G661), .ZN(G259) );
  NAND2_X1 U949 ( .A1(G3), .A2(G1), .ZN(n849) );
  NAND2_X1 U950 ( .A1(n850), .A2(n849), .ZN(G188) );
  XOR2_X1 U951 ( .A(G96), .B(KEYINPUT112), .Z(G221) );
  NOR2_X1 U952 ( .A1(n852), .A2(n851), .ZN(G325) );
  XNOR2_X1 U953 ( .A(KEYINPUT113), .B(G325), .ZN(G261) );
  XOR2_X1 U955 ( .A(n853), .B(KEYINPUT74), .Z(n857) );
  NAND2_X1 U956 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(G145) );
  INV_X1 U958 ( .A(G120), .ZN(G236) );
  INV_X1 U959 ( .A(G108), .ZN(G238) );
  INV_X1 U960 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U961 ( .A(G1971), .B(G2474), .ZN(n867) );
  XOR2_X1 U962 ( .A(G1976), .B(G1956), .Z(n859) );
  XNOR2_X1 U963 ( .A(G1986), .B(G1961), .ZN(n858) );
  XNOR2_X1 U964 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U965 ( .A(G1981), .B(G1966), .Z(n861) );
  XOR2_X1 U966 ( .A(n958), .B(G1991), .Z(n860) );
  XNOR2_X1 U967 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U968 ( .A(n863), .B(n862), .Z(n865) );
  XNOR2_X1 U969 ( .A(KEYINPUT114), .B(KEYINPUT41), .ZN(n864) );
  XNOR2_X1 U970 ( .A(n865), .B(n864), .ZN(n866) );
  XNOR2_X1 U971 ( .A(n867), .B(n866), .ZN(G229) );
  XNOR2_X1 U972 ( .A(n868), .B(G2096), .ZN(n870) );
  XNOR2_X1 U973 ( .A(KEYINPUT42), .B(G2678), .ZN(n869) );
  XNOR2_X1 U974 ( .A(n870), .B(n869), .ZN(n875) );
  INV_X1 U975 ( .A(G2072), .ZN(n871) );
  XNOR2_X1 U976 ( .A(KEYINPUT43), .B(n871), .ZN(n873) );
  XNOR2_X1 U977 ( .A(G2067), .B(G2090), .ZN(n872) );
  XNOR2_X1 U978 ( .A(n873), .B(n872), .ZN(n874) );
  XOR2_X1 U979 ( .A(n875), .B(n874), .Z(n877) );
  XNOR2_X1 U980 ( .A(G2084), .B(G2078), .ZN(n876) );
  XNOR2_X1 U981 ( .A(n877), .B(n876), .ZN(G227) );
  NAND2_X1 U982 ( .A1(G124), .A2(n903), .ZN(n878) );
  XNOR2_X1 U983 ( .A(n878), .B(KEYINPUT44), .ZN(n880) );
  NAND2_X1 U984 ( .A1(n902), .A2(G112), .ZN(n879) );
  NAND2_X1 U985 ( .A1(n880), .A2(n879), .ZN(n884) );
  NAND2_X1 U986 ( .A1(G136), .A2(n898), .ZN(n882) );
  NAND2_X1 U987 ( .A1(G100), .A2(n899), .ZN(n881) );
  NAND2_X1 U988 ( .A1(n882), .A2(n881), .ZN(n883) );
  NOR2_X1 U989 ( .A1(n884), .A2(n883), .ZN(G162) );
  XOR2_X1 U990 ( .A(n1021), .B(G162), .Z(n887) );
  XNOR2_X1 U991 ( .A(G160), .B(n885), .ZN(n886) );
  XNOR2_X1 U992 ( .A(n887), .B(n886), .ZN(n897) );
  NAND2_X1 U993 ( .A1(G118), .A2(n902), .ZN(n889) );
  NAND2_X1 U994 ( .A1(G130), .A2(n903), .ZN(n888) );
  NAND2_X1 U995 ( .A1(n889), .A2(n888), .ZN(n895) );
  NAND2_X1 U996 ( .A1(n898), .A2(G142), .ZN(n890) );
  XOR2_X1 U997 ( .A(KEYINPUT115), .B(n890), .Z(n892) );
  NAND2_X1 U998 ( .A1(n899), .A2(G106), .ZN(n891) );
  NAND2_X1 U999 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U1000 ( .A(n893), .B(KEYINPUT45), .Z(n894) );
  NOR2_X1 U1001 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U1002 ( .A(n897), .B(n896), .Z(n913) );
  XNOR2_X1 U1003 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n911) );
  NAND2_X1 U1004 ( .A1(G139), .A2(n898), .ZN(n901) );
  NAND2_X1 U1005 ( .A1(G103), .A2(n899), .ZN(n900) );
  NAND2_X1 U1006 ( .A1(n901), .A2(n900), .ZN(n908) );
  NAND2_X1 U1007 ( .A1(G115), .A2(n902), .ZN(n905) );
  NAND2_X1 U1008 ( .A1(G127), .A2(n903), .ZN(n904) );
  NAND2_X1 U1009 ( .A1(n905), .A2(n904), .ZN(n906) );
  XOR2_X1 U1010 ( .A(KEYINPUT47), .B(n906), .Z(n907) );
  NOR2_X1 U1011 ( .A1(n908), .A2(n907), .ZN(n1010) );
  XNOR2_X1 U1012 ( .A(n909), .B(n1010), .ZN(n910) );
  XNOR2_X1 U1013 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1014 ( .A(n913), .B(n912), .Z(n916) );
  XNOR2_X1 U1015 ( .A(G164), .B(n914), .ZN(n915) );
  XNOR2_X1 U1016 ( .A(n916), .B(n915), .ZN(n917) );
  NOR2_X1 U1017 ( .A1(G37), .A2(n917), .ZN(G395) );
  XNOR2_X1 U1018 ( .A(KEYINPUT116), .B(n985), .ZN(n919) );
  XOR2_X1 U1019 ( .A(G301), .B(n980), .Z(n918) );
  XNOR2_X1 U1020 ( .A(n919), .B(n918), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(n921), .B(n920), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(n922), .B(G286), .ZN(n923) );
  NOR2_X1 U1023 ( .A1(G37), .A2(n923), .ZN(G397) );
  XNOR2_X1 U1024 ( .A(KEYINPUT49), .B(KEYINPUT118), .ZN(n925) );
  NOR2_X1 U1025 ( .A1(G229), .A2(G227), .ZN(n924) );
  XNOR2_X1 U1026 ( .A(n925), .B(n924), .ZN(n928) );
  NOR2_X1 U1027 ( .A1(G401), .A2(n931), .ZN(n926) );
  XNOR2_X1 U1028 ( .A(KEYINPUT117), .B(n926), .ZN(n927) );
  NOR2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n930) );
  NOR2_X1 U1030 ( .A1(G395), .A2(G397), .ZN(n929) );
  NAND2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(G225) );
  INV_X1 U1032 ( .A(G225), .ZN(G308) );
  INV_X1 U1033 ( .A(n931), .ZN(G319) );
  XOR2_X1 U1034 ( .A(G1956), .B(G20), .Z(n934) );
  XNOR2_X1 U1035 ( .A(G6), .B(KEYINPUT123), .ZN(n932) );
  XNOR2_X1 U1036 ( .A(n932), .B(G1981), .ZN(n933) );
  NAND2_X1 U1037 ( .A1(n934), .A2(n933), .ZN(n937) );
  XOR2_X1 U1038 ( .A(G19), .B(n935), .Z(n936) );
  NOR2_X1 U1039 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1040 ( .A(KEYINPUT124), .B(n938), .ZN(n941) );
  XNOR2_X1 U1041 ( .A(G1348), .B(KEYINPUT59), .ZN(n939) );
  XNOR2_X1 U1042 ( .A(n939), .B(G4), .ZN(n940) );
  NAND2_X1 U1043 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1044 ( .A(n942), .B(KEYINPUT60), .ZN(n943) );
  XNOR2_X1 U1045 ( .A(KEYINPUT125), .B(n943), .ZN(n947) );
  XNOR2_X1 U1046 ( .A(G1966), .B(G21), .ZN(n945) );
  XNOR2_X1 U1047 ( .A(G5), .B(G1961), .ZN(n944) );
  NOR2_X1 U1048 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1049 ( .A1(n947), .A2(n946), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(G1971), .B(G22), .ZN(n949) );
  XNOR2_X1 U1051 ( .A(G23), .B(G1976), .ZN(n948) );
  NOR2_X1 U1052 ( .A1(n949), .A2(n948), .ZN(n951) );
  XOR2_X1 U1053 ( .A(G1986), .B(G24), .Z(n950) );
  NAND2_X1 U1054 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1055 ( .A(KEYINPUT58), .B(n952), .ZN(n953) );
  NOR2_X1 U1056 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1057 ( .A(n955), .B(KEYINPUT126), .Z(n956) );
  XNOR2_X1 U1058 ( .A(KEYINPUT61), .B(n956), .ZN(n957) );
  NOR2_X1 U1059 ( .A1(G16), .A2(n957), .ZN(n1036) );
  XNOR2_X1 U1060 ( .A(G2090), .B(G35), .ZN(n972) );
  XNOR2_X1 U1061 ( .A(G2067), .B(G26), .ZN(n960) );
  XOR2_X1 U1062 ( .A(G32), .B(n958), .Z(n959) );
  NOR2_X1 U1063 ( .A1(n960), .A2(n959), .ZN(n967) );
  XOR2_X1 U1064 ( .A(G33), .B(G2072), .Z(n961) );
  NAND2_X1 U1065 ( .A1(n961), .A2(G28), .ZN(n965) );
  XOR2_X1 U1066 ( .A(G27), .B(n962), .Z(n963) );
  XNOR2_X1 U1067 ( .A(KEYINPUT120), .B(n963), .ZN(n964) );
  NOR2_X1 U1068 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1069 ( .A1(n967), .A2(n966), .ZN(n969) );
  XNOR2_X1 U1070 ( .A(G25), .B(G1991), .ZN(n968) );
  NOR2_X1 U1071 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1072 ( .A(KEYINPUT53), .B(n970), .ZN(n971) );
  NOR2_X1 U1073 ( .A1(n972), .A2(n971), .ZN(n975) );
  XOR2_X1 U1074 ( .A(G2084), .B(G34), .Z(n973) );
  XNOR2_X1 U1075 ( .A(KEYINPUT54), .B(n973), .ZN(n974) );
  NAND2_X1 U1076 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1077 ( .A(KEYINPUT55), .B(n976), .Z(n978) );
  INV_X1 U1078 ( .A(G29), .ZN(n977) );
  NAND2_X1 U1079 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1080 ( .A1(G11), .A2(n979), .ZN(n1006) );
  XOR2_X1 U1081 ( .A(KEYINPUT56), .B(G16), .Z(n1004) );
  XOR2_X1 U1082 ( .A(n980), .B(G1341), .Z(n981) );
  NOR2_X1 U1083 ( .A1(n982), .A2(n981), .ZN(n984) );
  NAND2_X1 U1084 ( .A1(n984), .A2(n983), .ZN(n1002) );
  XOR2_X1 U1085 ( .A(n985), .B(G1348), .Z(n1000) );
  XOR2_X1 U1086 ( .A(G1971), .B(G303), .Z(n986) );
  XNOR2_X1 U1087 ( .A(n986), .B(KEYINPUT122), .ZN(n992) );
  XOR2_X1 U1088 ( .A(G301), .B(G1961), .Z(n988) );
  NAND2_X1 U1089 ( .A1(n988), .A2(n987), .ZN(n990) );
  XNOR2_X1 U1090 ( .A(G1956), .B(G299), .ZN(n989) );
  NOR2_X1 U1091 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1092 ( .A1(n992), .A2(n991), .ZN(n998) );
  XOR2_X1 U1093 ( .A(G1966), .B(G168), .Z(n993) );
  XNOR2_X1 U1094 ( .A(KEYINPUT121), .B(n993), .ZN(n995) );
  NAND2_X1 U1095 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1096 ( .A(KEYINPUT57), .B(n996), .Z(n997) );
  NOR2_X1 U1097 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1098 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NOR2_X1 U1099 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1100 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1101 ( .A1(n1006), .A2(n1005), .ZN(n1034) );
  XOR2_X1 U1102 ( .A(G2090), .B(G162), .Z(n1007) );
  NOR2_X1 U1103 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1104 ( .A(KEYINPUT51), .B(n1009), .Z(n1017) );
  XOR2_X1 U1105 ( .A(G164), .B(G2078), .Z(n1012) );
  XOR2_X1 U1106 ( .A(G2072), .B(n1010), .Z(n1011) );
  NOR2_X1 U1107 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1108 ( .A(KEYINPUT50), .B(n1013), .Z(n1014) );
  NOR2_X1 U1109 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1110 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1111 ( .A1(n1019), .A2(n1018), .ZN(n1027) );
  XOR2_X1 U1112 ( .A(G2084), .B(G160), .Z(n1020) );
  NOR2_X1 U1113 ( .A1(n1021), .A2(n1020), .ZN(n1023) );
  NAND2_X1 U1114 ( .A1(n1023), .A2(n1022), .ZN(n1025) );
  NOR2_X1 U1115 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1116 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1117 ( .A(KEYINPUT52), .B(n1028), .ZN(n1029) );
  XNOR2_X1 U1118 ( .A(KEYINPUT119), .B(n1029), .ZN(n1031) );
  INV_X1 U1119 ( .A(KEYINPUT55), .ZN(n1030) );
  NAND2_X1 U1120 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1121 ( .A1(n1032), .A2(G29), .ZN(n1033) );
  NAND2_X1 U1122 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  NOR2_X1 U1123 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  XOR2_X1 U1124 ( .A(KEYINPUT127), .B(n1037), .Z(n1038) );
  XOR2_X1 U1125 ( .A(KEYINPUT62), .B(n1038), .Z(G150) );
  INV_X1 U1126 ( .A(G150), .ZN(G311) );
endmodule

