//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n797, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G128), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT23), .A3(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G128), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT24), .B(G110), .Z(new_n194));
  XNOR2_X1  g008(.A(G119), .B(G128), .ZN(new_n195));
  OAI22_X1  g009(.A1(new_n193), .A2(G110), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT16), .ZN(new_n197));
  INV_X1    g011(.A(G140), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G125), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(G125), .ZN(new_n200));
  INV_X1    g014(.A(G125), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G140), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  OAI211_X1 g017(.A(G146), .B(new_n199), .C1(new_n203), .C2(new_n197), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n200), .A2(new_n202), .A3(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n196), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n199), .B1(new_n203), .B2(new_n197), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(new_n205), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(new_n204), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n194), .A2(new_n195), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n193), .A2(G110), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT79), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n213), .B(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n207), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT80), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT22), .B(G137), .ZN(new_n218));
  INV_X1    g032(.A(G221), .ZN(new_n219));
  INV_X1    g033(.A(G234), .ZN(new_n220));
  NOR3_X1   g034(.A1(new_n219), .A2(new_n220), .A3(G953), .ZN(new_n221));
  XOR2_X1   g035(.A(new_n218), .B(new_n221), .Z(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT80), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n224), .B(new_n207), .C1(new_n212), .C2(new_n215), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n217), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n216), .A2(KEYINPUT80), .A3(new_n222), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XOR2_X1   g042(.A(new_n228), .B(KEYINPUT81), .Z(new_n229));
  INV_X1    g043(.A(G217), .ZN(new_n230));
  XOR2_X1   g044(.A(KEYINPUT76), .B(G902), .Z(new_n231));
  AOI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(G234), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(G902), .ZN(new_n233));
  INV_X1    g047(.A(new_n231), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n234), .B1(new_n226), .B2(new_n227), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT25), .ZN(new_n236));
  OR2_X1    g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  XOR2_X1   g051(.A(new_n232), .B(KEYINPUT78), .Z(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n239), .B1(new_n235), .B2(new_n236), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n229), .A2(new_n233), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G143), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT1), .B1(new_n243), .B2(G146), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT69), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n205), .A2(G143), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(KEYINPUT1), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n190), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(G143), .B(G146), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n251), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n243), .A2(G146), .ZN(new_n254));
  AND4_X1   g068(.A1(new_n251), .A2(new_n252), .A3(new_n246), .A4(new_n254), .ZN(new_n255));
  OAI22_X1  g069(.A1(new_n249), .A2(new_n250), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n257));
  INV_X1    g071(.A(G137), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G134), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT65), .B(G137), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n259), .B1(new_n260), .B2(G134), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT11), .B1(new_n258), .B2(G134), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n259), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n258), .A2(KEYINPUT65), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT65), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G137), .ZN(new_n266));
  AND2_X1   g080(.A1(KEYINPUT11), .A2(G134), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(G131), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n263), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT66), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n263), .A2(new_n268), .A3(KEYINPUT66), .A4(new_n269), .ZN(new_n273));
  AOI221_X4 g087(.A(new_n257), .B1(G131), .B2(new_n261), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n273), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n261), .A2(G131), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT67), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n256), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n263), .A2(new_n268), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G131), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n260), .A2(new_n267), .B1(new_n262), .B2(new_n259), .ZN(new_n281));
  AOI21_X1  g095(.A(KEYINPUT66), .B1(new_n281), .B2(new_n269), .ZN(new_n282));
  INV_X1    g096(.A(new_n273), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n280), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(KEYINPUT0), .B(G128), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n246), .A2(new_n254), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(KEYINPUT64), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT64), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n289), .B1(new_n250), .B2(new_n285), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n250), .A2(KEYINPUT0), .A3(G128), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n284), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(KEYINPUT30), .B1(new_n278), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n296));
  INV_X1    g110(.A(G116), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n297), .A2(G119), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n188), .A2(G116), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT70), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT2), .B(G113), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n188), .A2(G116), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n297), .A2(G119), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT70), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n302), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n300), .A2(new_n301), .A3(new_n305), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n306), .A2(KEYINPUT71), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT71), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n300), .A2(new_n308), .A3(new_n301), .A4(new_n305), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n302), .A2(new_n303), .ZN(new_n310));
  OR2_X1    g124(.A1(new_n310), .A2(new_n301), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n296), .B1(new_n307), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n306), .A2(KEYINPUT71), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n314), .A2(KEYINPUT72), .A3(new_n309), .A4(new_n311), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n275), .A2(new_n276), .A3(new_n256), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n294), .A2(KEYINPUT30), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n295), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(G237), .A2(G953), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G210), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n322), .B(KEYINPUT27), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT26), .B(G101), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n323), .B(new_n324), .ZN(new_n325));
  AOI22_X1  g139(.A1(new_n272), .A2(new_n273), .B1(G131), .B2(new_n279), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n317), .B1(new_n326), .B2(new_n292), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n313), .A2(new_n315), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n325), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT73), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n294), .A2(new_n313), .A3(new_n315), .A4(new_n317), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT73), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n332), .A3(new_n325), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT31), .B1(new_n320), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n325), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT28), .ZN(new_n337));
  INV_X1    g151(.A(new_n256), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n276), .B1(new_n282), .B2(new_n283), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n257), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n275), .A2(KEYINPUT67), .A3(new_n276), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n338), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n292), .B1(new_n275), .B2(new_n280), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n328), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n337), .B1(new_n344), .B2(new_n331), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT74), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n275), .A2(new_n276), .A3(new_n256), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n346), .B1(new_n347), .B2(new_n343), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n294), .A2(KEYINPUT74), .A3(new_n317), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT28), .B1(new_n350), .B2(new_n316), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n336), .B1(new_n345), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n340), .A2(new_n341), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n343), .B1(new_n353), .B2(new_n256), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n318), .B(new_n328), .C1(new_n354), .C2(KEYINPUT30), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT31), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n355), .A2(new_n356), .A3(new_n330), .A4(new_n333), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n335), .A2(new_n352), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(G472), .A2(G902), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT32), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n358), .A2(KEYINPUT32), .A3(new_n359), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(KEYINPUT75), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT32), .B1(new_n358), .B2(new_n359), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT75), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n327), .A2(new_n328), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n337), .B1(new_n369), .B2(new_n331), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n351), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n336), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n234), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n316), .B1(new_n278), .B2(new_n294), .ZN(new_n375));
  INV_X1    g189(.A(new_n331), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT28), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR3_X1   g191(.A1(new_n347), .A2(new_n343), .A3(new_n346), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT74), .B1(new_n294), .B2(new_n317), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n316), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n337), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n377), .A2(new_n381), .A3(new_n325), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n372), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n325), .B1(new_n355), .B2(new_n331), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n374), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n385), .A2(G472), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT77), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(KEYINPUT77), .A3(G472), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n242), .B1(new_n368), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(G214), .B1(G237), .B2(G902), .ZN(new_n392));
  XOR2_X1   g206(.A(new_n392), .B(KEYINPUT88), .Z(new_n393));
  AND3_X1   g207(.A1(new_n292), .A2(KEYINPUT89), .A3(G125), .ZN(new_n394));
  AOI21_X1  g208(.A(KEYINPUT89), .B1(new_n292), .B2(G125), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT90), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n397), .B1(new_n256), .B2(G125), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n245), .A2(new_n248), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n287), .B1(new_n399), .B2(new_n190), .ZN(new_n400));
  OR2_X1    g214(.A1(new_n253), .A2(new_n255), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT90), .A4(new_n201), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G953), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n404), .A2(G224), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT7), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n396), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(G110), .B(G122), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(KEYINPUT8), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT91), .ZN(new_n411));
  INV_X1    g225(.A(G104), .ZN(new_n412));
  OAI21_X1  g226(.A(KEYINPUT3), .B1(new_n412), .B2(G107), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT3), .ZN(new_n414));
  INV_X1    g228(.A(G107), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n415), .A3(G104), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(G107), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n413), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(KEYINPUT84), .B(G101), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT85), .B1(new_n412), .B2(G107), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT85), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(new_n415), .A3(G104), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n423), .A3(new_n417), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G101), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n420), .A2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G113), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT5), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n427), .B1(new_n298), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n429), .B1(new_n428), .B2(new_n310), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n311), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n411), .B1(new_n426), .B2(new_n431), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n418), .A2(new_n419), .B1(new_n424), .B2(G101), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n433), .A2(KEYINPUT91), .A3(new_n311), .A4(new_n430), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n300), .A2(new_n305), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n429), .B1(new_n436), .B2(new_n428), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n433), .B1(new_n437), .B2(new_n311), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n410), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n408), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n413), .A2(new_n416), .A3(new_n417), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(G101), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n420), .A2(new_n442), .A3(KEYINPUT4), .ZN(new_n443));
  OR2_X1    g257(.A1(new_n442), .A2(KEYINPUT4), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n445), .B1(new_n313), .B2(new_n315), .ZN(new_n446));
  INV_X1    g260(.A(new_n409), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n437), .A2(new_n311), .A3(new_n433), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NOR3_X1   g263(.A1(new_n446), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n440), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n292), .A2(G125), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n407), .B1(new_n403), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT92), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n398), .A2(new_n402), .B1(G125), .B2(new_n292), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT92), .B1(new_n456), .B2(new_n407), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(G902), .B1(new_n451), .B2(new_n458), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n409), .B(new_n448), .C1(new_n316), .C2(new_n445), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n447), .B1(new_n446), .B2(new_n449), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(KEYINPUT6), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n463), .B(new_n447), .C1(new_n446), .C2(new_n449), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n396), .A2(new_n403), .A3(new_n405), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n405), .B1(new_n396), .B2(new_n403), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n462), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n459), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g283(.A(G210), .B1(G237), .B2(G902), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(KEYINPUT93), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n471), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n459), .A2(new_n468), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n393), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT9), .B(G234), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G902), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n219), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n253), .A2(new_n255), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n250), .B1(G128), .B2(new_n244), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n433), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n256), .B2(new_n433), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n326), .A2(KEYINPUT86), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT12), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n485), .B1(new_n483), .B2(new_n484), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT87), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n488), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT87), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n486), .ZN(new_n492));
  XNOR2_X1  g306(.A(G110), .B(G140), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(KEYINPUT82), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT83), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G227), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n496), .B1(new_n497), .B2(G953), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n494), .B(KEYINPUT83), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(G227), .A3(new_n404), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT10), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n482), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n293), .A2(new_n443), .A3(new_n444), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n256), .A2(KEYINPUT10), .A3(new_n433), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n503), .A2(new_n504), .A3(new_n326), .A4(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n501), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n489), .A2(new_n492), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n284), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n506), .ZN(new_n512));
  INV_X1    g326(.A(new_n501), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G469), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n516), .A3(new_n231), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n490), .A2(new_n506), .A3(new_n486), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n513), .A2(new_n518), .B1(new_n508), .B2(new_n511), .ZN(new_n519));
  OAI21_X1  g333(.A(G469), .B1(new_n519), .B2(G902), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n479), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT20), .ZN(new_n522));
  INV_X1    g336(.A(G237), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n523), .A2(new_n404), .A3(G143), .A4(G214), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT94), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT94), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n321), .A2(new_n526), .A3(G143), .A4(G214), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(G143), .B1(new_n321), .B2(G214), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n269), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT17), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n529), .B1(new_n525), .B2(new_n527), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n269), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n528), .A2(new_n530), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(KEYINPUT17), .A3(G131), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT96), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n210), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n531), .A2(KEYINPUT96), .A3(KEYINPUT17), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n536), .A2(new_n540), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  XOR2_X1   g357(.A(G113), .B(G122), .Z(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT95), .B(G104), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n537), .A2(KEYINPUT18), .A3(G131), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT18), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n534), .B1(new_n548), .B2(new_n269), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n203), .A2(G146), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n206), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n547), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n543), .A2(new_n546), .A3(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n203), .B(KEYINPUT19), .ZN(new_n554));
  AOI211_X1 g368(.A(G131), .B(new_n529), .C1(new_n525), .C2(new_n527), .ZN(new_n555));
  OAI221_X1 g369(.A(new_n204), .B1(new_n554), .B2(G146), .C1(new_n531), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n552), .ZN(new_n557));
  INV_X1    g371(.A(new_n546), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n553), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(G475), .A2(G902), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n522), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n561), .ZN(new_n563));
  AOI211_X1 g377(.A(KEYINPUT20), .B(new_n563), .C1(new_n553), .C2(new_n559), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n543), .A2(new_n552), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n558), .ZN(new_n566));
  AOI21_X1  g380(.A(G902), .B1(new_n566), .B2(new_n553), .ZN(new_n567));
  INV_X1    g381(.A(G475), .ZN(new_n568));
  OAI22_X1  g382(.A1(new_n562), .A2(new_n564), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G952), .ZN(new_n571));
  AOI211_X1 g385(.A(G953), .B(new_n571), .C1(G234), .C2(G237), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n234), .B(G953), .C1(new_n220), .C2(new_n523), .ZN(new_n574));
  XOR2_X1   g388(.A(KEYINPUT21), .B(G898), .Z(new_n575));
  OAI21_X1  g389(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n190), .A2(G143), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n243), .A2(G128), .ZN(new_n578));
  OAI21_X1  g392(.A(G134), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n243), .A2(G128), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n190), .A2(G143), .ZN(new_n581));
  INV_X1    g395(.A(G134), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(G122), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(G116), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n297), .A2(G122), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(new_n587), .A3(new_n415), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n586), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n587), .B1(new_n590), .B2(KEYINPUT14), .ZN(new_n591));
  OR2_X1    g405(.A1(new_n587), .A2(KEYINPUT14), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n415), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n588), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n415), .B1(new_n586), .B2(new_n587), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n583), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT13), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n580), .B1(new_n578), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n577), .A2(KEYINPUT13), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n582), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI22_X1  g414(.A1(new_n589), .A2(new_n593), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n476), .A2(new_n230), .A3(G953), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  OAI221_X1 g418(.A(new_n602), .B1(new_n596), .B2(new_n600), .C1(new_n589), .C2(new_n593), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(KEYINPUT97), .B1(new_n606), .B2(new_n231), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT97), .ZN(new_n608));
  AOI211_X1 g422(.A(new_n608), .B(new_n234), .C1(new_n604), .C2(new_n605), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(G478), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT98), .ZN(new_n613));
  OR2_X1    g427(.A1(new_n613), .A2(KEYINPUT15), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(KEYINPUT15), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n612), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n606), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n234), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n617), .B1(new_n619), .B2(new_n616), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n570), .A2(new_n576), .A3(new_n620), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n475), .A2(new_n521), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n391), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(new_n623), .B(new_n419), .Z(G3));
  INV_X1    g438(.A(new_n474), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n473), .B1(new_n459), .B2(new_n468), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n392), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n472), .A2(new_n474), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(KEYINPUT99), .A3(new_n392), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n231), .A2(G478), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n606), .A2(KEYINPUT33), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n604), .A2(new_n605), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n632), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n636), .B1(new_n610), .B2(new_n612), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n546), .B1(new_n556), .B2(new_n552), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n547), .A2(new_n549), .A3(new_n551), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n531), .A2(new_n555), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n210), .B1(new_n640), .B2(new_n533), .ZN(new_n641));
  AOI21_X1  g455(.A(KEYINPUT96), .B1(new_n531), .B2(KEYINPUT17), .ZN(new_n642));
  NOR4_X1   g456(.A1(new_n534), .A2(new_n539), .A3(new_n533), .A4(new_n269), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n639), .B1(new_n641), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n638), .B1(new_n645), .B2(new_n546), .ZN(new_n646));
  OAI21_X1  g460(.A(KEYINPUT20), .B1(new_n646), .B2(new_n563), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n560), .A2(new_n522), .A3(new_n561), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n553), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n546), .B1(new_n543), .B2(new_n552), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n478), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(G475), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n637), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  AND4_X1   g468(.A1(new_n576), .A2(new_n629), .A3(new_n631), .A4(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n358), .A2(new_n231), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(G472), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n658), .A2(new_n241), .A3(new_n360), .A4(new_n521), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT34), .B(G104), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G6));
  NOR2_X1   g476(.A1(new_n620), .A2(new_n569), .ZN(new_n663));
  AND4_X1   g477(.A1(new_n576), .A2(new_n629), .A3(new_n631), .A4(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n659), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT35), .B(G107), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  NAND2_X1  g482(.A1(new_n237), .A2(new_n240), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n223), .A2(KEYINPUT36), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n216), .B(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n233), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n475), .A2(new_n621), .A3(new_n521), .A4(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n658), .A2(new_n360), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT37), .B(G110), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G12));
  AND3_X1   g492(.A1(new_n358), .A2(KEYINPUT32), .A3(new_n359), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n679), .A2(new_n365), .A3(new_n366), .ZN(new_n680));
  INV_X1    g494(.A(new_n367), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n390), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n573), .B1(new_n574), .B2(G900), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT100), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n620), .A2(new_n569), .A3(new_n684), .ZN(new_n685));
  AND4_X1   g499(.A1(new_n629), .A2(new_n631), .A3(new_n673), .A4(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n682), .A2(new_n521), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G128), .ZN(G30));
  XNOR2_X1  g502(.A(new_n630), .B(KEYINPUT38), .ZN(new_n689));
  INV_X1    g503(.A(new_n673), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n570), .A2(new_n620), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n689), .A2(new_n392), .A3(new_n690), .A4(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n684), .B(KEYINPUT39), .Z(new_n693));
  NAND2_X1  g507(.A1(new_n521), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n694), .B(KEYINPUT101), .Z(new_n695));
  AOI21_X1  g509(.A(new_n692), .B1(new_n695), .B2(KEYINPUT40), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n320), .A2(new_n334), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n325), .B1(new_n369), .B2(new_n331), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n478), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(G472), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n700), .B1(new_n680), .B2(new_n681), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n696), .B(new_n701), .C1(KEYINPUT40), .C2(new_n695), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G143), .ZN(G45));
  INV_X1    g517(.A(new_n684), .ZN(new_n704));
  AOI21_X1  g518(.A(KEYINPUT102), .B1(new_n654), .B2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n637), .ZN(new_n706));
  AND4_X1   g520(.A1(KEYINPUT102), .A2(new_n569), .A3(new_n706), .A4(new_n704), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  AND4_X1   g522(.A1(new_n629), .A2(new_n708), .A3(new_n631), .A4(new_n673), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n682), .A2(new_n521), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G146), .ZN(G48));
  NAND2_X1  g525(.A1(new_n490), .A2(new_n486), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n507), .B1(new_n712), .B2(KEYINPUT87), .ZN(new_n713));
  AOI22_X1  g527(.A1(new_n713), .A2(new_n492), .B1(new_n512), .B2(new_n513), .ZN(new_n714));
  OAI21_X1  g528(.A(G469), .B1(new_n714), .B2(new_n234), .ZN(new_n715));
  INV_X1    g529(.A(new_n479), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n715), .A2(new_n716), .A3(new_n517), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT103), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n715), .A2(new_n517), .A3(KEYINPUT103), .A4(new_n716), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n682), .A2(new_n655), .A3(new_n241), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NAND4_X1  g538(.A1(new_n682), .A2(new_n664), .A3(new_n241), .A4(new_n721), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  AND4_X1   g540(.A1(new_n576), .A2(new_n673), .A3(new_n570), .A4(new_n620), .ZN(new_n727));
  INV_X1    g541(.A(new_n717), .ZN(new_n728));
  AND4_X1   g542(.A1(new_n629), .A2(new_n727), .A3(new_n728), .A4(new_n631), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n682), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  NAND3_X1  g545(.A1(new_n719), .A2(new_n576), .A3(new_n720), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n629), .A2(new_n631), .A3(new_n691), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g548(.A(G472), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n358), .B2(new_n231), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n336), .B1(new_n351), .B2(new_n370), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n357), .A2(new_n737), .ZN(new_n738));
  AND2_X1   g552(.A1(new_n330), .A2(new_n333), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n356), .B1(new_n739), .B2(new_n355), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n359), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(KEYINPUT104), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n335), .A2(new_n357), .A3(new_n737), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT104), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(new_n744), .A3(new_n359), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n736), .B1(new_n742), .B2(new_n745), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n746), .A2(new_n241), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n734), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G122), .ZN(G24));
  OAI21_X1  g563(.A(KEYINPUT105), .B1(new_n705), .B2(new_n707), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT102), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n569), .A2(new_n706), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n751), .B1(new_n752), .B2(new_n684), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT105), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n654), .A2(KEYINPUT102), .A3(new_n704), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n750), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(new_n745), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n744), .B1(new_n743), .B2(new_n359), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n658), .B(new_n673), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n629), .A2(new_n631), .A3(new_n728), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G125), .ZN(G27));
  INV_X1    g578(.A(KEYINPUT106), .ZN(new_n765));
  AOI22_X1  g579(.A1(new_n364), .A2(new_n367), .B1(new_n388), .B2(new_n389), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n750), .A2(new_n756), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n392), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n630), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n521), .ZN(new_n771));
  NOR4_X1   g585(.A1(new_n766), .A2(new_n768), .A3(new_n242), .A4(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n679), .A2(new_n365), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n242), .B1(new_n390), .B2(new_n773), .ZN(new_n774));
  AOI211_X1 g588(.A(G469), .B(new_n234), .C1(new_n509), .C2(new_n514), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n518), .A2(new_n513), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n508), .A2(new_n511), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n516), .B1(new_n778), .B2(new_n478), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n716), .B1(new_n775), .B2(new_n779), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n780), .A2(new_n630), .A3(new_n769), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n781), .A2(new_n750), .A3(new_n756), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n767), .B1(new_n774), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n765), .B1(new_n772), .B2(new_n783), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n385), .A2(KEYINPUT77), .A3(G472), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT77), .B1(new_n385), .B2(G472), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n362), .A2(new_n363), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n241), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n781), .A2(new_n750), .A3(new_n756), .ZN(new_n790));
  OAI21_X1  g604(.A(KEYINPUT42), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n768), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n682), .A2(new_n792), .A3(new_n241), .A4(new_n781), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n791), .A2(new_n793), .A3(KEYINPUT106), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n784), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(new_n269), .ZN(G33));
  NAND4_X1  g610(.A1(new_n682), .A2(new_n241), .A3(new_n685), .A4(new_n781), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G134), .ZN(G36));
  NAND2_X1  g612(.A1(new_n570), .A2(new_n706), .ZN(new_n799));
  XOR2_X1   g613(.A(new_n799), .B(KEYINPUT43), .Z(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n675), .A3(new_n673), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT44), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT107), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(new_n804), .A3(new_n770), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n778), .B(KEYINPUT45), .ZN(new_n806));
  OAI21_X1  g620(.A(G469), .B1(new_n806), .B2(G902), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n775), .B1(new_n807), .B2(KEYINPUT46), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n808), .B1(KEYINPUT46), .B2(new_n807), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n809), .A2(new_n716), .A3(new_n693), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n801), .A2(new_n802), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n805), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n804), .B1(new_n803), .B2(new_n770), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G137), .ZN(G39));
  NAND2_X1  g629(.A1(new_n809), .A2(new_n716), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT47), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n766), .A2(new_n242), .A3(new_n708), .A4(new_n770), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT108), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n819), .A2(KEYINPUT108), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n818), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT109), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n818), .A2(KEYINPUT109), .A3(new_n820), .A4(new_n821), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(new_n198), .ZN(G42));
  NAND3_X1  g641(.A1(new_n747), .A2(new_n572), .A3(new_n800), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n715), .A2(new_n517), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n830), .A2(new_n479), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n770), .B(new_n829), .C1(new_n818), .C2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT50), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n392), .B1(KEYINPUT115), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n728), .A2(new_n834), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n828), .A2(new_n689), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n833), .A2(KEYINPUT115), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n836), .B(new_n837), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n717), .A2(new_n630), .A3(new_n769), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n800), .A2(new_n572), .A3(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n832), .B(new_n838), .C1(new_n760), .C2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n839), .A2(new_n241), .A3(new_n572), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n701), .A2(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT116), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n844), .A2(new_n569), .A3(new_n706), .ZN(new_n845));
  OAI21_X1  g659(.A(KEYINPUT114), .B1(new_n841), .B2(new_n845), .ZN(new_n846));
  OR2_X1    g660(.A1(new_n846), .A2(KEYINPUT51), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(KEYINPUT51), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n844), .A2(new_n752), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n789), .A2(new_n840), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n850), .B(KEYINPUT48), .ZN(new_n851));
  INV_X1    g665(.A(new_n762), .ZN(new_n852));
  OAI211_X1 g666(.A(G952), .B(new_n404), .C1(new_n828), .C2(new_n852), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n849), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n847), .A2(new_n848), .A3(new_n854), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n766), .A2(new_n242), .A3(new_n771), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n746), .A2(new_n673), .A3(new_n750), .A4(new_n756), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n673), .A2(new_n570), .A3(new_n620), .A4(new_n704), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n857), .B1(new_n766), .B2(new_n858), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n685), .A2(new_n856), .B1(new_n859), .B2(new_n781), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n784), .A2(new_n860), .A3(new_n794), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n752), .B1(new_n620), .B2(new_n569), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n475), .A2(new_n576), .A3(new_n862), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n659), .A2(new_n863), .B1(new_n674), .B2(new_n675), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n864), .B1(new_n391), .B2(new_n622), .ZN(new_n865));
  AOI22_X1  g679(.A1(new_n734), .A2(new_n747), .B1(new_n682), .B2(new_n729), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n865), .A2(new_n866), .A3(new_n722), .A4(new_n725), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n861), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n869));
  INV_X1    g683(.A(new_n733), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n228), .A2(new_n236), .A3(new_n231), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n238), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n235), .A2(new_n236), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n672), .B(new_n704), .C1(new_n872), .C2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(KEYINPUT110), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT110), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n669), .A2(new_n876), .A3(new_n672), .A4(new_n704), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n521), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT111), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT111), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n521), .A2(new_n875), .A3(new_n880), .A4(new_n877), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n701), .A2(new_n870), .A3(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n687), .A2(new_n710), .A3(new_n883), .A4(new_n763), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT52), .ZN(new_n885));
  OR3_X1    g699(.A1(new_n884), .A2(KEYINPUT112), .A3(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n884), .A2(new_n885), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n780), .B1(new_n368), .B2(new_n390), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n888), .A2(new_n686), .B1(new_n761), .B2(new_n762), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n889), .A2(KEYINPUT52), .A3(new_n710), .A4(new_n883), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n887), .A2(KEYINPUT112), .A3(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n868), .A2(new_n869), .A3(new_n886), .A4(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n867), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n893), .A2(new_n784), .A3(new_n794), .A4(new_n860), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n887), .A2(new_n890), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n892), .B(KEYINPUT54), .C1(new_n897), .C2(new_n869), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n869), .B1(new_n894), .B2(new_n896), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT54), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n865), .A2(KEYINPUT53), .A3(new_n791), .A4(new_n793), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n722), .A2(new_n725), .A3(new_n730), .A4(new_n748), .ZN(new_n902));
  INV_X1    g716(.A(new_n858), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n750), .A2(new_n756), .ZN(new_n904));
  INV_X1    g718(.A(new_n760), .ZN(new_n905));
  AOI22_X1  g719(.A1(new_n682), .A2(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n797), .B1(new_n906), .B2(new_n771), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n901), .A2(new_n902), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n891), .A3(new_n886), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n899), .A2(new_n900), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT113), .B1(new_n898), .B2(new_n910), .ZN(new_n911));
  AND3_X1   g725(.A1(new_n898), .A2(KEYINPUT113), .A3(new_n910), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n855), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(G952), .A2(G953), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n830), .B(KEYINPUT49), .Z(new_n915));
  OR3_X1    g729(.A1(new_n242), .A2(new_n393), .A3(new_n479), .ZN(new_n916));
  OR4_X1    g730(.A1(new_n689), .A2(new_n915), .A3(new_n799), .A4(new_n916), .ZN(new_n917));
  OAI22_X1  g731(.A1(new_n913), .A2(new_n914), .B1(new_n701), .B2(new_n917), .ZN(G75));
  AOI21_X1  g732(.A(KEYINPUT53), .B1(new_n868), .B2(new_n895), .ZN(new_n919));
  AND3_X1   g733(.A1(new_n908), .A2(new_n891), .A3(new_n886), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n234), .B(new_n471), .C1(new_n919), .C2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT56), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n462), .A2(new_n464), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(new_n467), .Z(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT55), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT117), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT117), .ZN(new_n928));
  INV_X1    g742(.A(new_n926), .ZN(new_n929));
  AOI211_X1 g743(.A(new_n928), .B(new_n929), .C1(new_n921), .C2(new_n922), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n404), .A2(G952), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT118), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n921), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n926), .B(KEYINPUT119), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n922), .B(new_n937), .C1(new_n921), .C2(new_n934), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n933), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT120), .B1(new_n931), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n231), .B1(new_n899), .B2(new_n909), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT56), .B1(new_n941), .B2(new_n471), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n928), .B1(new_n942), .B2(new_n929), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n923), .A2(KEYINPUT117), .A3(new_n926), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n937), .A2(new_n922), .ZN(new_n946));
  INV_X1    g760(.A(new_n921), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(KEYINPUT118), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n932), .B1(new_n948), .B2(new_n935), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT120), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n945), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n940), .A2(new_n951), .ZN(G51));
  NAND2_X1  g766(.A1(G469), .A2(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT57), .ZN(new_n954));
  OAI21_X1  g768(.A(KEYINPUT54), .B1(new_n919), .B2(new_n920), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n954), .B1(new_n955), .B2(new_n910), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n956), .A2(new_n714), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n957), .A2(KEYINPUT121), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n941), .A2(G469), .A3(new_n806), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n959), .B1(new_n957), .B2(KEYINPUT121), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n932), .B1(new_n958), .B2(new_n960), .ZN(G54));
  AND3_X1   g775(.A1(new_n941), .A2(KEYINPUT58), .A3(G475), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n933), .B1(new_n962), .B2(new_n560), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(new_n560), .B2(new_n962), .ZN(G60));
  NAND2_X1  g778(.A1(new_n955), .A2(new_n910), .ZN(new_n965));
  NAND2_X1  g779(.A1(G478), .A2(G902), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT59), .ZN(new_n967));
  INV_X1    g781(.A(new_n633), .ZN(new_n968));
  INV_X1    g782(.A(new_n635), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n965), .B(new_n967), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n933), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n968), .A2(new_n969), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n967), .B1(new_n912), .B2(new_n911), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(G63));
  INV_X1    g788(.A(KEYINPUT61), .ZN(new_n975));
  NAND2_X1  g789(.A1(G217), .A2(G902), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT60), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n899), .B2(new_n909), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n932), .B1(new_n978), .B2(new_n671), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n975), .B1(new_n979), .B2(KEYINPUT122), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n979), .B1(new_n229), .B2(new_n978), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n980), .B(new_n981), .Z(G66));
  NAND3_X1  g796(.A1(new_n575), .A2(G224), .A3(G953), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n983), .B1(new_n867), .B2(G953), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT123), .Z(new_n985));
  OAI21_X1  g799(.A(new_n924), .B1(G898), .B2(new_n404), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(G69));
  NAND2_X1  g801(.A1(new_n889), .A2(new_n710), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT124), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n988), .B(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n814), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT126), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n810), .A2(new_n870), .A3(new_n774), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n797), .ZN(new_n994));
  NOR3_X1   g808(.A1(new_n826), .A2(new_n795), .A3(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n992), .A2(new_n404), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n318), .B1(new_n354), .B2(KEYINPUT30), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(new_n554), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n999), .B1(G900), .B2(G953), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT125), .ZN(new_n1002));
  INV_X1    g816(.A(new_n694), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n391), .A2(new_n1003), .A3(new_n770), .A4(new_n862), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1004), .B1(new_n812), .B2(new_n813), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1005), .B1(new_n824), .B2(new_n825), .ZN(new_n1006));
  AND3_X1   g820(.A1(new_n990), .A2(KEYINPUT62), .A3(new_n702), .ZN(new_n1007));
  AOI21_X1  g821(.A(KEYINPUT62), .B1(new_n990), .B2(new_n702), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n404), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1002), .B1(new_n1010), .B2(new_n999), .ZN(new_n1011));
  AOI211_X1 g825(.A(KEYINPUT125), .B(new_n998), .C1(new_n1009), .C2(new_n404), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1001), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n404), .B1(G227), .B2(G900), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1014), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n1001), .B(new_n1016), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1015), .A2(new_n1017), .ZN(G72));
  NOR2_X1   g832(.A1(new_n320), .A2(new_n376), .ZN(new_n1019));
  OR2_X1    g833(.A1(new_n1009), .A2(new_n867), .ZN(new_n1020));
  NAND2_X1  g834(.A1(G472), .A2(G902), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1021), .B(KEYINPUT63), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1022), .B(KEYINPUT127), .ZN(new_n1023));
  AOI211_X1 g837(.A(new_n336), .B(new_n1019), .C1(new_n1020), .C2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1019), .A2(new_n336), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n992), .A2(new_n893), .A3(new_n995), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1025), .B1(new_n1026), .B2(new_n1023), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n892), .B1(new_n897), .B2(new_n869), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n697), .A2(new_n384), .ZN(new_n1029));
  NOR3_X1   g843(.A1(new_n1028), .A2(new_n1022), .A3(new_n1029), .ZN(new_n1030));
  NOR4_X1   g844(.A1(new_n1024), .A2(new_n1027), .A3(new_n932), .A4(new_n1030), .ZN(G57));
endmodule


