//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 0 0 0 1 0 0 1 1 0 0 0 0 0 1 0 0 1 1 1 1 0 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1073, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NAND2_X1  g0005(.A1(G87), .A2(G250), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G50), .A2(G226), .ZN(new_n208));
  INV_X1    g0008(.A(G116), .ZN(new_n209));
  INV_X1    g0009(.A(G270), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n207), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n206), .B1(new_n211), .B2(KEYINPUT64), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(KEYINPUT64), .B2(new_n211), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G97), .A2(G257), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G58), .A2(G232), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G107), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n205), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(KEYINPUT65), .B2(KEYINPUT1), .ZN(new_n221));
  NOR2_X1   g0021(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n221), .B(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G68), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G50), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  NOR3_X1   g0029(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n205), .A2(G13), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n231), .B(G250), .C1(G257), .C2(G264), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT0), .Z(new_n233));
  NOR3_X1   g0033(.A1(new_n223), .A2(new_n230), .A3(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G264), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n210), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n238), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G13), .A3(G20), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G68), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT12), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(KEYINPUT71), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n256), .B1(new_n254), .B2(new_n253), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n229), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n228), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G50), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n261), .A2(G20), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n265), .A2(G77), .B1(G20), .B2(new_n225), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n260), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT70), .B(KEYINPUT11), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n267), .B(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n259), .B1(new_n251), .B2(G20), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n257), .B(new_n269), .C1(new_n225), .C2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G41), .A2(G45), .ZN(new_n273));
  INV_X1    g0073(.A(G274), .ZN(new_n274));
  NOR3_X1   g0074(.A1(new_n273), .A2(G1), .A3(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G226), .A2(G1698), .ZN(new_n276));
  INV_X1    g0076(.A(G232), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n276), .B1(new_n277), .B2(G1698), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G97), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n229), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G33), .A2(G41), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n275), .B1(new_n282), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT13), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT67), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n289), .B1(new_n273), .B2(G1), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n251), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n290), .A2(new_n291), .B1(new_n283), .B2(new_n284), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G238), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n287), .A2(new_n288), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n275), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n278), .A2(new_n279), .B1(G33), .B2(G97), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n295), .B1(new_n296), .B2(new_n285), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n292), .A2(G238), .ZN(new_n298));
  OAI21_X1  g0098(.A(KEYINPUT13), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G169), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT72), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT73), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n300), .A2(KEYINPUT72), .A3(new_n304), .A4(G169), .ZN(new_n305));
  AND3_X1   g0105(.A1(new_n303), .A2(KEYINPUT14), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n300), .A2(new_n304), .A3(G169), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  OAI22_X1  g0108(.A1(new_n307), .A2(KEYINPUT14), .B1(new_n308), .B2(new_n300), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n272), .B1(new_n306), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n272), .B1(G200), .B2(new_n300), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n294), .A2(new_n299), .A3(G190), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(KEYINPUT69), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n312), .A2(KEYINPUT69), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n311), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G1698), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(G222), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G223), .A2(G1698), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n279), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n320), .B(new_n286), .C1(G77), .C2(new_n279), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n295), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n322), .B1(G226), .B2(new_n292), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G190), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT9), .ZN(new_n325));
  OAI21_X1  g0125(.A(G20), .B1(new_n226), .B2(G50), .ZN(new_n326));
  INV_X1    g0126(.A(G150), .ZN(new_n327));
  INV_X1    g0127(.A(new_n265), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT8), .B(G58), .ZN(new_n329));
  OAI221_X1 g0129(.A(new_n326), .B1(new_n327), .B2(new_n262), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n330), .A2(new_n259), .B1(G50), .B2(new_n270), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(G50), .B2(new_n252), .ZN(new_n332));
  INV_X1    g0132(.A(G200), .ZN(new_n333));
  OAI221_X1 g0133(.A(new_n324), .B1(new_n325), .B2(new_n332), .C1(new_n333), .C2(new_n323), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(new_n325), .B2(new_n332), .ZN(new_n335));
  XOR2_X1   g0135(.A(new_n335), .B(KEYINPUT10), .Z(new_n336));
  NAND2_X1  g0136(.A1(new_n323), .A2(new_n308), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n337), .B(new_n332), .C1(G169), .C2(new_n323), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(G238), .A2(G1698), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n279), .B(new_n340), .C1(new_n277), .C2(G1698), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(new_n286), .C1(G107), .C2(new_n279), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n292), .A2(G244), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(new_n295), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G200), .ZN(new_n345));
  INV_X1    g0145(.A(new_n329), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n346), .A2(new_n263), .B1(G20), .B2(G77), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT15), .B(G87), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n347), .B1(new_n328), .B2(new_n348), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n349), .A2(new_n259), .B1(G77), .B2(new_n270), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(G77), .B2(new_n252), .ZN(new_n351));
  INV_X1    g0151(.A(G190), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT68), .B1(new_n344), .B2(new_n352), .ZN(new_n353));
  OR3_X1    g0153(.A1(new_n344), .A2(KEYINPUT68), .A3(new_n352), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n351), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI211_X1 g0155(.A(new_n316), .B(new_n339), .C1(new_n345), .C2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT77), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT75), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT74), .ZN(new_n359));
  AOI211_X1 g0159(.A(new_n359), .B(new_n275), .C1(new_n292), .C2(G232), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n290), .A2(new_n291), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(G232), .A3(new_n285), .ZN(new_n362));
  AOI21_X1  g0162(.A(KEYINPUT74), .B1(new_n362), .B2(new_n295), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n358), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  AOI221_X4 g0164(.A(new_n277), .B1(new_n283), .B2(new_n284), .C1(new_n290), .C2(new_n291), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n359), .B1(new_n365), .B2(new_n275), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n362), .A2(KEYINPUT74), .A3(new_n295), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(KEYINPUT75), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n279), .B1(G226), .B2(new_n317), .ZN(new_n370));
  NOR2_X1   g0170(.A1(G223), .A2(G1698), .ZN(new_n371));
  INV_X1    g0171(.A(G87), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n370), .A2(new_n371), .B1(new_n261), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n286), .ZN(new_n374));
  XNOR2_X1  g0174(.A(KEYINPUT76), .B(G190), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n366), .A2(new_n374), .A3(new_n367), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n369), .A2(new_n378), .B1(new_n333), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT16), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G58), .A2(G68), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n228), .B1(new_n226), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT7), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n279), .B2(G20), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT3), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G33), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n389), .A2(KEYINPUT7), .A3(new_n228), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n383), .B1(new_n391), .B2(G68), .ZN(new_n392));
  INV_X1    g0192(.A(G159), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n262), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n381), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n225), .B1(new_n385), .B2(new_n390), .ZN(new_n397));
  NOR4_X1   g0197(.A1(new_n397), .A2(KEYINPUT16), .A3(new_n394), .A4(new_n383), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n259), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n252), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n329), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n271), .B2(new_n329), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n357), .B1(new_n380), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT7), .B1(new_n389), .B2(new_n228), .ZN(new_n406));
  AOI211_X1 g0206(.A(new_n384), .B(G20), .C1(new_n386), .C2(new_n388), .ZN(new_n407));
  OAI21_X1  g0207(.A(G68), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n383), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n395), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT16), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n392), .A2(new_n381), .A3(new_n395), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n402), .B1(new_n413), .B2(new_n259), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n377), .B1(new_n364), .B2(new_n368), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n360), .A2(new_n363), .ZN(new_n416));
  AOI21_X1  g0216(.A(G200), .B1(new_n416), .B2(new_n374), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n414), .B(KEYINPUT77), .C1(new_n415), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n405), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT17), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n399), .B(new_n403), .C1(new_n415), .C2(new_n417), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n421), .A2(KEYINPUT17), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n369), .A2(new_n308), .A3(new_n374), .ZN(new_n425));
  INV_X1    g0225(.A(G169), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n379), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n404), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  XNOR2_X1  g0228(.A(new_n428), .B(KEYINPUT18), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n344), .A2(new_n426), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n344), .A2(G179), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n351), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n424), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n356), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  XNOR2_X1  g0238(.A(KEYINPUT85), .B(KEYINPUT24), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n279), .A2(new_n228), .A3(G87), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT83), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n279), .A2(KEYINPUT83), .A3(new_n228), .A4(G87), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n442), .A2(KEYINPUT22), .A3(new_n443), .ZN(new_n444));
  OR2_X1    g0244(.A1(new_n440), .A2(KEYINPUT22), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(KEYINPUT84), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT84), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n442), .A2(new_n448), .A3(KEYINPUT22), .A4(new_n443), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n228), .A2(G107), .ZN(new_n450));
  XNOR2_X1  g0250(.A(new_n450), .B(KEYINPUT23), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n228), .A2(G33), .A3(G116), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n439), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n449), .A2(new_n452), .ZN(new_n455));
  INV_X1    g0255(.A(new_n439), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n455), .A2(new_n456), .A3(new_n446), .A4(new_n451), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n454), .A2(new_n457), .A3(new_n259), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT25), .ZN(new_n459));
  NOR3_X1   g0259(.A1(new_n252), .A2(new_n459), .A3(G107), .ZN(new_n460));
  XNOR2_X1  g0260(.A(new_n460), .B(KEYINPUT86), .ZN(new_n461));
  XOR2_X1   g0261(.A(new_n461), .B(KEYINPUT87), .Z(new_n462));
  OAI21_X1  g0262(.A(new_n459), .B1(new_n252), .B2(G107), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n251), .A2(G33), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n400), .B1(KEYINPUT79), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n464), .A2(KEYINPUT79), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(new_n259), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n462), .A2(new_n463), .B1(G107), .B2(new_n469), .ZN(new_n470));
  OR2_X1    g0270(.A1(G250), .A2(G1698), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n279), .B(new_n471), .C1(G257), .C2(new_n317), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G33), .A2(G294), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(new_n286), .ZN(new_n475));
  INV_X1    g0275(.A(G45), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(G1), .ZN(new_n477));
  AND2_X1   g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  NOR2_X1   g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OR2_X1    g0280(.A1(new_n480), .A2(new_n274), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n480), .A2(new_n285), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT88), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n483), .A3(G264), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n480), .A2(new_n285), .ZN(new_n485));
  OAI21_X1  g0285(.A(KEYINPUT88), .B1(new_n485), .B2(new_n218), .ZN(new_n486));
  AND4_X1   g0286(.A1(new_n475), .A2(new_n481), .A3(new_n484), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G190), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n475), .A2(new_n481), .A3(new_n484), .A4(new_n486), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G200), .ZN(new_n490));
  AND4_X1   g0290(.A1(new_n458), .A2(new_n470), .A3(new_n488), .A4(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT89), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n489), .A2(new_n492), .A3(G169), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n492), .B1(new_n489), .B2(G169), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n487), .A2(G179), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n458), .A2(new_n470), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(G257), .A2(G1698), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n317), .A2(G264), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n279), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n501), .B1(G303), .B2(new_n279), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT82), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n501), .B(KEYINPUT82), .C1(G303), .C2(new_n279), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(new_n286), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n480), .A2(G270), .A3(new_n285), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT81), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n507), .B(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n506), .A2(new_n509), .A3(new_n481), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n400), .A2(new_n209), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G283), .ZN(new_n512));
  INV_X1    g0312(.A(G97), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n512), .B(new_n228), .C1(G33), .C2(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n514), .B(new_n259), .C1(new_n228), .C2(G116), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT20), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n515), .A2(new_n516), .ZN(new_n518));
  OAI221_X1 g0318(.A(new_n511), .B1(new_n468), .B2(new_n209), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n510), .A2(G169), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT21), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OR2_X1    g0322(.A1(new_n520), .A2(new_n521), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n506), .A2(new_n509), .A3(G179), .A4(new_n481), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n519), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n510), .A2(G200), .ZN(new_n527));
  INV_X1    g0327(.A(new_n519), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n527), .B(new_n528), .C1(new_n376), .C2(new_n510), .ZN(new_n529));
  AND4_X1   g0329(.A1(new_n522), .A2(new_n523), .A3(new_n526), .A4(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT4), .ZN(new_n531));
  INV_X1    g0331(.A(G244), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n531), .B1(new_n389), .B2(new_n532), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n279), .A2(KEYINPUT4), .A3(G244), .A4(new_n317), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n533), .A2(new_n534), .A3(new_n512), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n279), .A2(G250), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n317), .B1(new_n536), .B2(KEYINPUT4), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n286), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n482), .A2(G257), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n538), .A2(G190), .A3(new_n481), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n539), .ZN(new_n541));
  INV_X1    g0341(.A(new_n481), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n540), .B1(new_n543), .B2(new_n333), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT6), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n513), .A2(new_n217), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n546), .B2(new_n202), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n217), .A2(KEYINPUT6), .A3(G97), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n391), .A2(G107), .B1(G20), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n263), .A2(G77), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n259), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n469), .A2(G97), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n252), .A2(G97), .ZN(new_n555));
  XNOR2_X1  g0355(.A(new_n555), .B(KEYINPUT78), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT80), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n552), .A2(new_n259), .B1(G97), .B2(new_n469), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n560), .A2(KEYINPUT80), .A3(new_n556), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n544), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n469), .A2(G87), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT19), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n328), .B2(new_n513), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n279), .A2(new_n228), .A3(G68), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n228), .B1(new_n281), .B2(new_n564), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(G87), .B2(new_n203), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n569), .A2(new_n259), .B1(new_n400), .B2(new_n348), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n285), .B1(G250), .B2(new_n477), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n476), .A2(G1), .A3(G274), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OR2_X1    g0374(.A1(new_n317), .A2(G244), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(G238), .B2(G1698), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n576), .A2(new_n389), .B1(new_n261), .B2(new_n209), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n574), .B1(new_n286), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G190), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n571), .B(new_n579), .C1(new_n333), .C2(new_n578), .ZN(new_n580));
  INV_X1    g0380(.A(new_n578), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n426), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n578), .A2(new_n308), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n570), .B1(new_n348), .B2(new_n468), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n543), .A2(G179), .ZN(new_n587));
  OAI21_X1  g0387(.A(G169), .B1(new_n541), .B2(new_n542), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n587), .A2(new_n588), .B1(new_n560), .B2(new_n556), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n562), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  AND4_X1   g0390(.A1(new_n438), .A2(new_n498), .A3(new_n530), .A4(new_n590), .ZN(G372));
  INV_X1    g0391(.A(new_n310), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n315), .B2(new_n433), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n422), .B1(new_n419), .B2(KEYINPUT17), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n430), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n336), .ZN(new_n596));
  AND2_X1   g0396(.A1(new_n596), .A2(new_n338), .ZN(new_n597));
  INV_X1    g0397(.A(new_n585), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n559), .A2(new_n561), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n588), .B2(new_n587), .ZN(new_n600));
  XNOR2_X1  g0400(.A(new_n600), .B(KEYINPUT90), .ZN(new_n601));
  INV_X1    g0401(.A(new_n586), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT26), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n602), .A2(new_n589), .A3(KEYINPUT26), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n598), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n523), .A2(new_n522), .A3(new_n526), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n608), .A2(new_n497), .ZN(new_n609));
  NOR4_X1   g0409(.A1(new_n609), .A2(new_n491), .A3(new_n589), .A4(new_n562), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n602), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n597), .B1(new_n613), .B2(new_n437), .ZN(G369));
  INV_X1    g0414(.A(G13), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n615), .A2(G20), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n251), .ZN(new_n617));
  OR2_X1    g0417(.A1(new_n617), .A2(KEYINPUT27), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(KEYINPUT27), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n618), .A2(G213), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n620), .B(KEYINPUT91), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(G343), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n625), .A2(new_n528), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n608), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n626), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n627), .B1(new_n530), .B2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(G330), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n458), .A2(new_n470), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n624), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n498), .A2(new_n633), .B1(new_n497), .B2(new_n624), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n608), .A2(new_n625), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n498), .A2(new_n608), .A3(new_n625), .ZN(new_n638));
  AND2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n497), .A2(new_n625), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(G399));
  INV_X1    g0441(.A(new_n231), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n642), .A2(G41), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(G1), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n202), .A2(new_n372), .A3(new_n209), .ZN(new_n646));
  OAI22_X1  g0446(.A1(new_n645), .A2(new_n646), .B1(new_n227), .B2(new_n644), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n647), .B(KEYINPUT28), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n624), .B1(new_n607), .B2(new_n611), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT29), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n601), .A2(new_n580), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n598), .B1(new_n652), .B2(KEYINPUT26), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n589), .A2(new_n604), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n580), .B1(new_n610), .B2(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n624), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n651), .B1(new_n650), .B2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT30), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n487), .A2(new_n578), .A3(new_n538), .A4(new_n539), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n524), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n541), .A2(new_n581), .A3(new_n489), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n662), .A2(new_n525), .A3(KEYINPUT30), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n510), .A2(new_n308), .A3(new_n489), .A4(new_n581), .ZN(new_n664));
  OAI211_X1 g0464(.A(new_n661), .B(new_n663), .C1(new_n543), .C2(new_n664), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n665), .A2(KEYINPUT31), .A3(new_n624), .ZN(new_n666));
  AOI21_X1  g0466(.A(KEYINPUT31), .B1(new_n665), .B2(new_n624), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n498), .A2(new_n590), .A3(new_n530), .A4(new_n625), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G330), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT92), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n658), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n648), .B1(new_n673), .B2(G1), .ZN(G364));
  AOI21_X1  g0474(.A(new_n645), .B1(G45), .B2(new_n616), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(G13), .A2(G33), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(G20), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n676), .B1(new_n629), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(G20), .B1(KEYINPUT95), .B2(G169), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n681), .B1(KEYINPUT95), .B2(G169), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n229), .ZN(new_n683));
  OR3_X1    g0483(.A1(new_n333), .A2(KEYINPUT96), .A3(G179), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n228), .A2(G190), .ZN(new_n685));
  OAI21_X1  g0485(.A(KEYINPUT96), .B1(new_n333), .B2(G179), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n279), .B1(new_n688), .B2(G283), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n685), .A2(G179), .A3(G200), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  XNOR2_X1  g0491(.A(KEYINPUT33), .B(G317), .ZN(new_n692));
  NOR2_X1   g0492(.A1(G179), .A2(G200), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n685), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n691), .A2(new_n692), .B1(new_n695), .B2(G329), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n684), .A2(G20), .A3(G190), .A4(new_n686), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n698), .A2(KEYINPUT97), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(KEYINPUT97), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G303), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n689), .B(new_n696), .C1(new_n701), .C2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n375), .A2(G20), .A3(G179), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n333), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n685), .A2(G179), .A3(new_n333), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n705), .A2(G326), .B1(G311), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(G294), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n228), .B1(new_n693), .B2(G190), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT98), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n704), .A2(G200), .ZN(new_n713));
  AOI211_X1 g0513(.A(new_n703), .B(new_n712), .C1(G322), .C2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n688), .A2(G107), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n715), .B1(new_n701), .B2(new_n372), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n690), .A2(new_n225), .ZN(new_n717));
  INV_X1    g0517(.A(G77), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n706), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n694), .A2(new_n393), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT32), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n389), .B1(new_n713), .B2(G58), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n705), .A2(G50), .ZN(new_n723));
  INV_X1    g0523(.A(new_n710), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G97), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n721), .A2(new_n722), .A3(new_n723), .A4(new_n725), .ZN(new_n726));
  NOR4_X1   g0526(.A1(new_n716), .A2(new_n717), .A3(new_n719), .A4(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n683), .B1(new_n714), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n642), .A2(new_n389), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT94), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(G355), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n226), .A2(new_n476), .A3(G50), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n642), .A2(new_n279), .ZN(new_n733));
  OAI211_X1 g0533(.A(new_n732), .B(new_n733), .C1(new_n246), .C2(new_n476), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n731), .B(new_n734), .C1(G116), .C2(new_n231), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n683), .A2(new_n679), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n680), .A2(new_n728), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(KEYINPUT93), .B1(new_n629), .B2(new_n630), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n629), .A2(new_n630), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n739), .B(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n738), .B1(new_n741), .B2(new_n675), .ZN(G396));
  AOI22_X1  g0542(.A1(new_n713), .A2(G143), .B1(G150), .B2(new_n691), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(new_n393), .B2(new_n706), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(G137), .B2(new_n705), .ZN(new_n745));
  OAI22_X1  g0545(.A1(new_n745), .A2(KEYINPUT34), .B1(new_n224), .B2(new_n710), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(KEYINPUT34), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n279), .ZN(new_n748));
  AOI211_X1 g0548(.A(new_n746), .B(new_n748), .C1(G68), .C2(new_n688), .ZN(new_n749));
  INV_X1    g0549(.A(G50), .ZN(new_n750));
  INV_X1    g0550(.A(G132), .ZN(new_n751));
  OAI221_X1 g0551(.A(new_n749), .B1(new_n750), .B2(new_n701), .C1(new_n751), .C2(new_n694), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n687), .A2(new_n372), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n695), .A2(G311), .ZN(new_n754));
  INV_X1    g0554(.A(new_n705), .ZN(new_n755));
  OAI211_X1 g0555(.A(new_n725), .B(new_n754), .C1(new_n755), .C2(new_n702), .ZN(new_n756));
  XOR2_X1   g0556(.A(KEYINPUT99), .B(G283), .Z(new_n757));
  AOI211_X1 g0557(.A(new_n753), .B(new_n756), .C1(new_n691), .C2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n713), .A2(G294), .ZN(new_n759));
  INV_X1    g0559(.A(new_n701), .ZN(new_n760));
  AOI22_X1  g0560(.A1(new_n760), .A2(G107), .B1(G116), .B2(new_n707), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n758), .A2(new_n389), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT100), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n752), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n676), .B1(new_n764), .B2(new_n683), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n433), .A2(new_n625), .ZN(new_n766));
  AOI22_X1  g0566(.A1(new_n355), .A2(new_n345), .B1(new_n351), .B2(new_n624), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n766), .B1(new_n767), .B2(new_n433), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n765), .B1(new_n769), .B2(new_n678), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n683), .A2(new_n677), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n770), .B1(new_n718), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT101), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n672), .B(new_n769), .ZN(new_n774));
  XNOR2_X1  g0574(.A(new_n774), .B(new_n649), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n773), .B1(new_n775), .B2(new_n676), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(G384));
  NAND2_X1  g0577(.A1(new_n624), .A2(new_n272), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n310), .A2(new_n315), .A3(new_n778), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n272), .B(new_n624), .C1(new_n306), .C2(new_n309), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n767), .A2(new_n433), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n649), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n782), .B1(new_n784), .B2(new_n766), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT38), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n260), .B1(new_n411), .B2(new_n412), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n621), .B1(new_n787), .B2(new_n402), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(new_n424), .B2(new_n430), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n399), .A2(new_n403), .B1(new_n426), .B2(new_n379), .ZN(new_n790));
  AOI221_X4 g0590(.A(KEYINPUT37), .B1(new_n790), .B2(new_n425), .C1(new_n405), .C2(new_n418), .ZN(new_n791));
  INV_X1    g0591(.A(KEYINPUT102), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n788), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n404), .A2(KEYINPUT102), .A3(new_n621), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n421), .A2(new_n357), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n360), .A2(new_n363), .A3(new_n358), .ZN(new_n798));
  AOI21_X1  g0598(.A(KEYINPUT75), .B1(new_n366), .B2(new_n367), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n378), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n379), .A2(new_n333), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(KEYINPUT77), .B1(new_n802), .B2(new_n414), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n428), .B(new_n788), .C1(new_n797), .C2(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n791), .A2(new_n796), .B1(new_n804), .B2(KEYINPUT37), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n786), .B1(new_n789), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(KEYINPUT37), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT37), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n796), .A2(new_n419), .A3(new_n808), .A4(new_n428), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n788), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n594), .B2(new_n429), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n810), .A2(new_n812), .A3(KEYINPUT38), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n806), .A2(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n785), .A2(new_n814), .B1(new_n429), .B2(new_n622), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n310), .A2(new_n624), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  AND3_X1   g0617(.A1(new_n428), .A2(KEYINPUT103), .A3(new_n421), .ZN(new_n818));
  AOI21_X1  g0618(.A(KEYINPUT103), .B1(new_n428), .B2(new_n421), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n818), .A2(new_n819), .A3(new_n795), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n809), .B1(new_n820), .B2(new_n808), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n795), .B1(new_n594), .B2(new_n429), .ZN(new_n822));
  AOI21_X1  g0622(.A(KEYINPUT38), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AND3_X1   g0623(.A1(new_n810), .A2(new_n812), .A3(KEYINPUT38), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT39), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n806), .A2(KEYINPUT39), .A3(new_n813), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n815), .B1(new_n817), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n597), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(new_n658), .B2(new_n438), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n830), .B(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n437), .B1(new_n669), .B2(new_n668), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n768), .B1(new_n779), .B2(new_n780), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n670), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(KEYINPUT38), .B1(new_n810), .B2(new_n812), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n836), .B1(new_n824), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT40), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OAI211_X1 g0640(.A(KEYINPUT40), .B(new_n836), .C1(new_n823), .C2(new_n824), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n834), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(G330), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n833), .B(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n251), .B2(new_n616), .ZN(new_n846));
  OAI211_X1 g0646(.A(G20), .B(new_n283), .C1(new_n549), .C2(KEYINPUT35), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n209), .B(new_n847), .C1(KEYINPUT35), .C2(new_n549), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT36), .Z(new_n849));
  NAND2_X1  g0649(.A1(new_n382), .A2(G77), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n227), .A2(new_n850), .B1(G50), .B2(new_n225), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n851), .A2(G1), .A3(new_n615), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n846), .A2(new_n849), .A3(new_n852), .ZN(G367));
  AOI21_X1  g0653(.A(new_n251), .B1(new_n616), .B2(G45), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n673), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n639), .B1(new_n631), .B2(new_n636), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n562), .A2(new_n589), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n859), .B1(new_n599), .B2(new_n625), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n600), .A2(new_n624), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n638), .A2(new_n640), .ZN(new_n863));
  OR3_X1    g0663(.A1(new_n862), .A2(new_n863), .A3(KEYINPUT106), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT106), .B1(new_n862), .B2(new_n863), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n866), .A2(KEYINPUT45), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n862), .A2(new_n863), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT44), .Z(new_n869));
  NAND2_X1  g0669(.A1(new_n866), .A2(KEYINPUT45), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n637), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n858), .A2(KEYINPUT107), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n673), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n643), .B(KEYINPUT41), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n855), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OR2_X1    g0677(.A1(new_n638), .A2(new_n860), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT42), .ZN(new_n879));
  INV_X1    g0679(.A(new_n862), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n589), .B1(new_n880), .B2(new_n497), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n879), .B1(new_n881), .B2(new_n624), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n882), .B(KEYINPUT104), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n878), .A2(KEYINPUT42), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n872), .A2(new_n880), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n886), .B(KEYINPUT105), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n625), .A2(new_n571), .ZN(new_n889));
  OR2_X1    g0689(.A1(new_n889), .A2(new_n585), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n602), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT43), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n885), .A2(new_n888), .A3(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n888), .B1(new_n885), .B2(new_n894), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n892), .A2(KEYINPUT43), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n898), .B(new_n900), .ZN(new_n901));
  OR3_X1    g0701(.A1(new_n877), .A2(new_n901), .A3(KEYINPUT108), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT108), .B1(new_n877), .B2(new_n901), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n688), .A2(G77), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n695), .A2(G137), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n905), .B(new_n906), .C1(new_n750), .C2(new_n706), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n389), .B(new_n907), .C1(new_n760), .C2(G58), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n713), .A2(G150), .B1(G68), .B2(new_n724), .ZN(new_n909));
  INV_X1    g0709(.A(G143), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n908), .B(new_n909), .C1(new_n910), .C2(new_n755), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(G159), .B2(new_n691), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT46), .B1(new_n760), .B2(G116), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n760), .A2(KEYINPUT46), .A3(G116), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n713), .A2(G303), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n690), .A2(new_n709), .B1(new_n710), .B2(new_n217), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n687), .A2(new_n513), .ZN(new_n917));
  AOI211_X1 g0717(.A(new_n916), .B(new_n917), .C1(G317), .C2(new_n695), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n279), .B1(new_n705), .B2(G311), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n914), .A2(new_n915), .A3(new_n918), .A4(new_n919), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n913), .B(new_n920), .C1(new_n707), .C2(new_n757), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n912), .A2(new_n921), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT47), .Z(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n683), .ZN(new_n924));
  INV_X1    g0724(.A(new_n733), .ZN(new_n925));
  OAI221_X1 g0725(.A(new_n736), .B1(new_n231), .B2(new_n348), .C1(new_n237), .C2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n890), .A2(new_n679), .A3(new_n891), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n924), .A2(new_n675), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n904), .A2(new_n928), .ZN(G387));
  XOR2_X1   g0729(.A(KEYINPUT109), .B(G322), .Z(new_n930));
  NOR2_X1   g0730(.A1(new_n755), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(G311), .B2(new_n691), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n702), .B2(new_n706), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(G317), .B2(new_n713), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT48), .Z(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n709), .B2(new_n701), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n724), .B2(new_n757), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT49), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n389), .B1(new_n687), .B2(new_n209), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(G326), .B2(new_n695), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT110), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n701), .A2(new_n718), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n713), .A2(G50), .B1(new_n346), .B2(new_n691), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n327), .B2(new_n694), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n710), .A2(new_n348), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n389), .B1(new_n707), .B2(G68), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n946), .B(new_n947), .C1(new_n755), .C2(new_n393), .ZN(new_n948));
  NOR4_X1   g0748(.A1(new_n943), .A2(new_n917), .A3(new_n945), .A4(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n683), .B1(new_n942), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n733), .B1(new_n242), .B2(new_n476), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n730), .A2(new_n646), .ZN(new_n952));
  AOI211_X1 g0752(.A(G45), .B(new_n646), .C1(G68), .C2(G77), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n329), .A2(G50), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT50), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n951), .A2(new_n952), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n231), .A2(G107), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n736), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n676), .B1(new_n634), .B2(new_n679), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n950), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n857), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n643), .B1(new_n673), .B2(new_n961), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n960), .B1(new_n854), .B2(new_n857), .C1(new_n858), .C2(new_n962), .ZN(G393));
  NAND2_X1  g0763(.A1(new_n873), .A2(KEYINPUT111), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n871), .A2(new_n872), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n964), .B(new_n965), .Z(new_n966));
  OAI211_X1 g0766(.A(new_n643), .B(new_n874), .C1(new_n966), .C2(new_n858), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n930), .A2(new_n694), .ZN(new_n968));
  AOI22_X1  g0768(.A1(G311), .A2(new_n713), .B1(new_n705), .B2(G317), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT112), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT52), .Z(new_n971));
  OAI221_X1 g0771(.A(new_n715), .B1(new_n709), .B2(new_n706), .C1(new_n702), .C2(new_n690), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n972), .B1(new_n760), .B2(new_n757), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n971), .A2(new_n389), .A3(new_n973), .ZN(new_n974));
  AOI211_X1 g0774(.A(new_n968), .B(new_n974), .C1(G116), .C2(new_n724), .ZN(new_n975));
  AOI22_X1  g0775(.A1(G150), .A2(new_n705), .B1(new_n713), .B2(G159), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n976), .B(KEYINPUT51), .Z(new_n977));
  OAI221_X1 g0777(.A(new_n977), .B1(new_n910), .B2(new_n694), .C1(new_n329), .C2(new_n706), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n710), .A2(new_n718), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n701), .A2(new_n225), .B1(new_n372), .B2(new_n687), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n279), .B1(new_n690), .B2(new_n750), .ZN(new_n981));
  NOR4_X1   g0781(.A1(new_n978), .A2(new_n979), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n683), .B1(new_n975), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n862), .A2(new_n679), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n736), .B1(new_n513), .B2(new_n231), .C1(new_n249), .C2(new_n925), .ZN(new_n985));
  AND4_X1   g0785(.A1(new_n675), .A2(new_n983), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(new_n966), .B2(new_n855), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n967), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT113), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n967), .A2(KEYINPUT113), .A3(new_n987), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(G390));
  OAI21_X1  g0792(.A(new_n829), .B1(new_n785), .B2(new_n816), .ZN(new_n993));
  INV_X1    g0793(.A(new_n766), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(new_n657), .B2(new_n783), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n995), .A2(new_n782), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n825), .A2(new_n817), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n993), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n670), .A2(new_n835), .A3(G330), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT114), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n672), .A2(new_n835), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1000), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT115), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n834), .A2(G330), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n832), .A2(new_n1010), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n649), .A2(new_n783), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n781), .B1(new_n672), .B2(new_n769), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n1012), .A2(new_n994), .B1(new_n1002), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n782), .B1(new_n671), .B2(new_n768), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n995), .A2(new_n1005), .A3(new_n1015), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1011), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1008), .B1(new_n1009), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1018), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1020), .B(KEYINPUT115), .C1(new_n1004), .C2(new_n1007), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1019), .A2(new_n643), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n771), .A2(new_n329), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n760), .A2(G150), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT53), .ZN(new_n1025));
  XOR2_X1   g0825(.A(KEYINPUT54), .B(G143), .Z(new_n1026));
  AOI211_X1 g0826(.A(new_n389), .B(new_n1025), .C1(new_n707), .C2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n695), .A2(G125), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n691), .A2(G137), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n713), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n1030), .A2(new_n751), .B1(new_n687), .B2(new_n750), .ZN(new_n1031));
  INV_X1    g0831(.A(G128), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n755), .A2(new_n1032), .B1(new_n393), .B2(new_n710), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n694), .A2(new_n709), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n760), .A2(G87), .B1(G68), .B2(new_n688), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n979), .B1(G107), .B2(new_n691), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n1030), .B2(new_n209), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n279), .B(new_n1039), .C1(G97), .C2(new_n707), .ZN(new_n1040));
  INV_X1    g0840(.A(G283), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1037), .B(new_n1040), .C1(new_n1041), .C2(new_n755), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1035), .B1(new_n1036), .B2(new_n1042), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n1043), .A2(new_n683), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n676), .B(new_n1044), .C1(new_n829), .C2(new_n677), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n1008), .A2(new_n855), .B1(new_n1023), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1022), .A2(new_n1046), .ZN(G378));
  XOR2_X1   g0847(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n336), .B2(new_n338), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n336), .A2(new_n338), .A3(new_n1049), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1051), .A2(new_n332), .A3(new_n621), .A4(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n621), .A2(new_n332), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1052), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1054), .B1(new_n1055), .B2(new_n1050), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n677), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n771), .A2(new_n750), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(G33), .A2(G41), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT116), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1062), .B(new_n750), .C1(G41), .C2(new_n279), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n760), .A2(new_n1026), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n691), .A2(G132), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n705), .A2(G125), .B1(G137), .B2(new_n707), .ZN(new_n1066));
  AND3_X1   g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n1032), .B2(new_n1030), .C1(new_n327), .C2(new_n710), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1068), .A2(KEYINPUT59), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1062), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n695), .A2(G124), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1068), .A2(KEYINPUT59), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n687), .A2(new_n393), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1063), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n687), .A2(new_n224), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT117), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n701), .B2(new_n718), .ZN(new_n1078));
  AOI211_X1 g0878(.A(G41), .B(new_n279), .C1(new_n724), .C2(G68), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n1041), .B2(new_n694), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n755), .A2(new_n209), .B1(new_n513), .B2(new_n690), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n1078), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n217), .B2(new_n1030), .C1(new_n348), .C2(new_n706), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT58), .Z(new_n1084));
  OAI21_X1  g0884(.A(new_n683), .B1(new_n1075), .B2(new_n1084), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1059), .A2(new_n675), .A3(new_n1060), .A4(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n670), .A2(new_n835), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n806), .B2(new_n813), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n841), .B(G330), .C1(KEYINPUT40), .C2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT118), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n840), .A2(KEYINPUT118), .A3(G330), .A4(new_n841), .ZN(new_n1093));
  AND4_X1   g0893(.A1(KEYINPUT119), .A2(new_n1092), .A3(new_n1058), .A4(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1057), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1095));
  AOI21_X1  g0895(.A(KEYINPUT119), .B1(new_n1095), .B2(new_n1093), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1058), .A2(new_n1090), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT120), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1092), .A2(new_n1058), .A3(new_n1093), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT119), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1095), .A2(KEYINPUT119), .A3(new_n1093), .ZN(new_n1103));
  AND4_X1   g0903(.A1(KEYINPUT120), .A2(new_n1102), .A3(new_n1098), .A4(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n830), .B1(new_n1099), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT121), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1102), .A2(new_n1098), .A3(new_n1103), .ZN(new_n1108));
  OR2_X1    g0908(.A1(new_n830), .A2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g0909(.A(KEYINPUT121), .B(new_n830), .C1(new_n1099), .C2(new_n1104), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1087), .B1(new_n1111), .B2(new_n855), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1011), .A2(KEYINPUT122), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n1011), .A2(KEYINPUT122), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1003), .B1(new_n1006), .B2(new_n1000), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1113), .B(new_n1114), .C1(new_n1115), .C2(new_n1020), .ZN(new_n1116));
  AOI21_X1  g0916(.A(KEYINPUT57), .B1(new_n1111), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT123), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n830), .B2(new_n1108), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n1109), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1109), .A2(new_n1119), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1116), .A2(new_n1120), .A3(KEYINPUT57), .A4(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n643), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1112), .B1(new_n1117), .B2(new_n1123), .ZN(G375));
  NAND2_X1  g0924(.A1(new_n905), .A2(new_n389), .ZN(new_n1125));
  XOR2_X1   g0925(.A(new_n1125), .B(KEYINPUT124), .Z(new_n1126));
  OAI221_X1 g0926(.A(new_n1126), .B1(new_n513), .B2(new_n701), .C1(new_n217), .C2(new_n706), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n755), .A2(new_n709), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n1030), .A2(new_n1041), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n946), .B1(new_n209), .B2(new_n690), .C1(new_n702), .C2(new_n694), .ZN(new_n1130));
  NOR4_X1   g0930(.A1(new_n1127), .A2(new_n1128), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n691), .A2(new_n1026), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n701), .B2(new_n393), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n713), .A2(G137), .B1(G128), .B2(new_n695), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n389), .B1(new_n707), .B2(G150), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1077), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n710), .A2(new_n750), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n755), .A2(new_n751), .ZN(new_n1138));
  NOR4_X1   g0938(.A1(new_n1133), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n683), .B1(new_n1131), .B2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n675), .B(new_n1140), .C1(new_n781), .C2(new_n678), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(new_n225), .B2(new_n771), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1017), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1142), .B1(new_n1143), .B2(new_n855), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1011), .A2(new_n1017), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n876), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1144), .B1(new_n1146), .B2(new_n1018), .ZN(G381));
  NAND4_X1  g0947(.A1(new_n904), .A2(new_n990), .A3(new_n928), .A4(new_n991), .ZN(new_n1148));
  OR2_X1    g0948(.A1(G381), .A2(G384), .ZN(new_n1149));
  NOR4_X1   g0949(.A1(new_n1148), .A2(G396), .A3(G393), .A4(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(G378), .ZN(new_n1151));
  INV_X1    g0951(.A(G375), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(G407));
  NAND2_X1  g0953(.A1(new_n623), .A2(G213), .ZN(new_n1154));
  XOR2_X1   g0954(.A(new_n1154), .B(KEYINPUT125), .Z(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1150), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1152), .A2(new_n1151), .ZN(new_n1158));
  OAI21_X1  g0958(.A(G213), .B1(new_n1157), .B2(new_n1158), .ZN(G409));
  INV_X1    g0959(.A(KEYINPUT61), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1111), .A2(new_n876), .A3(new_n1116), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1120), .A2(new_n855), .A3(new_n1121), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1161), .A2(new_n1086), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1163), .A2(new_n1151), .ZN(new_n1164));
  OAI211_X1 g0964(.A(G378), .B(new_n1112), .C1(new_n1117), .C2(new_n1123), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1156), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT60), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n644), .B1(new_n1145), .B2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1168), .B(new_n1020), .C1(new_n1167), .C2(new_n1145), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n1144), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n776), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1169), .A2(G384), .A3(new_n1144), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1173), .A2(G2897), .A3(new_n1156), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1154), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1175), .A2(G2897), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1174), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1160), .B1(new_n1166), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(KEYINPUT126), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1173), .ZN(new_n1180));
  AND2_X1   g0980(.A1(new_n1180), .A2(KEYINPUT62), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1166), .A2(new_n1181), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1175), .B(new_n1173), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1182), .B1(new_n1183), .B2(KEYINPUT62), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT126), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1185), .B(new_n1160), .C1(new_n1166), .C2(new_n1177), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1179), .A2(new_n1184), .A3(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(G393), .B(G396), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1148), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n904), .A2(new_n928), .B1(new_n990), .B2(new_n991), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1189), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1191), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1193), .A2(new_n1148), .A3(new_n1188), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1187), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1183), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1175), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1198));
  OAI21_X1  g0998(.A(KEYINPUT63), .B1(new_n1198), .B2(new_n1177), .ZN(new_n1199));
  AOI21_X1  g0999(.A(KEYINPUT61), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1195), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1166), .A2(KEYINPUT63), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(new_n1180), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1200), .A2(new_n1201), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1196), .A2(new_n1204), .ZN(G405));
  NAND2_X1  g1005(.A1(G375), .A2(new_n1151), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1180), .A2(KEYINPUT127), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1206), .A2(new_n1165), .A3(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1180), .A2(KEYINPUT127), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1208), .B(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(new_n1201), .ZN(G402));
endmodule


