

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U552 ( .A1(G164), .A2(G1384), .ZN(n693) );
  INV_X1 U553 ( .A(KEYINPUT27), .ZN(n709) );
  XNOR2_X1 U554 ( .A(n710), .B(n709), .ZN(n712) );
  INV_X1 U555 ( .A(n740), .ZN(n720) );
  INV_X1 U556 ( .A(KEYINPUT28), .ZN(n730) );
  XNOR2_X1 U557 ( .A(KEYINPUT31), .B(KEYINPUT97), .ZN(n705) );
  XNOR2_X1 U558 ( .A(n706), .B(n705), .ZN(n739) );
  NAND2_X1 U559 ( .A1(n694), .A2(n693), .ZN(n740) );
  INV_X1 U560 ( .A(n779), .ZN(n764) );
  XNOR2_X1 U561 ( .A(n699), .B(KEYINPUT90), .ZN(n779) );
  NAND2_X1 U562 ( .A1(G160), .A2(G40), .ZN(n692) );
  NOR2_X1 U563 ( .A1(G651), .A2(G543), .ZN(n633) );
  NOR2_X1 U564 ( .A1(G2104), .A2(n520), .ZN(n868) );
  NOR2_X1 U565 ( .A1(n545), .A2(n544), .ZN(G160) );
  XNOR2_X1 U566 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n517) );
  NOR2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n516) );
  XNOR2_X2 U568 ( .A(n517), .B(n516), .ZN(n873) );
  NAND2_X1 U569 ( .A1(G138), .A2(n873), .ZN(n519) );
  INV_X1 U570 ( .A(G2105), .ZN(n520) );
  AND2_X4 U571 ( .A1(n520), .A2(G2104), .ZN(n872) );
  NAND2_X1 U572 ( .A1(G102), .A2(n872), .ZN(n518) );
  NAND2_X1 U573 ( .A1(n519), .A2(n518), .ZN(n524) );
  NAND2_X1 U574 ( .A1(G126), .A2(n868), .ZN(n522) );
  AND2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n869) );
  NAND2_X1 U576 ( .A1(G114), .A2(n869), .ZN(n521) );
  NAND2_X1 U577 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U578 ( .A1(n524), .A2(n523), .ZN(G164) );
  INV_X1 U579 ( .A(G651), .ZN(n531) );
  NOR2_X1 U580 ( .A1(G543), .A2(n531), .ZN(n525) );
  XOR2_X1 U581 ( .A(KEYINPUT1), .B(n525), .Z(n638) );
  NAND2_X1 U582 ( .A1(G63), .A2(n638), .ZN(n528) );
  XOR2_X1 U583 ( .A(KEYINPUT0), .B(G543), .Z(n617) );
  NOR2_X1 U584 ( .A1(G651), .A2(n617), .ZN(n526) );
  XNOR2_X1 U585 ( .A(KEYINPUT64), .B(n526), .ZN(n635) );
  NAND2_X1 U586 ( .A1(G51), .A2(n635), .ZN(n527) );
  NAND2_X1 U587 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U588 ( .A(KEYINPUT6), .B(n529), .ZN(n537) );
  NAND2_X1 U589 ( .A1(n633), .A2(G89), .ZN(n530) );
  XNOR2_X1 U590 ( .A(n530), .B(KEYINPUT4), .ZN(n533) );
  NOR2_X1 U591 ( .A1(n617), .A2(n531), .ZN(n631) );
  NAND2_X1 U592 ( .A1(G76), .A2(n631), .ZN(n532) );
  NAND2_X1 U593 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U594 ( .A(KEYINPUT5), .B(n534), .ZN(n535) );
  XNOR2_X1 U595 ( .A(KEYINPUT71), .B(n535), .ZN(n536) );
  NOR2_X1 U596 ( .A1(n537), .A2(n536), .ZN(n538) );
  XOR2_X1 U597 ( .A(KEYINPUT7), .B(n538), .Z(G168) );
  XOR2_X1 U598 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U599 ( .A1(n873), .A2(G137), .ZN(n541) );
  NAND2_X1 U600 ( .A1(G101), .A2(n872), .ZN(n539) );
  XOR2_X1 U601 ( .A(KEYINPUT23), .B(n539), .Z(n540) );
  NAND2_X1 U602 ( .A1(n541), .A2(n540), .ZN(n545) );
  NAND2_X1 U603 ( .A1(G125), .A2(n868), .ZN(n543) );
  NAND2_X1 U604 ( .A1(G113), .A2(n869), .ZN(n542) );
  NAND2_X1 U605 ( .A1(n543), .A2(n542), .ZN(n544) );
  NAND2_X1 U606 ( .A1(G85), .A2(n633), .ZN(n547) );
  NAND2_X1 U607 ( .A1(G60), .A2(n638), .ZN(n546) );
  NAND2_X1 U608 ( .A1(n547), .A2(n546), .ZN(n551) );
  NAND2_X1 U609 ( .A1(G72), .A2(n631), .ZN(n549) );
  NAND2_X1 U610 ( .A1(G47), .A2(n635), .ZN(n548) );
  NAND2_X1 U611 ( .A1(n549), .A2(n548), .ZN(n550) );
  OR2_X1 U612 ( .A1(n551), .A2(n550), .ZN(G290) );
  AND2_X1 U613 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U614 ( .A(G82), .ZN(G220) );
  INV_X1 U615 ( .A(G57), .ZN(G237) );
  NAND2_X1 U616 ( .A1(G64), .A2(n638), .ZN(n553) );
  NAND2_X1 U617 ( .A1(G52), .A2(n635), .ZN(n552) );
  NAND2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n558) );
  NAND2_X1 U619 ( .A1(G77), .A2(n631), .ZN(n555) );
  NAND2_X1 U620 ( .A1(G90), .A2(n633), .ZN(n554) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U622 ( .A(KEYINPUT9), .B(n556), .Z(n557) );
  NOR2_X1 U623 ( .A1(n558), .A2(n557), .ZN(G171) );
  XOR2_X1 U624 ( .A(KEYINPUT10), .B(KEYINPUT67), .Z(n560) );
  NAND2_X1 U625 ( .A1(G7), .A2(G661), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(G223) );
  INV_X1 U627 ( .A(G223), .ZN(n816) );
  NAND2_X1 U628 ( .A1(n816), .A2(G567), .ZN(n561) );
  XOR2_X1 U629 ( .A(KEYINPUT11), .B(n561), .Z(G234) );
  XOR2_X1 U630 ( .A(G860), .B(KEYINPUT68), .Z(n590) );
  NAND2_X1 U631 ( .A1(G56), .A2(n638), .ZN(n562) );
  XOR2_X1 U632 ( .A(KEYINPUT14), .B(n562), .Z(n568) );
  NAND2_X1 U633 ( .A1(n633), .A2(G81), .ZN(n563) );
  XNOR2_X1 U634 ( .A(n563), .B(KEYINPUT12), .ZN(n565) );
  NAND2_X1 U635 ( .A1(G68), .A2(n631), .ZN(n564) );
  NAND2_X1 U636 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U637 ( .A(KEYINPUT13), .B(n566), .Z(n567) );
  NOR2_X1 U638 ( .A1(n568), .A2(n567), .ZN(n570) );
  NAND2_X1 U639 ( .A1(G43), .A2(n635), .ZN(n569) );
  NAND2_X1 U640 ( .A1(n570), .A2(n569), .ZN(n997) );
  OR2_X1 U641 ( .A1(n590), .A2(n997), .ZN(G153) );
  INV_X1 U642 ( .A(G171), .ZN(G301) );
  INV_X1 U643 ( .A(G868), .ZN(n652) );
  NOR2_X1 U644 ( .A1(G301), .A2(n652), .ZN(n580) );
  NAND2_X1 U645 ( .A1(n635), .A2(G54), .ZN(n577) );
  NAND2_X1 U646 ( .A1(G92), .A2(n633), .ZN(n572) );
  NAND2_X1 U647 ( .A1(G66), .A2(n638), .ZN(n571) );
  NAND2_X1 U648 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U649 ( .A1(G79), .A2(n631), .ZN(n573) );
  XNOR2_X1 U650 ( .A(KEYINPUT69), .B(n573), .ZN(n574) );
  NOR2_X1 U651 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U652 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U653 ( .A(n578), .B(KEYINPUT15), .ZN(n1009) );
  AND2_X1 U654 ( .A1(n652), .A2(n1009), .ZN(n579) );
  NOR2_X1 U655 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U656 ( .A(KEYINPUT70), .B(n581), .ZN(G284) );
  NAND2_X1 U657 ( .A1(G65), .A2(n638), .ZN(n583) );
  NAND2_X1 U658 ( .A1(G53), .A2(n635), .ZN(n582) );
  NAND2_X1 U659 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U660 ( .A1(G78), .A2(n631), .ZN(n585) );
  NAND2_X1 U661 ( .A1(G91), .A2(n633), .ZN(n584) );
  NAND2_X1 U662 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U663 ( .A1(n587), .A2(n586), .ZN(n988) );
  INV_X1 U664 ( .A(n988), .ZN(G299) );
  NOR2_X1 U665 ( .A1(G286), .A2(n652), .ZN(n589) );
  NOR2_X1 U666 ( .A1(G868), .A2(G299), .ZN(n588) );
  NOR2_X1 U667 ( .A1(n589), .A2(n588), .ZN(G297) );
  NAND2_X1 U668 ( .A1(n590), .A2(G559), .ZN(n591) );
  NAND2_X1 U669 ( .A1(n591), .A2(n1009), .ZN(n592) );
  XNOR2_X1 U670 ( .A(n592), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U671 ( .A1(G868), .A2(n997), .ZN(n595) );
  NAND2_X1 U672 ( .A1(G868), .A2(n1009), .ZN(n593) );
  NOR2_X1 U673 ( .A1(G559), .A2(n593), .ZN(n594) );
  NOR2_X1 U674 ( .A1(n595), .A2(n594), .ZN(G282) );
  NAND2_X1 U675 ( .A1(G123), .A2(n868), .ZN(n596) );
  XNOR2_X1 U676 ( .A(n596), .B(KEYINPUT72), .ZN(n597) );
  XNOR2_X1 U677 ( .A(KEYINPUT18), .B(n597), .ZN(n600) );
  NAND2_X1 U678 ( .A1(G111), .A2(n869), .ZN(n598) );
  XOR2_X1 U679 ( .A(KEYINPUT73), .B(n598), .Z(n599) );
  NAND2_X1 U680 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U681 ( .A1(G99), .A2(n872), .ZN(n602) );
  NAND2_X1 U682 ( .A1(G135), .A2(n873), .ZN(n601) );
  NAND2_X1 U683 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U684 ( .A1(n604), .A2(n603), .ZN(n918) );
  XOR2_X1 U685 ( .A(n918), .B(G2096), .Z(n605) );
  NOR2_X1 U686 ( .A1(G2100), .A2(n605), .ZN(n606) );
  XOR2_X1 U687 ( .A(KEYINPUT74), .B(n606), .Z(G156) );
  NAND2_X1 U688 ( .A1(G67), .A2(n638), .ZN(n607) );
  XNOR2_X1 U689 ( .A(n607), .B(KEYINPUT76), .ZN(n614) );
  NAND2_X1 U690 ( .A1(G80), .A2(n631), .ZN(n609) );
  NAND2_X1 U691 ( .A1(G55), .A2(n635), .ZN(n608) );
  NAND2_X1 U692 ( .A1(n609), .A2(n608), .ZN(n612) );
  NAND2_X1 U693 ( .A1(G93), .A2(n633), .ZN(n610) );
  XNOR2_X1 U694 ( .A(KEYINPUT75), .B(n610), .ZN(n611) );
  NOR2_X1 U695 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U696 ( .A1(n614), .A2(n613), .ZN(n653) );
  NAND2_X1 U697 ( .A1(n1009), .A2(G559), .ZN(n650) );
  XNOR2_X1 U698 ( .A(n997), .B(n650), .ZN(n615) );
  NOR2_X1 U699 ( .A1(G860), .A2(n615), .ZN(n616) );
  XOR2_X1 U700 ( .A(n653), .B(n616), .Z(G145) );
  NAND2_X1 U701 ( .A1(n617), .A2(G87), .ZN(n618) );
  XNOR2_X1 U702 ( .A(n618), .B(KEYINPUT78), .ZN(n620) );
  NAND2_X1 U703 ( .A1(G74), .A2(G651), .ZN(n619) );
  NAND2_X1 U704 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U705 ( .A1(n638), .A2(n621), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n635), .A2(G49), .ZN(n622) );
  XOR2_X1 U707 ( .A(KEYINPUT77), .B(n622), .Z(n623) );
  NAND2_X1 U708 ( .A1(n624), .A2(n623), .ZN(G288) );
  NAND2_X1 U709 ( .A1(G75), .A2(n631), .ZN(n626) );
  NAND2_X1 U710 ( .A1(G88), .A2(n633), .ZN(n625) );
  NAND2_X1 U711 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U712 ( .A1(G62), .A2(n638), .ZN(n628) );
  NAND2_X1 U713 ( .A1(G50), .A2(n635), .ZN(n627) );
  NAND2_X1 U714 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U715 ( .A1(n630), .A2(n629), .ZN(G166) );
  NAND2_X1 U716 ( .A1(n631), .A2(G73), .ZN(n632) );
  XNOR2_X1 U717 ( .A(KEYINPUT2), .B(n632), .ZN(n643) );
  NAND2_X1 U718 ( .A1(G86), .A2(n633), .ZN(n634) );
  XNOR2_X1 U719 ( .A(n634), .B(KEYINPUT80), .ZN(n637) );
  NAND2_X1 U720 ( .A1(G48), .A2(n635), .ZN(n636) );
  NAND2_X1 U721 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U722 ( .A1(G61), .A2(n638), .ZN(n639) );
  XNOR2_X1 U723 ( .A(KEYINPUT79), .B(n639), .ZN(n640) );
  NOR2_X1 U724 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U725 ( .A1(n643), .A2(n642), .ZN(G305) );
  XNOR2_X1 U726 ( .A(G290), .B(KEYINPUT19), .ZN(n645) );
  XNOR2_X1 U727 ( .A(n988), .B(G166), .ZN(n644) );
  XNOR2_X1 U728 ( .A(n645), .B(n644), .ZN(n646) );
  XOR2_X1 U729 ( .A(n646), .B(n997), .Z(n647) );
  XNOR2_X1 U730 ( .A(G288), .B(n647), .ZN(n649) );
  XOR2_X1 U731 ( .A(G305), .B(n653), .Z(n648) );
  XNOR2_X1 U732 ( .A(n649), .B(n648), .ZN(n890) );
  XOR2_X1 U733 ( .A(n890), .B(n650), .Z(n651) );
  NAND2_X1 U734 ( .A1(G868), .A2(n651), .ZN(n655) );
  NAND2_X1 U735 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U736 ( .A1(n655), .A2(n654), .ZN(G295) );
  NAND2_X1 U737 ( .A1(G2078), .A2(G2084), .ZN(n656) );
  XOR2_X1 U738 ( .A(KEYINPUT20), .B(n656), .Z(n657) );
  NAND2_X1 U739 ( .A1(G2090), .A2(n657), .ZN(n658) );
  XNOR2_X1 U740 ( .A(KEYINPUT21), .B(n658), .ZN(n659) );
  NAND2_X1 U741 ( .A1(n659), .A2(G2072), .ZN(G158) );
  XOR2_X1 U742 ( .A(KEYINPUT66), .B(G132), .Z(G219) );
  XNOR2_X1 U743 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U744 ( .A1(G69), .A2(G120), .ZN(n660) );
  NOR2_X1 U745 ( .A1(G237), .A2(n660), .ZN(n661) );
  NAND2_X1 U746 ( .A1(G108), .A2(n661), .ZN(n820) );
  NAND2_X1 U747 ( .A1(G567), .A2(n820), .ZN(n662) );
  XNOR2_X1 U748 ( .A(n662), .B(KEYINPUT82), .ZN(n668) );
  NOR2_X1 U749 ( .A1(G219), .A2(G220), .ZN(n664) );
  XNOR2_X1 U750 ( .A(KEYINPUT22), .B(KEYINPUT81), .ZN(n663) );
  XNOR2_X1 U751 ( .A(n664), .B(n663), .ZN(n665) );
  NOR2_X1 U752 ( .A1(n665), .A2(G218), .ZN(n666) );
  NAND2_X1 U753 ( .A1(G96), .A2(n666), .ZN(n821) );
  NAND2_X1 U754 ( .A1(G2106), .A2(n821), .ZN(n667) );
  NAND2_X1 U755 ( .A1(n668), .A2(n667), .ZN(n822) );
  NAND2_X1 U756 ( .A1(G661), .A2(G483), .ZN(n669) );
  NOR2_X1 U757 ( .A1(n822), .A2(n669), .ZN(n819) );
  NAND2_X1 U758 ( .A1(n819), .A2(G36), .ZN(G176) );
  INV_X1 U759 ( .A(G166), .ZN(G303) );
  NOR2_X1 U760 ( .A1(n693), .A2(n692), .ZN(n670) );
  XOR2_X1 U761 ( .A(KEYINPUT83), .B(n670), .Z(n811) );
  INV_X1 U762 ( .A(n811), .ZN(n691) );
  NAND2_X1 U763 ( .A1(G105), .A2(n872), .ZN(n671) );
  XOR2_X1 U764 ( .A(KEYINPUT38), .B(n671), .Z(n676) );
  NAND2_X1 U765 ( .A1(G129), .A2(n868), .ZN(n673) );
  NAND2_X1 U766 ( .A1(G117), .A2(n869), .ZN(n672) );
  NAND2_X1 U767 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U768 ( .A(KEYINPUT87), .B(n674), .Z(n675) );
  NOR2_X1 U769 ( .A1(n676), .A2(n675), .ZN(n678) );
  NAND2_X1 U770 ( .A1(n873), .A2(G141), .ZN(n677) );
  NAND2_X1 U771 ( .A1(n678), .A2(n677), .ZN(n866) );
  NAND2_X1 U772 ( .A1(G1996), .A2(n866), .ZN(n679) );
  XNOR2_X1 U773 ( .A(n679), .B(KEYINPUT88), .ZN(n688) );
  NAND2_X1 U774 ( .A1(G95), .A2(n872), .ZN(n681) );
  NAND2_X1 U775 ( .A1(G131), .A2(n873), .ZN(n680) );
  NAND2_X1 U776 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U777 ( .A(KEYINPUT86), .B(n682), .Z(n686) );
  NAND2_X1 U778 ( .A1(G119), .A2(n868), .ZN(n684) );
  NAND2_X1 U779 ( .A1(G107), .A2(n869), .ZN(n683) );
  AND2_X1 U780 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U781 ( .A1(n686), .A2(n685), .ZN(n865) );
  NAND2_X1 U782 ( .A1(G1991), .A2(n865), .ZN(n687) );
  NAND2_X1 U783 ( .A1(n688), .A2(n687), .ZN(n689) );
  XOR2_X1 U784 ( .A(KEYINPUT89), .B(n689), .Z(n929) );
  XNOR2_X1 U785 ( .A(G1986), .B(G290), .ZN(n996) );
  NOR2_X1 U786 ( .A1(n929), .A2(n996), .ZN(n690) );
  NOR2_X1 U787 ( .A1(n691), .A2(n690), .ZN(n786) );
  XNOR2_X1 U788 ( .A(G1981), .B(G305), .ZN(n1001) );
  INV_X1 U789 ( .A(n692), .ZN(n694) );
  NOR2_X1 U790 ( .A1(n720), .A2(G1961), .ZN(n695) );
  XNOR2_X1 U791 ( .A(n695), .B(KEYINPUT91), .ZN(n697) );
  XNOR2_X1 U792 ( .A(G2078), .B(KEYINPUT25), .ZN(n971) );
  NAND2_X1 U793 ( .A1(n720), .A2(n971), .ZN(n696) );
  NAND2_X1 U794 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U795 ( .A(KEYINPUT92), .B(n698), .Z(n707) );
  AND2_X1 U796 ( .A1(G301), .A2(n707), .ZN(n704) );
  NAND2_X1 U797 ( .A1(n740), .A2(G8), .ZN(n699) );
  NOR2_X1 U798 ( .A1(n779), .A2(G1966), .ZN(n753) );
  NOR2_X1 U799 ( .A1(G2084), .A2(n740), .ZN(n750) );
  NOR2_X1 U800 ( .A1(n753), .A2(n750), .ZN(n700) );
  NAND2_X1 U801 ( .A1(G8), .A2(n700), .ZN(n701) );
  XNOR2_X1 U802 ( .A(n701), .B(KEYINPUT30), .ZN(n702) );
  NOR2_X1 U803 ( .A1(G168), .A2(n702), .ZN(n703) );
  NOR2_X1 U804 ( .A1(n704), .A2(n703), .ZN(n706) );
  NOR2_X1 U805 ( .A1(G301), .A2(n707), .ZN(n708) );
  XNOR2_X1 U806 ( .A(KEYINPUT93), .B(n708), .ZN(n737) );
  NAND2_X1 U807 ( .A1(n720), .A2(G2072), .ZN(n710) );
  NAND2_X1 U808 ( .A1(G1956), .A2(n740), .ZN(n711) );
  NAND2_X1 U809 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U810 ( .A(KEYINPUT94), .B(n713), .Z(n729) );
  NAND2_X1 U811 ( .A1(n988), .A2(n729), .ZN(n728) );
  AND2_X1 U812 ( .A1(n720), .A2(G1996), .ZN(n714) );
  XOR2_X1 U813 ( .A(n714), .B(KEYINPUT26), .Z(n716) );
  NAND2_X1 U814 ( .A1(n740), .A2(G1341), .ZN(n715) );
  NAND2_X1 U815 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U816 ( .A1(n997), .A2(n717), .ZN(n718) );
  OR2_X1 U817 ( .A1(n1009), .A2(n718), .ZN(n726) );
  NAND2_X1 U818 ( .A1(n1009), .A2(n718), .ZN(n724) );
  INV_X1 U819 ( .A(G1348), .ZN(n1008) );
  NOR2_X1 U820 ( .A1(n720), .A2(n1008), .ZN(n719) );
  XNOR2_X1 U821 ( .A(n719), .B(KEYINPUT95), .ZN(n722) );
  NAND2_X1 U822 ( .A1(n720), .A2(G2067), .ZN(n721) );
  NAND2_X1 U823 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U824 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U825 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U826 ( .A1(n728), .A2(n727), .ZN(n733) );
  NOR2_X1 U827 ( .A1(n988), .A2(n729), .ZN(n731) );
  XNOR2_X1 U828 ( .A(n731), .B(n730), .ZN(n732) );
  NAND2_X1 U829 ( .A1(n733), .A2(n732), .ZN(n735) );
  XOR2_X1 U830 ( .A(KEYINPUT29), .B(KEYINPUT96), .Z(n734) );
  XNOR2_X1 U831 ( .A(n735), .B(n734), .ZN(n736) );
  NAND2_X1 U832 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U833 ( .A1(n739), .A2(n738), .ZN(n751) );
  NAND2_X1 U834 ( .A1(n751), .A2(G286), .ZN(n745) );
  NOR2_X1 U835 ( .A1(n779), .A2(G1971), .ZN(n742) );
  NOR2_X1 U836 ( .A1(G2090), .A2(n740), .ZN(n741) );
  NOR2_X1 U837 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U838 ( .A1(n743), .A2(G303), .ZN(n744) );
  NAND2_X1 U839 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U840 ( .A(KEYINPUT98), .B(n746), .ZN(n747) );
  NAND2_X1 U841 ( .A1(n747), .A2(G8), .ZN(n749) );
  XOR2_X1 U842 ( .A(KEYINPUT99), .B(KEYINPUT32), .Z(n748) );
  XNOR2_X1 U843 ( .A(n749), .B(n748), .ZN(n774) );
  NAND2_X1 U844 ( .A1(G8), .A2(n750), .ZN(n755) );
  INV_X1 U845 ( .A(n751), .ZN(n752) );
  NOR2_X1 U846 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U847 ( .A1(n755), .A2(n754), .ZN(n775) );
  NAND2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n993) );
  AND2_X1 U849 ( .A1(n775), .A2(n993), .ZN(n757) );
  INV_X1 U850 ( .A(KEYINPUT33), .ZN(n756) );
  AND2_X1 U851 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U852 ( .A1(n774), .A2(n758), .ZN(n763) );
  INV_X1 U853 ( .A(n993), .ZN(n760) );
  NOR2_X1 U854 ( .A1(G1976), .A2(G288), .ZN(n766) );
  NOR2_X1 U855 ( .A1(G1971), .A2(G303), .ZN(n759) );
  NOR2_X1 U856 ( .A1(n766), .A2(n759), .ZN(n999) );
  OR2_X1 U857 ( .A1(n760), .A2(n999), .ZN(n761) );
  OR2_X1 U858 ( .A1(KEYINPUT33), .A2(n761), .ZN(n762) );
  NAND2_X1 U859 ( .A1(n763), .A2(n762), .ZN(n765) );
  NAND2_X1 U860 ( .A1(n765), .A2(n764), .ZN(n769) );
  NAND2_X1 U861 ( .A1(n766), .A2(n764), .ZN(n767) );
  NAND2_X1 U862 ( .A1(n767), .A2(KEYINPUT33), .ZN(n768) );
  NAND2_X1 U863 ( .A1(n769), .A2(n768), .ZN(n770) );
  XOR2_X1 U864 ( .A(KEYINPUT100), .B(n770), .Z(n771) );
  NOR2_X1 U865 ( .A1(n1001), .A2(n771), .ZN(n784) );
  NOR2_X1 U866 ( .A1(G1981), .A2(G305), .ZN(n772) );
  XNOR2_X1 U867 ( .A(KEYINPUT24), .B(n772), .ZN(n773) );
  NAND2_X1 U868 ( .A1(n773), .A2(n764), .ZN(n782) );
  NAND2_X1 U869 ( .A1(n775), .A2(n774), .ZN(n778) );
  NOR2_X1 U870 ( .A1(G2090), .A2(G303), .ZN(n776) );
  NAND2_X1 U871 ( .A1(G8), .A2(n776), .ZN(n777) );
  NAND2_X1 U872 ( .A1(n778), .A2(n777), .ZN(n780) );
  NAND2_X1 U873 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n783) );
  NOR2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U876 ( .A1(n786), .A2(n785), .ZN(n798) );
  XNOR2_X1 U877 ( .A(KEYINPUT85), .B(KEYINPUT36), .ZN(n797) );
  NAND2_X1 U878 ( .A1(G128), .A2(n868), .ZN(n788) );
  NAND2_X1 U879 ( .A1(G116), .A2(n869), .ZN(n787) );
  NAND2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U881 ( .A(KEYINPUT35), .B(n789), .ZN(n795) );
  NAND2_X1 U882 ( .A1(G104), .A2(n872), .ZN(n791) );
  NAND2_X1 U883 ( .A1(G140), .A2(n873), .ZN(n790) );
  NAND2_X1 U884 ( .A1(n791), .A2(n790), .ZN(n793) );
  XOR2_X1 U885 ( .A(KEYINPUT84), .B(KEYINPUT34), .Z(n792) );
  XNOR2_X1 U886 ( .A(n793), .B(n792), .ZN(n794) );
  NAND2_X1 U887 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U888 ( .A(n797), .B(n796), .Z(n886) );
  XOR2_X1 U889 ( .A(G2067), .B(KEYINPUT37), .Z(n807) );
  AND2_X1 U890 ( .A1(n886), .A2(n807), .ZN(n910) );
  NAND2_X1 U891 ( .A1(n910), .A2(n811), .ZN(n805) );
  NAND2_X1 U892 ( .A1(n798), .A2(n805), .ZN(n814) );
  NOR2_X1 U893 ( .A1(G1996), .A2(n866), .ZN(n922) );
  NOR2_X1 U894 ( .A1(G1986), .A2(G290), .ZN(n800) );
  NOR2_X1 U895 ( .A1(G1991), .A2(n865), .ZN(n799) );
  XOR2_X1 U896 ( .A(KEYINPUT101), .B(n799), .Z(n909) );
  NOR2_X1 U897 ( .A1(n800), .A2(n909), .ZN(n801) );
  XNOR2_X1 U898 ( .A(n801), .B(KEYINPUT102), .ZN(n802) );
  NOR2_X1 U899 ( .A1(n929), .A2(n802), .ZN(n803) );
  NOR2_X1 U900 ( .A1(n922), .A2(n803), .ZN(n804) );
  XNOR2_X1 U901 ( .A(KEYINPUT39), .B(n804), .ZN(n806) );
  NAND2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n809) );
  NOR2_X1 U903 ( .A1(n807), .A2(n886), .ZN(n808) );
  XNOR2_X1 U904 ( .A(n808), .B(KEYINPUT103), .ZN(n930) );
  NAND2_X1 U905 ( .A1(n809), .A2(n930), .ZN(n810) );
  NAND2_X1 U906 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U907 ( .A(n812), .B(KEYINPUT104), .ZN(n813) );
  NAND2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U909 ( .A(n815), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n816), .ZN(G217) );
  AND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n817) );
  NAND2_X1 U912 ( .A1(G661), .A2(n817), .ZN(G259) );
  NAND2_X1 U913 ( .A1(G3), .A2(G1), .ZN(n818) );
  NAND2_X1 U914 ( .A1(n819), .A2(n818), .ZN(G188) );
  INV_X1 U916 ( .A(G120), .ZN(G236) );
  INV_X1 U917 ( .A(G96), .ZN(G221) );
  INV_X1 U918 ( .A(G69), .ZN(G235) );
  NOR2_X1 U919 ( .A1(n821), .A2(n820), .ZN(G325) );
  INV_X1 U920 ( .A(G325), .ZN(G261) );
  XOR2_X1 U921 ( .A(KEYINPUT106), .B(n822), .Z(G319) );
  XNOR2_X1 U922 ( .A(G2067), .B(G2084), .ZN(n823) );
  XNOR2_X1 U923 ( .A(n823), .B(KEYINPUT42), .ZN(n833) );
  XOR2_X1 U924 ( .A(G2678), .B(KEYINPUT43), .Z(n825) );
  XNOR2_X1 U925 ( .A(KEYINPUT108), .B(G2096), .ZN(n824) );
  XNOR2_X1 U926 ( .A(n825), .B(n824), .ZN(n829) );
  XOR2_X1 U927 ( .A(G2100), .B(G2090), .Z(n827) );
  XNOR2_X1 U928 ( .A(G2072), .B(G2078), .ZN(n826) );
  XNOR2_X1 U929 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U930 ( .A(n829), .B(n828), .Z(n831) );
  XNOR2_X1 U931 ( .A(KEYINPUT109), .B(KEYINPUT107), .ZN(n830) );
  XNOR2_X1 U932 ( .A(n831), .B(n830), .ZN(n832) );
  XNOR2_X1 U933 ( .A(n833), .B(n832), .ZN(G227) );
  XOR2_X1 U934 ( .A(G1976), .B(G1956), .Z(n835) );
  XNOR2_X1 U935 ( .A(G1981), .B(G1966), .ZN(n834) );
  XNOR2_X1 U936 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U937 ( .A(n836), .B(KEYINPUT41), .Z(n838) );
  XNOR2_X1 U938 ( .A(G1996), .B(G1991), .ZN(n837) );
  XNOR2_X1 U939 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U940 ( .A(G2474), .B(G1986), .Z(n840) );
  XNOR2_X1 U941 ( .A(G1961), .B(G1971), .ZN(n839) );
  XNOR2_X1 U942 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(G229) );
  NAND2_X1 U944 ( .A1(G124), .A2(n868), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n843), .B(KEYINPUT44), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n844), .B(KEYINPUT110), .ZN(n846) );
  NAND2_X1 U947 ( .A1(G112), .A2(n869), .ZN(n845) );
  NAND2_X1 U948 ( .A1(n846), .A2(n845), .ZN(n850) );
  NAND2_X1 U949 ( .A1(G100), .A2(n872), .ZN(n848) );
  NAND2_X1 U950 ( .A1(n873), .A2(G136), .ZN(n847) );
  NAND2_X1 U951 ( .A1(n848), .A2(n847), .ZN(n849) );
  NOR2_X1 U952 ( .A1(n850), .A2(n849), .ZN(G162) );
  XOR2_X1 U953 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n852) );
  XNOR2_X1 U954 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n851) );
  XNOR2_X1 U955 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U956 ( .A(n853), .B(KEYINPUT114), .Z(n863) );
  NAND2_X1 U957 ( .A1(G103), .A2(n872), .ZN(n855) );
  NAND2_X1 U958 ( .A1(G139), .A2(n873), .ZN(n854) );
  NAND2_X1 U959 ( .A1(n855), .A2(n854), .ZN(n861) );
  NAND2_X1 U960 ( .A1(G127), .A2(n868), .ZN(n857) );
  NAND2_X1 U961 ( .A1(G115), .A2(n869), .ZN(n856) );
  NAND2_X1 U962 ( .A1(n857), .A2(n856), .ZN(n858) );
  XOR2_X1 U963 ( .A(KEYINPUT112), .B(n858), .Z(n859) );
  XNOR2_X1 U964 ( .A(KEYINPUT47), .B(n859), .ZN(n860) );
  NOR2_X1 U965 ( .A1(n861), .A2(n860), .ZN(n911) );
  XNOR2_X1 U966 ( .A(n911), .B(KEYINPUT113), .ZN(n862) );
  XNOR2_X1 U967 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U968 ( .A(G164), .B(n864), .ZN(n885) );
  XNOR2_X1 U969 ( .A(n918), .B(n865), .ZN(n867) );
  XNOR2_X1 U970 ( .A(n867), .B(n866), .ZN(n881) );
  NAND2_X1 U971 ( .A1(G130), .A2(n868), .ZN(n871) );
  NAND2_X1 U972 ( .A1(G118), .A2(n869), .ZN(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n879) );
  NAND2_X1 U974 ( .A1(G106), .A2(n872), .ZN(n875) );
  NAND2_X1 U975 ( .A1(G142), .A2(n873), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U977 ( .A(KEYINPUT111), .B(n876), .ZN(n877) );
  XNOR2_X1 U978 ( .A(KEYINPUT45), .B(n877), .ZN(n878) );
  NOR2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U980 ( .A(n881), .B(n880), .Z(n883) );
  XNOR2_X1 U981 ( .A(G160), .B(G162), .ZN(n882) );
  XNOR2_X1 U982 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U983 ( .A(n885), .B(n884), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n887), .B(n886), .ZN(n888) );
  NOR2_X1 U985 ( .A1(G37), .A2(n888), .ZN(G395) );
  XNOR2_X1 U986 ( .A(n1009), .B(G171), .ZN(n889) );
  XNOR2_X1 U987 ( .A(n889), .B(G286), .ZN(n891) );
  XNOR2_X1 U988 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U989 ( .A1(G37), .A2(n892), .ZN(G397) );
  XOR2_X1 U990 ( .A(G2430), .B(G2451), .Z(n894) );
  XNOR2_X1 U991 ( .A(G2446), .B(G2427), .ZN(n893) );
  XNOR2_X1 U992 ( .A(n894), .B(n893), .ZN(n901) );
  XOR2_X1 U993 ( .A(G2438), .B(G2435), .Z(n896) );
  XNOR2_X1 U994 ( .A(G2443), .B(KEYINPUT105), .ZN(n895) );
  XNOR2_X1 U995 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U996 ( .A(n897), .B(G2454), .Z(n899) );
  XNOR2_X1 U997 ( .A(G1348), .B(G1341), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n902) );
  NAND2_X1 U1000 ( .A1(n902), .A2(G14), .ZN(n908) );
  NAND2_X1 U1001 ( .A1(n908), .A2(G319), .ZN(n905) );
  NOR2_X1 U1002 ( .A1(G227), .A2(G229), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(KEYINPUT49), .B(n903), .ZN(n904) );
  NOR2_X1 U1004 ( .A1(n905), .A2(n904), .ZN(n907) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n906) );
  NAND2_X1 U1006 ( .A1(n907), .A2(n906), .ZN(G225) );
  INV_X1 U1007 ( .A(G225), .ZN(G308) );
  INV_X1 U1008 ( .A(G108), .ZN(G238) );
  INV_X1 U1009 ( .A(n908), .ZN(G401) );
  XNOR2_X1 U1010 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n978) );
  NOR2_X1 U1011 ( .A1(n910), .A2(n909), .ZN(n927) );
  XOR2_X1 U1012 ( .A(G2072), .B(n911), .Z(n913) );
  XOR2_X1 U1013 ( .A(G164), .B(G2078), .Z(n912) );
  NOR2_X1 U1014 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1015 ( .A(KEYINPUT118), .B(n914), .ZN(n915) );
  XNOR2_X1 U1016 ( .A(n915), .B(KEYINPUT50), .ZN(n920) );
  XNOR2_X1 U1017 ( .A(G2084), .B(G160), .ZN(n916) );
  XNOR2_X1 U1018 ( .A(KEYINPUT117), .B(n916), .ZN(n917) );
  NOR2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n925) );
  XOR2_X1 U1021 ( .A(G2090), .B(G162), .Z(n921) );
  NOR2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(n923), .B(KEYINPUT51), .ZN(n924) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n931) );
  NAND2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1028 ( .A(KEYINPUT52), .B(n932), .Z(n933) );
  NAND2_X1 U1029 ( .A1(n978), .A2(n933), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n934), .A2(G29), .ZN(n987) );
  XNOR2_X1 U1031 ( .A(G1348), .B(KEYINPUT59), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(n935), .B(G4), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(G1981), .B(G6), .ZN(n937) );
  XNOR2_X1 U1034 ( .A(G1341), .B(G19), .ZN(n936) );
  NOR2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n942) );
  XOR2_X1 U1037 ( .A(KEYINPUT125), .B(G1956), .Z(n940) );
  XNOR2_X1 U1038 ( .A(G20), .B(n940), .ZN(n941) );
  NOR2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1040 ( .A(KEYINPUT60), .B(n943), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(n944), .B(KEYINPUT126), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(G1966), .B(G21), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(G5), .B(G1961), .ZN(n945) );
  NOR2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n956) );
  XOR2_X1 U1046 ( .A(G1976), .B(G23), .Z(n952) );
  XNOR2_X1 U1047 ( .A(G1971), .B(G22), .ZN(n950) );
  XNOR2_X1 U1048 ( .A(G24), .B(G1986), .ZN(n949) );
  NOR2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1050 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1051 ( .A(KEYINPUT58), .B(n953), .Z(n954) );
  XNOR2_X1 U1052 ( .A(KEYINPUT127), .B(n954), .ZN(n955) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  XOR2_X1 U1054 ( .A(KEYINPUT61), .B(n957), .Z(n958) );
  NOR2_X1 U1055 ( .A1(G16), .A2(n958), .ZN(n985) );
  XOR2_X1 U1056 ( .A(G2090), .B(G35), .Z(n961) );
  XOR2_X1 U1057 ( .A(KEYINPUT54), .B(G34), .Z(n959) );
  XNOR2_X1 U1058 ( .A(n959), .B(G2084), .ZN(n960) );
  NAND2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n977) );
  XNOR2_X1 U1060 ( .A(KEYINPUT121), .B(G1996), .ZN(n962) );
  XNOR2_X1 U1061 ( .A(n962), .B(G32), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(G2067), .B(G26), .ZN(n964) );
  XNOR2_X1 U1063 ( .A(G33), .B(G2072), .ZN(n963) );
  NOR2_X1 U1064 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1065 ( .A1(G28), .A2(n965), .ZN(n968) );
  XNOR2_X1 U1066 ( .A(G25), .B(G1991), .ZN(n966) );
  XNOR2_X1 U1067 ( .A(KEYINPUT120), .B(n966), .ZN(n967) );
  NOR2_X1 U1068 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1069 ( .A1(n970), .A2(n969), .ZN(n973) );
  XOR2_X1 U1070 ( .A(G27), .B(n971), .Z(n972) );
  NOR2_X1 U1071 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1072 ( .A(KEYINPUT53), .B(n974), .ZN(n975) );
  XNOR2_X1 U1073 ( .A(KEYINPUT122), .B(n975), .ZN(n976) );
  NOR2_X1 U1074 ( .A1(n977), .A2(n976), .ZN(n980) );
  XNOR2_X1 U1075 ( .A(KEYINPUT123), .B(n978), .ZN(n979) );
  XNOR2_X1 U1076 ( .A(n980), .B(n979), .ZN(n982) );
  INV_X1 U1077 ( .A(G29), .ZN(n981) );
  NAND2_X1 U1078 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1079 ( .A1(n983), .A2(G11), .ZN(n984) );
  NOR2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n1015) );
  XNOR2_X1 U1082 ( .A(n988), .B(G1956), .ZN(n990) );
  NAND2_X1 U1083 ( .A1(G1971), .A2(G303), .ZN(n989) );
  NAND2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n992) );
  XNOR2_X1 U1085 ( .A(G1961), .B(G301), .ZN(n991) );
  NOR2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n994) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n1007) );
  XOR2_X1 U1089 ( .A(G1341), .B(n997), .Z(n998) );
  NAND2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1005) );
  XOR2_X1 U1091 ( .A(G1966), .B(G168), .Z(n1000) );
  XNOR2_X1 U1092 ( .A(KEYINPUT124), .B(n1000), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1094 ( .A(KEYINPUT57), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(n1009), .B(n1008), .ZN(n1010) );
  NOR2_X1 U1098 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XOR2_X1 U1099 ( .A(G16), .B(KEYINPUT56), .Z(n1012) );
  NOR2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1102 ( .A(n1016), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1103 ( .A(G311), .ZN(G150) );
endmodule

