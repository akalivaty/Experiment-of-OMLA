//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT79), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n190), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n196));
  OR2_X1    g010(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT67), .A2(KEYINPUT1), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n193), .A2(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n191), .A2(G146), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n200), .A2(new_n201), .A3(G128), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n195), .B(new_n196), .C1(new_n199), .C2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G107), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT78), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT78), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G107), .ZN(new_n208));
  AOI21_X1  g022(.A(G104), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(G104), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(G101), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n213), .B1(G104), .B2(new_n205), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G104), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(KEYINPUT3), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(new_n206), .A3(new_n208), .ZN(new_n218));
  AOI21_X1  g032(.A(G101), .B1(new_n216), .B2(G107), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n215), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n212), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n189), .B1(new_n204), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT78), .B(G107), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n210), .B1(new_n223), .B2(G104), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n214), .B1(new_n223), .B2(new_n217), .ZN(new_n225));
  AOI22_X1  g039(.A1(G101), .A2(new_n224), .B1(new_n225), .B2(new_n219), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(KEYINPUT79), .A3(new_n203), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT10), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT0), .B(G128), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n192), .B2(new_n194), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n200), .A2(new_n201), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n216), .A2(G107), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n215), .A2(new_n218), .A3(new_n234), .ZN(new_n235));
  AOI22_X1  g049(.A1(KEYINPUT4), .A2(new_n220), .B1(new_n235), .B2(G101), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n235), .A2(KEYINPUT4), .A3(G101), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n233), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G143), .B(G146), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n239), .A2(G128), .A3(new_n197), .A4(new_n198), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n199), .A2(new_n191), .A3(G146), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n240), .A2(new_n241), .A3(new_n195), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n226), .A2(KEYINPUT10), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n228), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G131), .ZN(new_n246));
  INV_X1    g060(.A(G137), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(G134), .ZN(new_n248));
  INV_X1    g062(.A(G134), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT65), .B1(new_n249), .B2(G137), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n248), .B1(new_n250), .B2(KEYINPUT11), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT11), .ZN(new_n252));
  OAI211_X1 g066(.A(KEYINPUT65), .B(new_n252), .C1(new_n249), .C2(G137), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n246), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT66), .B(G131), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n251), .A2(new_n256), .A3(new_n253), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n245), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(G110), .B(G140), .ZN(new_n261));
  INV_X1    g075(.A(G953), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n262), .A2(G227), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n261), .B(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT12), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n242), .B1(new_n220), .B2(new_n212), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n268), .B1(new_n222), .B2(new_n227), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT80), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n258), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n221), .A2(new_n241), .A3(new_n195), .A4(new_n240), .ZN(new_n272));
  AOI21_X1  g086(.A(KEYINPUT79), .B1(new_n226), .B2(new_n203), .ZN(new_n273));
  AND4_X1   g087(.A1(KEYINPUT79), .A2(new_n203), .A3(new_n220), .A4(new_n212), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n270), .B(new_n272), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n267), .B1(new_n271), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT81), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT81), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n279), .B(new_n267), .C1(new_n271), .C2(new_n276), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n269), .A2(new_n267), .A3(new_n259), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n266), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n245), .A2(new_n259), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n265), .B1(new_n286), .B2(new_n260), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n187), .B(new_n188), .C1(new_n284), .C2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n187), .A2(new_n188), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n282), .B1(new_n278), .B2(new_n280), .ZN(new_n291));
  INV_X1    g105(.A(new_n260), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n264), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n266), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n286), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n288), .B(new_n290), .C1(new_n296), .C2(new_n187), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT9), .B(G234), .ZN(new_n298));
  OAI21_X1  g112(.A(G221), .B1(new_n298), .B2(G902), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(G116), .B(G122), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT14), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G122), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(G116), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n205), .B1(new_n305), .B2(KEYINPUT14), .ZN(new_n306));
  AOI22_X1  g120(.A1(new_n303), .A2(new_n306), .B1(new_n223), .B2(new_n301), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n190), .A2(G143), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(KEYINPUT91), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n190), .A2(G143), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n249), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n249), .B1(new_n309), .B2(new_n310), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n307), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT92), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n309), .A2(KEYINPUT92), .A3(new_n249), .A4(new_n310), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n223), .B(new_n301), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT13), .ZN(new_n320));
  OR2_X1    g134(.A1(new_n309), .A2(new_n320), .ZN(new_n321));
  AOI22_X1  g135(.A1(new_n309), .A2(new_n320), .B1(new_n190), .B2(G143), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n249), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n314), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G217), .ZN(new_n325));
  NOR3_X1   g139(.A1(new_n298), .A2(new_n325), .A3(G953), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(KEYINPUT93), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT94), .ZN(new_n329));
  INV_X1    g143(.A(new_n327), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n314), .B(new_n330), .C1(new_n319), .C2(new_n323), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n328), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  OR3_X1    g146(.A1(new_n324), .A2(new_n329), .A3(new_n327), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n333), .A3(new_n188), .ZN(new_n334));
  INV_X1    g148(.A(G478), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n335), .A2(KEYINPUT15), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n334), .B(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT20), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT90), .ZN(new_n339));
  XNOR2_X1  g153(.A(G125), .B(G140), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT74), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G140), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G125), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT74), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n342), .A2(KEYINPUT16), .A3(new_n346), .ZN(new_n347));
  OR2_X1    g161(.A1(new_n345), .A2(KEYINPUT16), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n193), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n193), .B1(new_n347), .B2(new_n348), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n339), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n347), .A2(new_n348), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G146), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(KEYINPUT90), .A3(new_n349), .ZN(new_n355));
  INV_X1    g169(.A(G237), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(new_n262), .A3(G214), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(KEYINPUT88), .A3(new_n191), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n191), .A2(KEYINPUT88), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n359), .A2(G214), .A3(new_n356), .A4(new_n262), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(new_n256), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT17), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n256), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n361), .A2(KEYINPUT17), .A3(new_n365), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n352), .A2(new_n355), .A3(new_n364), .A4(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(G113), .B(G122), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(new_n216), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT89), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n370), .A2(KEYINPUT18), .A3(G131), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n361), .B(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n340), .A2(new_n193), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n342), .A2(new_n346), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n373), .B1(new_n374), .B2(new_n193), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n367), .A2(new_n369), .A3(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n361), .B(new_n365), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n354), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n340), .A2(KEYINPUT19), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(new_n374), .B2(KEYINPUT19), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(G146), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n376), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n369), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n377), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(G475), .A2(G902), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n338), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n387), .ZN(new_n389));
  AOI211_X1 g203(.A(KEYINPUT20), .B(new_n389), .C1(new_n377), .C2(new_n385), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n367), .A2(new_n376), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n384), .ZN(new_n392));
  AOI21_X1  g206(.A(G902), .B1(new_n392), .B2(new_n377), .ZN(new_n393));
  INV_X1    g207(.A(G475), .ZN(new_n394));
  OAI22_X1  g208(.A1(new_n388), .A2(new_n390), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n337), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(G234), .A2(G237), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n397), .A2(G952), .A3(new_n262), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n397), .A2(G902), .A3(G953), .ZN(new_n399));
  XNOR2_X1  g213(.A(KEYINPUT21), .B(G898), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n396), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n300), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(G214), .B1(G237), .B2(G902), .ZN(new_n405));
  OAI21_X1  g219(.A(G210), .B1(G237), .B2(G902), .ZN(new_n406));
  XNOR2_X1  g220(.A(G116), .B(G119), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT2), .B(G113), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT69), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XOR2_X1   g224(.A(KEYINPUT2), .B(G113), .Z(new_n411));
  INV_X1    g225(.A(KEYINPUT69), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n412), .A3(new_n407), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n411), .A2(KEYINPUT68), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT68), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n409), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n415), .A2(new_n408), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n419), .B1(new_n236), .B2(new_n237), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n407), .A2(KEYINPUT5), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT5), .ZN(new_n422));
  INV_X1    g236(.A(G119), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(G116), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n424), .A2(G113), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n226), .A2(new_n414), .A3(new_n426), .ZN(new_n427));
  XNOR2_X1  g241(.A(G110), .B(G122), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n420), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT6), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n428), .B(KEYINPUT82), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n432), .B1(new_n420), .B2(new_n427), .ZN(new_n433));
  OAI21_X1  g247(.A(KEYINPUT83), .B1(new_n430), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(G125), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n242), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n233), .A2(G125), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n262), .A2(G224), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n438), .B(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT6), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n433), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n235), .A2(G101), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n220), .A2(KEYINPUT4), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n235), .A2(KEYINPUT4), .A3(G101), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n445), .A2(new_n446), .B1(new_n414), .B2(new_n418), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n226), .A2(new_n414), .A3(new_n426), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n431), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT83), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n449), .A2(new_n429), .A3(new_n450), .A4(KEYINPUT6), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n434), .A2(new_n440), .A3(new_n442), .A4(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT84), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n451), .A2(new_n442), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n455), .A2(KEYINPUT84), .A3(new_n440), .A4(new_n434), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n439), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n440), .B1(KEYINPUT7), .B2(new_n458), .ZN(new_n459));
  XOR2_X1   g273(.A(new_n425), .B(KEYINPUT86), .Z(new_n460));
  XNOR2_X1  g274(.A(new_n421), .B(KEYINPUT85), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n414), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n226), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n428), .B(KEYINPUT8), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n414), .A2(new_n426), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n463), .B(new_n464), .C1(new_n226), .C2(new_n465), .ZN(new_n466));
  OR3_X1    g280(.A1(new_n438), .A2(KEYINPUT7), .A3(new_n458), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n459), .A2(new_n466), .A3(new_n429), .A4(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n188), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n406), .B1(new_n457), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n406), .ZN(new_n472));
  AOI211_X1 g286(.A(new_n472), .B(new_n469), .C1(new_n454), .C2(new_n456), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n405), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT87), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(KEYINPUT87), .B(new_n405), .C1(new_n471), .C2(new_n473), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G472), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n188), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n251), .A2(new_n256), .A3(new_n253), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n233), .B1(new_n481), .B2(new_n254), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n249), .A2(G137), .ZN(new_n483));
  OAI21_X1  g297(.A(G131), .B1(new_n483), .B2(new_n248), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n242), .A2(new_n257), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n482), .A2(new_n485), .A3(KEYINPUT30), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT64), .ZN(new_n487));
  XOR2_X1   g301(.A(KEYINPUT0), .B(G128), .Z(new_n488));
  OAI211_X1 g302(.A(new_n487), .B(new_n232), .C1(new_n488), .C2(new_n239), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n487), .B1(new_n230), .B2(new_n232), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n257), .A2(new_n484), .ZN(new_n493));
  AOI22_X1  g307(.A1(new_n492), .A2(new_n258), .B1(new_n493), .B2(new_n242), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n419), .B(new_n486), .C1(new_n494), .C2(KEYINPUT30), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n407), .B1(new_n411), .B2(KEYINPUT68), .ZN(new_n496));
  AOI22_X1  g310(.A1(new_n410), .A2(new_n413), .B1(new_n496), .B2(new_n417), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n482), .A2(new_n485), .A3(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n499));
  INV_X1    g313(.A(G210), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n500), .A2(G237), .A3(G953), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n499), .B(new_n501), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT26), .B(G101), .Z(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT71), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT71), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n498), .A2(new_n507), .A3(new_n504), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n495), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT31), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n495), .A2(new_n506), .A3(KEYINPUT31), .A4(new_n508), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OR2_X1    g327(.A1(new_n494), .A2(new_n497), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n498), .A2(KEYINPUT28), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT28), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n482), .A2(new_n485), .A3(new_n497), .A4(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n504), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n480), .B1(new_n513), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT32), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n482), .A2(new_n485), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n419), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n518), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n504), .A2(KEYINPUT29), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n188), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n495), .A2(new_n498), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT29), .B1(new_n529), .B2(new_n520), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n514), .A2(new_n518), .A3(new_n504), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(KEYINPUT72), .B1(new_n532), .B2(new_n479), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT32), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n511), .A2(new_n512), .B1(new_n519), .B2(new_n520), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n534), .B1(new_n535), .B2(new_n480), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT72), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n514), .A2(new_n518), .A3(new_n504), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n504), .B1(new_n495), .B2(new_n498), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n538), .A2(new_n539), .A3(KEYINPUT29), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n537), .B(G472), .C1(new_n540), .C2(new_n528), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n523), .A2(new_n533), .A3(new_n536), .A4(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n262), .A2(G221), .A3(G234), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT75), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT22), .B(G137), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT24), .B(G110), .ZN(new_n547));
  OR3_X1    g361(.A1(new_n423), .A2(KEYINPUT73), .A3(G128), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT73), .B1(new_n423), .B2(G128), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n423), .A2(G128), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT23), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(new_n423), .B2(G128), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n190), .A2(KEYINPUT23), .A3(G119), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n553), .A2(new_n550), .A3(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(G110), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n547), .A2(new_n551), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(new_n193), .B2(new_n340), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n354), .ZN(new_n559));
  OR2_X1    g373(.A1(new_n551), .A2(new_n547), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n555), .A2(new_n556), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n560), .B(new_n561), .C1(new_n350), .C2(new_n351), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT76), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n559), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n563), .B1(new_n559), .B2(new_n562), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n546), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n546), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n559), .A2(new_n562), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n567), .B1(new_n568), .B2(KEYINPUT76), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n325), .B1(G234), .B2(new_n188), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(G902), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT77), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n566), .A2(new_n188), .A3(new_n569), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT25), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT25), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n566), .A2(new_n578), .A3(new_n188), .A4(new_n569), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n577), .A2(new_n579), .A3(new_n571), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n570), .A2(KEYINPUT77), .A3(new_n572), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n575), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n542), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n404), .A2(new_n478), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(new_n585), .B(G101), .ZN(G3));
  OR2_X1    g400(.A1(new_n535), .A2(G902), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n522), .B1(new_n587), .B2(G472), .ZN(new_n588));
  AND4_X1   g402(.A1(new_n582), .A2(new_n297), .A3(new_n299), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n457), .A2(new_n470), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n472), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n457), .A2(new_n406), .A3(new_n470), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(new_n405), .A3(new_n402), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT33), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n332), .A2(new_n333), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n328), .A2(KEYINPUT33), .A3(new_n331), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n335), .A2(G902), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n334), .A2(new_n335), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n395), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(new_n602), .B(KEYINPUT95), .Z(new_n603));
  NOR2_X1   g417(.A1(new_n594), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n589), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(KEYINPUT96), .ZN(new_n606));
  XOR2_X1   g420(.A(KEYINPUT34), .B(G104), .Z(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G6));
  INV_X1    g422(.A(new_n405), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n591), .B2(new_n592), .ZN(new_n610));
  INV_X1    g424(.A(new_n336), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n334), .B(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n612), .A2(new_n395), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n589), .A2(new_n610), .A3(new_n402), .A4(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT35), .B(G107), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G9));
  NOR2_X1   g430(.A1(new_n567), .A2(KEYINPUT36), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n568), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n572), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n580), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n588), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT97), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n404), .A2(new_n478), .A3(new_n622), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT37), .B(G110), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT98), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n623), .B(new_n625), .ZN(G12));
  INV_X1    g440(.A(G900), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n399), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n398), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AND4_X1   g444(.A1(new_n542), .A2(new_n613), .A3(new_n620), .A4(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n631), .A2(new_n610), .A3(new_n299), .A4(new_n297), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT99), .B(G128), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G30));
  NAND2_X1  g448(.A1(new_n525), .A2(new_n498), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n520), .ZN(new_n636));
  AOI21_X1  g450(.A(G902), .B1(new_n509), .B2(new_n636), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n523), .B(new_n536), .C1(new_n479), .C2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n620), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n337), .A2(new_n395), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n640), .A2(new_n609), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n593), .A2(KEYINPUT38), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n471), .A2(new_n473), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT38), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n643), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n647), .B1(new_n643), .B2(new_n646), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n642), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n630), .B(KEYINPUT39), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n297), .A2(new_n299), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT40), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n297), .A2(new_n654), .A3(new_n299), .A4(new_n651), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(new_n191), .ZN(G45));
  NAND2_X1  g472(.A1(new_n542), .A2(new_n620), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n395), .A2(new_n601), .A3(new_n630), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n661), .A2(new_n610), .A3(new_n299), .A4(new_n297), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G146), .ZN(G48));
  INV_X1    g477(.A(new_n280), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(KEYINPUT80), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n258), .A3(new_n275), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n279), .B1(new_n667), .B2(new_n267), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n283), .B1(new_n664), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n287), .B1(new_n669), .B2(new_n294), .ZN(new_n670));
  OAI21_X1  g484(.A(G469), .B1(new_n670), .B2(G902), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n299), .A3(new_n288), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT102), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n671), .A2(KEYINPUT102), .A3(new_n288), .A4(new_n299), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(KEYINPUT103), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n674), .A2(new_n678), .A3(new_n675), .ZN(new_n679));
  AND2_X1   g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n594), .A2(new_n603), .A3(new_n583), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT41), .B(G113), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G15));
  INV_X1    g498(.A(new_n613), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n594), .A2(new_n583), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G116), .ZN(G18));
  AND3_X1   g502(.A1(new_n674), .A2(new_n610), .A3(new_n675), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n659), .A2(new_n403), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G119), .ZN(G21));
  AOI22_X1  g506(.A1(new_n511), .A2(new_n512), .B1(new_n520), .B2(new_n526), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n693), .A2(new_n480), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT104), .B(G472), .Z(new_n695));
  NAND2_X1  g509(.A1(new_n587), .A2(new_n695), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n582), .A2(new_n694), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n402), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n699));
  INV_X1    g513(.A(new_n388), .ZN(new_n700));
  INV_X1    g514(.A(new_n390), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n392), .A2(new_n377), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n188), .ZN(new_n703));
  AOI22_X1  g517(.A1(new_n700), .A2(new_n701), .B1(new_n703), .B2(G475), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n699), .B1(new_n704), .B2(new_n612), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n337), .A2(new_n395), .A3(KEYINPUT105), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n708), .A2(new_n610), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g524(.A(KEYINPUT106), .B1(new_n474), .B2(new_n707), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n698), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n677), .A3(new_n679), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G122), .ZN(G24));
  NAND3_X1  g528(.A1(new_n696), .A2(new_n620), .A3(new_n694), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n715), .A2(new_n660), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n674), .A2(new_n610), .A3(new_n675), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G125), .ZN(G27));
  NAND2_X1  g532(.A1(new_n669), .A2(new_n294), .ZN(new_n719));
  INV_X1    g533(.A(new_n287), .ZN(new_n720));
  AOI21_X1  g534(.A(G902), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n289), .B1(new_n721), .B2(new_n187), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n293), .A2(KEYINPUT107), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n724), .B(new_n264), .C1(new_n291), .C2(new_n292), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n723), .A2(G469), .A3(new_n295), .A4(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n299), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n609), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n591), .A2(new_n592), .A3(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n575), .A2(new_n580), .A3(new_n581), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT108), .B1(new_n522), .B2(KEYINPUT32), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n735));
  NOR4_X1   g549(.A1(new_n535), .A2(new_n735), .A3(new_n534), .A4(new_n480), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n533), .A2(new_n536), .A3(new_n541), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n733), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n660), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(KEYINPUT42), .B1(new_n732), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n730), .B1(new_n722), .B2(new_n726), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n660), .A2(KEYINPUT42), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(new_n584), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n742), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n246), .ZN(G33));
  INV_X1    g561(.A(new_n630), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n685), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n727), .A2(new_n731), .A3(new_n584), .A4(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G134), .ZN(G36));
  AOI21_X1  g565(.A(new_n395), .B1(new_n600), .B2(new_n599), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n752), .B(KEYINPUT43), .Z(new_n753));
  NOR3_X1   g567(.A1(new_n753), .A2(new_n588), .A3(new_n639), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(KEYINPUT44), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n471), .A2(new_n473), .A3(new_n609), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n288), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n187), .B1(new_n296), .B2(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n723), .A2(KEYINPUT45), .A3(new_n295), .A4(new_n725), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n761), .A2(new_n762), .A3(KEYINPUT109), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT109), .B1(new_n761), .B2(new_n762), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n290), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n759), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  OAI211_X1 g581(.A(KEYINPUT46), .B(new_n290), .C1(new_n763), .C2(new_n764), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n728), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n769), .A2(KEYINPUT110), .A3(new_n651), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT110), .B1(new_n769), .B2(new_n651), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n758), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G137), .ZN(G39));
  NOR4_X1   g587(.A1(new_n757), .A2(new_n542), .A3(new_n582), .A4(new_n660), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n769), .A2(KEYINPUT47), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n769), .A2(KEYINPUT47), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  XOR2_X1   g591(.A(KEYINPUT111), .B(G140), .Z(new_n778));
  XNOR2_X1  g592(.A(new_n777), .B(new_n778), .ZN(G42));
  OR2_X1    g593(.A1(new_n648), .A2(new_n649), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n582), .A2(new_n729), .A3(new_n752), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n671), .A2(new_n288), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n781), .B1(new_n782), .B2(KEYINPUT49), .ZN(new_n783));
  XOR2_X1   g597(.A(new_n783), .B(KEYINPUT112), .Z(new_n784));
  NOR2_X1   g598(.A1(new_n782), .A2(KEYINPUT49), .ZN(new_n785));
  OR4_X1    g599(.A1(new_n780), .A2(new_n784), .A3(new_n638), .A4(new_n785), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n677), .B(new_n679), .C1(new_n681), .C2(new_n686), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n401), .B1(new_n685), .B2(new_n602), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n476), .A2(new_n477), .A3(new_n788), .ZN(new_n789));
  AOI22_X1  g603(.A1(new_n689), .A2(new_n690), .B1(new_n789), .B2(new_n589), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n404), .B(new_n478), .C1(new_n622), .C2(new_n584), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n787), .A2(new_n790), .A3(new_n713), .A4(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n727), .A2(new_n716), .A3(new_n731), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT113), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n743), .A2(new_n795), .A3(new_n716), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  AND4_X1   g611(.A1(new_n542), .A2(new_n396), .A3(new_n620), .A4(new_n630), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(new_n299), .A3(new_n297), .A4(new_n756), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n750), .A2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n797), .A2(new_n800), .A3(new_n742), .A4(new_n745), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n792), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(KEYINPUT114), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n717), .A2(new_n662), .A3(new_n632), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n748), .A2(new_n728), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n638), .A2(new_n639), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n727), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n710), .B2(new_n711), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n804), .B1(new_n805), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n709), .B1(new_n708), .B2(new_n610), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n474), .A2(new_n707), .A3(KEYINPUT106), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n727), .B(new_n807), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n300), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n814), .B(new_n610), .C1(new_n631), .C2(new_n661), .ZN(new_n815));
  XNOR2_X1  g629(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n813), .A2(new_n815), .A3(new_n717), .A4(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n810), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT53), .B1(new_n802), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT115), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n803), .B1(new_n805), .B2(new_n809), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n813), .A2(new_n815), .A3(KEYINPUT52), .A4(new_n717), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n802), .A2(KEYINPUT53), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n819), .A2(KEYINPUT115), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT54), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n582), .A2(new_n694), .A3(new_n696), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n753), .A2(new_n629), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(new_n757), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n769), .B(KEYINPUT47), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n782), .A2(new_n299), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n676), .A2(new_n757), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n638), .A2(new_n733), .A3(new_n629), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n839), .A2(new_n395), .A3(new_n601), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n753), .A2(new_n629), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n842), .A2(new_n715), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n830), .A2(new_n609), .A3(new_n674), .A4(new_n675), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n845), .B1(new_n846), .B2(new_n780), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT50), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n845), .B(KEYINPUT50), .C1(new_n846), .C2(new_n780), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n849), .A2(KEYINPUT117), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT117), .B1(new_n849), .B2(new_n850), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n844), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n828), .B1(new_n836), .B2(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n787), .A2(new_n713), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n790), .A2(new_n791), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n742), .A2(new_n745), .A3(new_n750), .A4(new_n799), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n794), .A2(new_n796), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n823), .A2(new_n855), .A3(new_n856), .A4(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n802), .A2(KEYINPUT53), .A3(new_n818), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  AND4_X1   g679(.A1(KEYINPUT51), .A2(new_n844), .A3(new_n849), .A4(new_n850), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n839), .A2(new_n603), .ZN(new_n867));
  INV_X1    g681(.A(G952), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n830), .A2(new_n689), .ZN(new_n869));
  NOR4_X1   g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .A4(G953), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n837), .A2(new_n739), .A3(new_n841), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT48), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT118), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT118), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n870), .A2(new_n875), .A3(new_n872), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n835), .A2(new_n866), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  AND4_X1   g691(.A1(new_n827), .A2(new_n854), .A3(new_n865), .A4(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(G952), .A2(G953), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n786), .B1(new_n878), .B2(new_n879), .ZN(G75));
  NAND2_X1  g694(.A1(new_n455), .A2(new_n434), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(new_n440), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT55), .Z(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n500), .A2(new_n188), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT53), .B1(new_n802), .B2(new_n823), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n810), .A2(new_n817), .ZN(new_n887));
  NOR4_X1   g701(.A1(new_n887), .A2(new_n792), .A3(new_n861), .A4(new_n801), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n885), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT56), .B1(new_n889), .B2(KEYINPUT119), .ZN(new_n890));
  INV_X1    g704(.A(new_n885), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n891), .B1(new_n862), .B2(new_n863), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT119), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n884), .B1(new_n890), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n868), .A2(G953), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT120), .Z(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n883), .A2(KEYINPUT56), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n898), .B1(new_n889), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT121), .B1(new_n895), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n894), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT56), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n904), .B1(new_n892), .B2(new_n893), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n883), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT121), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n906), .A2(new_n907), .A3(new_n900), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n902), .A2(new_n908), .ZN(G51));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n862), .A2(new_n863), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n763), .A2(new_n764), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n911), .A2(G902), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n289), .B(KEYINPUT57), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n862), .A2(new_n864), .A3(new_n863), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n864), .B1(new_n862), .B2(new_n863), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n914), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n670), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n913), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n910), .B1(new_n919), .B2(new_n898), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT54), .B1(new_n886), .B2(new_n888), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(new_n865), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n670), .B1(new_n922), .B2(new_n914), .ZN(new_n923));
  OAI211_X1 g737(.A(KEYINPUT122), .B(new_n897), .C1(new_n923), .C2(new_n913), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n920), .A2(new_n924), .ZN(G54));
  AND4_X1   g739(.A1(KEYINPUT58), .A2(new_n911), .A3(G475), .A4(G902), .ZN(new_n926));
  INV_X1    g740(.A(new_n386), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n898), .B1(new_n928), .B2(new_n929), .ZN(G60));
  AND2_X1   g744(.A1(new_n596), .A2(new_n597), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT123), .ZN(new_n932));
  NAND2_X1  g746(.A1(G478), .A2(G902), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT59), .Z(new_n934));
  NOR2_X1   g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n922), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n897), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n827), .A2(new_n865), .ZN(new_n938));
  INV_X1    g752(.A(new_n934), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n937), .B1(new_n940), .B2(new_n932), .ZN(G63));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT60), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n862), .B2(new_n863), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n898), .B1(new_n944), .B2(new_n618), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n570), .B2(new_n944), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT124), .B1(new_n944), .B2(new_n618), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n947), .A2(KEYINPUT61), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n946), .B(new_n948), .ZN(G66));
  INV_X1    g763(.A(new_n400), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n262), .B1(new_n950), .B2(G224), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n951), .B1(new_n792), .B2(new_n262), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n881), .B1(G898), .B2(new_n262), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n952), .B(new_n953), .Z(G69));
  OAI21_X1  g768(.A(new_n486), .B1(new_n494), .B2(KEYINPUT30), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(new_n381), .Z(new_n956));
  OAI211_X1 g770(.A(new_n717), .B(new_n815), .C1(new_n650), .C2(new_n656), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n685), .A2(new_n602), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n584), .A2(new_n756), .A3(new_n958), .ZN(new_n959));
  OAI22_X1  g773(.A1(new_n957), .A2(KEYINPUT62), .B1(new_n652), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n957), .A2(KEYINPUT62), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n957), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n960), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n772), .A2(new_n777), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n956), .B1(new_n966), .B2(G953), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n956), .B1(G900), .B2(G953), .ZN(new_n968));
  INV_X1    g782(.A(new_n739), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n710), .B2(new_n711), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n770), .B2(new_n771), .ZN(new_n971));
  INV_X1    g785(.A(new_n750), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n746), .A2(new_n805), .A3(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n772), .A2(new_n971), .A3(new_n777), .A4(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n968), .B1(new_n974), .B2(G953), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n967), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n262), .B1(G227), .B2(G900), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n977), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n967), .A2(new_n975), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n980), .ZN(G72));
  INV_X1    g795(.A(new_n826), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n982), .A2(new_n824), .A3(new_n820), .ZN(new_n983));
  XNOR2_X1  g797(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n479), .A2(new_n188), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n984), .B(new_n985), .Z(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n539), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n987), .B1(new_n988), .B2(new_n509), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n898), .B1(new_n983), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n986), .B1(new_n974), .B2(new_n792), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n529), .A2(new_n504), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n529), .A2(new_n504), .ZN(new_n994));
  INV_X1    g808(.A(new_n792), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n772), .A2(new_n777), .A3(new_n965), .A4(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n994), .B1(new_n996), .B2(new_n986), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n997), .A2(KEYINPUT127), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT127), .ZN(new_n999));
  AOI211_X1 g813(.A(new_n999), .B(new_n994), .C1(new_n996), .C2(new_n986), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n990), .B(new_n993), .C1(new_n998), .C2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(G57));
endmodule


