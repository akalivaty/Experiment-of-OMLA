//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n549, new_n551, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT66), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT67), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n451), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  NAND2_X1  g032(.A1(G113), .A2(G2104), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n458), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n459), .A2(G2105), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n465), .A2(G2105), .B1(G101), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g042(.A(KEYINPUT69), .B1(new_n459), .B2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(new_n461), .A3(G2104), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n473), .B1(new_n461), .B2(G2104), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n459), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n471), .A2(G137), .A3(new_n472), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n467), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  NAND3_X1  g054(.A1(new_n471), .A2(G2105), .A3(new_n476), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NAND4_X1  g057(.A1(new_n476), .A2(new_n472), .A3(new_n468), .A4(new_n470), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  NOR3_X1   g060(.A1(KEYINPUT70), .A2(G100), .A3(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(KEYINPUT70), .B1(G100), .B2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n482), .B(new_n485), .C1(new_n486), .C2(new_n488), .ZN(new_n489));
  OR2_X1    g064(.A1(new_n489), .A2(KEYINPUT71), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(KEYINPUT71), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(G162));
  OR2_X1    g068(.A1(new_n472), .A2(G114), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G126), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n480), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR4_X1   g075(.A1(new_n463), .A2(KEYINPUT4), .A3(new_n500), .A4(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT4), .B1(new_n483), .B2(new_n500), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(KEYINPUT72), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n471), .A2(G138), .A3(new_n472), .A4(new_n476), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT72), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT4), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n499), .B1(new_n503), .B2(new_n506), .ZN(G164));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G651), .ZN(new_n518));
  AND3_X1   g093(.A1(new_n516), .A2(new_n518), .A3(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G50), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n516), .A2(new_n518), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n512), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n515), .A2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  AND2_X1   g101(.A1(G63), .A2(G651), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n512), .A2(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n530), .B1(new_n528), .B2(new_n529), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n519), .A2(G51), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n522), .B2(new_n533), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n531), .A2(new_n534), .ZN(G286));
  INV_X1    g110(.A(G286), .ZN(G168));
  AOI22_X1  g111(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n514), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n519), .A2(G52), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n522), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(G171));
  INV_X1    g117(.A(G81), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n522), .A2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n514), .ZN(new_n546));
  AOI211_X1 g121(.A(new_n544), .B(new_n546), .C1(G43), .C2(new_n519), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  XOR2_X1   g125(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n551));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n549), .A2(new_n553), .ZN(G188));
  AND3_X1   g129(.A1(new_n512), .A2(new_n521), .A3(KEYINPUT76), .ZN(new_n555));
  AOI21_X1  g130(.A(KEYINPUT76), .B1(new_n512), .B2(new_n521), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n509), .A2(new_n511), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n557), .A2(G91), .B1(G651), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n519), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT9), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(KEYINPUT74), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n519), .A2(new_n567), .A3(G53), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(KEYINPUT75), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(KEYINPUT75), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT74), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n571), .B(KEYINPUT9), .C1(new_n563), .C2(new_n564), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n566), .A2(new_n569), .A3(new_n570), .A4(new_n572), .ZN(new_n573));
  AOI21_X1  g148(.A(KEYINPUT77), .B1(new_n562), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n562), .A2(KEYINPUT77), .A3(new_n573), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(G299));
  INV_X1    g152(.A(G171), .ZN(G301));
  INV_X1    g153(.A(G49), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT78), .B1(new_n563), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR3_X1   g157(.A1(new_n563), .A2(KEYINPUT78), .A3(new_n579), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n557), .A2(G87), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(G288));
  OAI21_X1  g161(.A(G86), .B1(new_n555), .B2(new_n556), .ZN(new_n587));
  NAND2_X1  g162(.A1(G73), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n559), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(new_n519), .B2(G48), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT79), .ZN(G305));
  AOI22_X1  g168(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(new_n514), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n519), .A2(G47), .ZN(new_n596));
  INV_X1    g171(.A(G85), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n522), .B2(new_n597), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n595), .A2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n557), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n555), .A2(new_n556), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n559), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(new_n519), .B2(G54), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n600), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n600), .B1(new_n612), .B2(G868), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  INV_X1    g190(.A(G299), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G297));
  XOR2_X1   g192(.A(G297), .B(KEYINPUT80), .Z(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(G148));
  NAND2_X1  g195(.A1(new_n612), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n547), .ZN(G323));
  XOR2_X1   g198(.A(KEYINPUT81), .B(KEYINPUT11), .Z(new_n624));
  XNOR2_X1  g199(.A(G323), .B(new_n624), .ZN(G282));
  OR2_X1    g200(.A1(G99), .A2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n626), .B(G2104), .C1(G111), .C2(new_n472), .ZN(new_n627));
  INV_X1    g202(.A(G135), .ZN(new_n628));
  INV_X1    g203(.A(G123), .ZN(new_n629));
  OAI221_X1 g204(.A(new_n627), .B1(new_n483), .B2(new_n628), .C1(new_n480), .C2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(G2096), .Z(new_n631));
  NAND3_X1  g206(.A1(new_n472), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2100), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n631), .A2(new_n635), .ZN(G156));
  INV_X1    g211(.A(KEYINPUT14), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2435), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n640), .B2(new_n639), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT16), .B(G1341), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n645), .B(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(G14), .B1(new_n642), .B2(new_n648), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n649), .B1(new_n642), .B2(new_n648), .ZN(G401));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT17), .Z(new_n652));
  XOR2_X1   g227(.A(G2084), .B(G2090), .Z(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2067), .B(G2678), .Z(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  OR3_X1    g233(.A1(new_n652), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  NOR3_X1   g234(.A1(new_n654), .A2(new_n651), .A3(new_n655), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT18), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n651), .A2(KEYINPUT82), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n651), .A2(KEYINPUT82), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n658), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n659), .A2(new_n661), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT83), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n665), .B(new_n667), .ZN(G227));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT84), .ZN(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT85), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n676), .A2(KEYINPUT20), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(KEYINPUT20), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n670), .A2(new_n671), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n680), .A2(new_n674), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n680), .A2(new_n674), .A3(new_n672), .ZN(new_n682));
  NAND4_X1  g257(.A1(new_n677), .A2(new_n678), .A3(new_n681), .A4(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1991), .B(G1996), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT87), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT86), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1981), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(new_n691), .ZN(G229));
  MUX2_X1   g267(.A(G6), .B(G305), .S(G16), .Z(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT90), .Z(new_n694));
  XOR2_X1   g269(.A(KEYINPUT32), .B(G1981), .Z(new_n695));
  OR2_X1    g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n694), .A2(new_n695), .ZN(new_n697));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G22), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G166), .B2(new_n698), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G1971), .ZN(new_n701));
  NOR2_X1   g276(.A1(G16), .A2(G23), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n584), .A2(new_n585), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(G16), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT33), .B(G1976), .Z(new_n705));
  AND2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n704), .A2(new_n705), .ZN(new_n707));
  NOR3_X1   g282(.A1(new_n701), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n696), .A2(new_n697), .A3(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT34), .Z(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G25), .ZN(new_n712));
  OAI21_X1  g287(.A(KEYINPUT88), .B1(G95), .B2(G2105), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NOR3_X1   g289(.A1(KEYINPUT88), .A2(G95), .A3(G2105), .ZN(new_n715));
  OAI221_X1 g290(.A(G2104), .B1(G107), .B2(new_n472), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT89), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n484), .A2(G131), .ZN(new_n718));
  INV_X1    g293(.A(G119), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n717), .B(new_n718), .C1(new_n719), .C2(new_n480), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n712), .B1(new_n721), .B2(new_n711), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT35), .B(G1991), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n698), .A2(G24), .ZN(new_n726));
  INV_X1    g301(.A(G290), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(new_n698), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G1986), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT92), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n730), .A2(KEYINPUT36), .ZN(new_n731));
  NOR4_X1   g306(.A1(new_n724), .A2(new_n725), .A3(new_n729), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n710), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n730), .B1(KEYINPUT91), .B2(KEYINPUT36), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n547), .A2(new_n698), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n698), .B2(G19), .ZN(new_n737));
  INV_X1    g312(.A(G1341), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G16), .A2(G21), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G168), .B2(G16), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n739), .B1(G1966), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G1966), .B2(new_n741), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n630), .A2(new_n711), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT95), .ZN(new_n745));
  OR2_X1    g320(.A1(G29), .A2(G32), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n481), .A2(G129), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n484), .A2(G141), .ZN(new_n748));
  NAND3_X1  g323(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT26), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n751), .A2(new_n752), .B1(G105), .B2(new_n466), .ZN(new_n753));
  NAND3_X1  g328(.A1(new_n747), .A2(new_n748), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n746), .B1(new_n754), .B2(new_n711), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT27), .B(G1996), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  NOR3_X1   g333(.A1(new_n745), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n484), .A2(G139), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n466), .A2(G103), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT25), .Z(new_n762));
  AND2_X1   g337(.A1(new_n460), .A2(new_n462), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n763), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n760), .B(new_n762), .C1(new_n472), .C2(new_n764), .ZN(new_n765));
  MUX2_X1   g340(.A(G33), .B(new_n765), .S(G29), .Z(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G2072), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT24), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n711), .B1(new_n768), .B2(G34), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT94), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n769), .A2(new_n770), .B1(new_n768), .B2(G34), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n770), .B2(new_n769), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n478), .B2(new_n711), .ZN(new_n773));
  INV_X1    g348(.A(G2084), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n767), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(G28), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n777), .A2(KEYINPUT30), .ZN(new_n778));
  AOI21_X1  g353(.A(G29), .B1(new_n777), .B2(KEYINPUT30), .ZN(new_n779));
  OR2_X1    g354(.A1(KEYINPUT31), .A2(G11), .ZN(new_n780));
  NAND2_X1  g355(.A1(KEYINPUT31), .A2(G11), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n778), .A2(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n737), .B2(new_n738), .ZN(new_n783));
  NOR2_X1   g358(.A1(G5), .A2(G16), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G171), .B2(G16), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1961), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n743), .A2(new_n759), .A3(new_n776), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n481), .A2(G128), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n484), .A2(G140), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n472), .A2(G116), .ZN(new_n791));
  OAI21_X1  g366(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n789), .B(new_n790), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n793), .A2(G29), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT93), .Z(new_n795));
  NAND2_X1  g370(.A1(new_n711), .A2(G26), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT28), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2067), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n698), .A2(G4), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n612), .B2(new_n698), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(G1348), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(G1348), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n773), .A2(new_n774), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT96), .Z(new_n805));
  NAND3_X1  g380(.A1(new_n802), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  NOR3_X1   g381(.A1(new_n788), .A2(new_n799), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n711), .A2(G35), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G162), .B2(new_n711), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT29), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G2090), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n698), .A2(G20), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT23), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(KEYINPUT23), .B1(new_n616), .B2(new_n698), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(new_n812), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G1956), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n711), .A2(G27), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G164), .B2(new_n711), .ZN(new_n819));
  MUX2_X1   g394(.A(new_n818), .B(new_n819), .S(KEYINPUT97), .Z(new_n820));
  INV_X1    g395(.A(G2078), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n807), .A2(new_n811), .A3(new_n817), .A4(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n735), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n733), .A2(new_n734), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n825), .A2(new_n826), .ZN(G311));
  INV_X1    g402(.A(new_n826), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n828), .A2(new_n735), .A3(new_n824), .ZN(G150));
  NAND2_X1  g404(.A1(G80), .A2(G543), .ZN(new_n830));
  INV_X1    g405(.A(G67), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n559), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G651), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(KEYINPUT99), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n519), .A2(G55), .ZN(new_n835));
  INV_X1    g410(.A(G93), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n834), .B(new_n835), .C1(new_n836), .C2(new_n522), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n833), .A2(KEYINPUT99), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(G860), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT37), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n611), .A2(new_n619), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT39), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT98), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT38), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n839), .B(new_n547), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n840), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n846), .A2(new_n848), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n842), .B1(new_n850), .B2(new_n851), .ZN(G145));
  NAND2_X1  g427(.A1(new_n502), .A2(KEYINPUT72), .ZN(new_n853));
  INV_X1    g428(.A(new_n501), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n853), .A2(new_n506), .A3(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n499), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n793), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n765), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n754), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n720), .B(new_n633), .Z(new_n861));
  OR2_X1    g436(.A1(G106), .A2(G2105), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n862), .B(G2104), .C1(G118), .C2(new_n472), .ZN(new_n863));
  INV_X1    g438(.A(G142), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n483), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(G130), .B2(new_n481), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n861), .B(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n860), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n860), .A2(new_n868), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n630), .B(new_n478), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n492), .B(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n868), .A2(KEYINPUT100), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n872), .B1(new_n874), .B2(new_n860), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n860), .B2(new_n874), .ZN(new_n876));
  INV_X1    g451(.A(G37), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n873), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g454(.A(new_n576), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n612), .B1(new_n880), .B2(new_n574), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n575), .A2(new_n576), .A3(new_n611), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(G299), .A2(KEYINPUT101), .A3(new_n612), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(KEYINPUT41), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n616), .A2(KEYINPUT102), .A3(new_n611), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n881), .A2(new_n890), .A3(new_n883), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n887), .A2(KEYINPUT103), .A3(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n621), .B(new_n848), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n886), .A2(new_n896), .A3(KEYINPUT41), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n893), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n886), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n894), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(G305), .B(G303), .ZN(new_n902));
  XNOR2_X1  g477(.A(G288), .B(new_n727), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n902), .B(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(new_n904), .B(KEYINPUT42), .Z(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(KEYINPUT104), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n901), .B2(new_n905), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT104), .B1(new_n901), .B2(new_n905), .ZN(new_n908));
  OAI21_X1  g483(.A(G868), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n839), .A2(G868), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(G295));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n909), .A2(new_n912), .A3(new_n910), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n912), .B1(new_n909), .B2(new_n910), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(G331));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n916));
  OAI21_X1  g491(.A(G286), .B1(new_n916), .B2(G171), .ZN(new_n917));
  NAND2_X1  g492(.A1(G171), .A2(new_n916), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n917), .B(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n848), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n849), .A2(new_n919), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n893), .A2(new_n897), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT108), .ZN(new_n925));
  INV_X1    g500(.A(new_n904), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT108), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n893), .A2(new_n927), .A3(new_n897), .A4(new_n923), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n921), .A2(new_n922), .A3(KEYINPUT109), .ZN(new_n929));
  OR3_X1    g504(.A1(new_n849), .A2(new_n919), .A3(KEYINPUT109), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n899), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n925), .A2(new_n926), .A3(new_n928), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT110), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n925), .A2(new_n928), .A3(new_n932), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(new_n904), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n924), .A2(KEYINPUT108), .B1(new_n899), .B2(new_n931), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT110), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n937), .A2(new_n938), .A3(new_n926), .A4(new_n928), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n934), .A2(new_n936), .A3(new_n877), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n941));
  AOI21_X1  g516(.A(G37), .B1(new_n933), .B2(KEYINPUT110), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n899), .A2(KEYINPUT41), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n888), .A2(KEYINPUT41), .A3(new_n891), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n944), .A2(new_n929), .A3(new_n930), .ZN(new_n945));
  OAI22_X1  g520(.A1(new_n943), .A2(new_n945), .B1(new_n886), .B2(new_n923), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n904), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT43), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n942), .A2(new_n947), .A3(new_n948), .A4(new_n939), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n941), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g525(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n942), .A2(new_n948), .A3(new_n939), .A4(new_n936), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n942), .A2(new_n939), .A3(new_n947), .ZN(new_n954));
  OAI211_X1 g529(.A(KEYINPUT44), .B(new_n953), .C1(new_n954), .C2(new_n948), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n952), .A2(new_n955), .ZN(G397));
  INV_X1    g531(.A(G1384), .ZN(new_n957));
  AND3_X1   g532(.A1(new_n504), .A2(new_n505), .A3(KEYINPUT4), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n505), .B1(new_n504), .B2(KEYINPUT4), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n958), .A2(new_n959), .A3(new_n501), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n957), .B1(new_n960), .B2(new_n499), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT45), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n467), .A2(G40), .A3(new_n477), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT111), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n793), .B(G2067), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g543(.A1(new_n968), .A2(KEYINPUT112), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(KEYINPUT112), .ZN(new_n970));
  INV_X1    g545(.A(new_n966), .ZN(new_n971));
  XOR2_X1   g546(.A(new_n754), .B(G1996), .Z(new_n972));
  OAI211_X1 g547(.A(new_n969), .B(new_n970), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n720), .B(new_n723), .ZN(new_n974));
  XOR2_X1   g549(.A(new_n974), .B(KEYINPUT113), .Z(new_n975));
  NOR2_X1   g550(.A1(new_n975), .A2(new_n971), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n727), .A2(new_n687), .ZN(new_n977));
  NAND2_X1  g552(.A1(G290), .A2(G1986), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n971), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n973), .A2(new_n976), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(G1384), .B1(new_n855), .B2(new_n856), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT45), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT111), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n964), .B(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n963), .A2(new_n821), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n857), .A2(new_n988), .A3(new_n957), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(new_n990), .A3(new_n984), .ZN(new_n991));
  INV_X1    g566(.A(G1961), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NOR3_X1   g568(.A1(new_n964), .A2(new_n986), .A3(G2078), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n963), .A2(new_n982), .A3(new_n994), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n987), .A2(G301), .A3(new_n993), .A4(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT125), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n965), .B1(new_n961), .B2(new_n962), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n999), .A2(KEYINPUT53), .A3(new_n821), .A4(new_n982), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n987), .A2(new_n1000), .A3(new_n993), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(G171), .ZN(new_n1002));
  AOI22_X1  g577(.A1(new_n985), .A2(new_n986), .B1(new_n992), .B2(new_n991), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n1003), .A2(KEYINPUT125), .A3(G301), .A4(new_n995), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n998), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  XOR2_X1   g580(.A(KEYINPUT124), .B(KEYINPUT54), .Z(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n987), .A2(new_n993), .A3(new_n995), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT126), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT126), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1003), .A2(new_n1010), .A3(new_n995), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1009), .A2(G171), .A3(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1003), .A2(G301), .A3(new_n1000), .ZN(new_n1013));
  AND2_X1   g588(.A1(new_n1013), .A2(KEYINPUT54), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1966), .B1(new_n999), .B2(new_n982), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n989), .A2(new_n990), .A3(new_n774), .A4(new_n984), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(G8), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(G286), .A2(G8), .ZN(new_n1020));
  XOR2_X1   g595(.A(new_n1020), .B(KEYINPUT123), .Z(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n963), .A2(new_n982), .A3(new_n984), .ZN(new_n1025));
  INV_X1    g600(.A(G1966), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1021), .B1(new_n1027), .B2(new_n1017), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1028), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1024), .B1(new_n1029), .B2(new_n1023), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n981), .A2(new_n984), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n703), .A2(G1976), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(G8), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT52), .ZN(new_n1034));
  INV_X1    g609(.A(G1976), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT52), .B1(G288), .B2(new_n1035), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1031), .A2(new_n1032), .A3(new_n1036), .A4(G8), .ZN(new_n1037));
  INV_X1    g612(.A(new_n591), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n512), .A2(new_n521), .A3(G86), .ZN(new_n1039));
  OAI21_X1  g614(.A(G1981), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G1981), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n587), .A2(new_n1041), .A3(new_n591), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1040), .A2(new_n1042), .A3(KEYINPUT49), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT49), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1045), .A2(G8), .A3(new_n1031), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1034), .A2(new_n1037), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G8), .ZN(new_n1048));
  INV_X1    g623(.A(G1971), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n984), .B1(new_n981), .B2(KEYINPUT45), .ZN(new_n1050));
  NOR3_X1   g625(.A1(G164), .A2(new_n962), .A3(G1384), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1049), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g627(.A(KEYINPUT114), .B(G2090), .Z(new_n1053));
  NAND4_X1  g628(.A1(new_n989), .A2(new_n990), .A3(new_n984), .A4(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1048), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1056), .B1(G166), .B2(new_n1048), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1057), .A2(KEYINPUT116), .ZN(new_n1058));
  NAND3_X1  g633(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1057), .A2(KEYINPUT116), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1058), .A2(new_n1061), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1047), .B1(new_n1055), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1066), .A2(G8), .A3(new_n1064), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1055), .A2(KEYINPUT117), .A3(new_n1064), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1065), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1007), .A2(new_n1015), .A3(new_n1030), .A4(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n562), .A2(new_n573), .ZN(new_n1073));
  NAND2_X1  g648(.A1(KEYINPUT121), .A2(KEYINPUT57), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g650(.A1(KEYINPUT121), .A2(KEYINPUT57), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1075), .B(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G1956), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n991), .A2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT56), .B(G2072), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n999), .A2(new_n982), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1078), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT122), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1078), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1078), .A2(new_n1080), .A3(new_n1082), .A4(KEYINPUT122), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1085), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT61), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G1348), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1031), .ZN(new_n1094));
  INV_X1    g669(.A(G2067), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n991), .A2(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n612), .B1(new_n1096), .B2(KEYINPUT60), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(KEYINPUT60), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1097), .B(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT58), .B(G1341), .ZN(new_n1100));
  OAI22_X1  g675(.A1(new_n1025), .A2(G1996), .B1(new_n1094), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n547), .ZN(new_n1102));
  XNOR2_X1  g677(.A(new_n1102), .B(KEYINPUT59), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1088), .A2(KEYINPUT61), .A3(new_n1083), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1092), .A2(new_n1099), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1088), .B1(new_n611), .B2(new_n1096), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1106), .A2(new_n1085), .A3(new_n1089), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1072), .A2(KEYINPUT127), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1030), .A2(new_n1071), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT127), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1109), .A2(new_n1110), .A3(new_n1007), .A4(new_n1015), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1071), .A2(G171), .A3(new_n1001), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(KEYINPUT62), .B2(new_n1030), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1030), .A2(KEYINPUT62), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1108), .A2(new_n1111), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1046), .A2(new_n1035), .A3(new_n703), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1042), .ZN(new_n1117));
  OAI211_X1 g692(.A(G8), .B(new_n1031), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1034), .A2(new_n1037), .A3(new_n1046), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(G1971), .B1(new_n999), .B2(new_n982), .ZN(new_n1122));
  AND4_X1   g697(.A1(new_n984), .A2(new_n989), .A3(new_n990), .A4(new_n1053), .ZN(new_n1123));
  OAI21_X1  g698(.A(G8), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1064), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1120), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1019), .A2(G286), .ZN(new_n1127));
  AND4_X1   g702(.A1(KEYINPUT117), .A2(new_n1066), .A3(G8), .A4(new_n1064), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT117), .B1(new_n1055), .B2(new_n1064), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1126), .B(new_n1127), .C1(new_n1128), .C2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT63), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1130), .A2(KEYINPUT118), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT118), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1119), .A2(new_n1134), .A3(new_n1126), .A4(new_n1127), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1133), .A2(new_n1131), .A3(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1132), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1133), .A2(new_n1135), .A3(KEYINPUT119), .A4(new_n1131), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1121), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1115), .B1(new_n1140), .B2(KEYINPUT120), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n1142));
  AOI211_X1 g717(.A(new_n1142), .B(new_n1121), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n980), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n971), .A2(new_n977), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT48), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n1146), .A2(new_n973), .A3(new_n976), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT46), .ZN(new_n1148));
  OR3_X1    g723(.A1(new_n971), .A2(new_n1148), .A3(G1996), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n966), .B1(new_n754), .B2(new_n967), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1148), .B1(new_n971), .B2(G1996), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  XOR2_X1   g727(.A(new_n1152), .B(KEYINPUT47), .Z(new_n1153));
  OR2_X1    g728(.A1(new_n720), .A2(new_n723), .ZN(new_n1154));
  OAI22_X1  g729(.A1(new_n973), .A2(new_n1154), .B1(G2067), .B2(new_n793), .ZN(new_n1155));
  AOI211_X1 g730(.A(new_n1147), .B(new_n1153), .C1(new_n966), .C2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1144), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g732(.A(G319), .ZN(new_n1159));
  NOR4_X1   g733(.A1(G229), .A2(new_n1159), .A3(G401), .A4(G227), .ZN(new_n1160));
  NAND3_X1  g734(.A1(new_n950), .A2(new_n878), .A3(new_n1160), .ZN(G225));
  INV_X1    g735(.A(G225), .ZN(G308));
endmodule


