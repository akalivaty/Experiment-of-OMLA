//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n844, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957, new_n958;
  INV_X1    g000(.A(G22gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT2), .ZN(new_n204));
  OR2_X1    g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n203), .A2(KEYINPUT73), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G155gat), .B(G162gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n207), .A2(new_n210), .A3(new_n208), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT29), .ZN(new_n215));
  XNOR2_X1  g014(.A(G197gat), .B(G204gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(G211gat), .B(G218gat), .ZN(new_n217));
  INV_X1    g016(.A(G211gat), .ZN(new_n218));
  OR2_X1    g017(.A1(KEYINPUT68), .A2(G218gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(KEYINPUT68), .A2(G218gat), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n216), .B(new_n217), .C1(new_n221), .C2(KEYINPUT22), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  AND2_X1   g022(.A1(KEYINPUT68), .A2(G218gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(KEYINPUT68), .A2(G218gat), .ZN(new_n225));
  OAI21_X1  g024(.A(G211gat), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT22), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n217), .B1(new_n228), .B2(new_n216), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n215), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n214), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n216), .B1(new_n221), .B2(KEYINPUT22), .ZN(new_n233));
  INV_X1    g032(.A(new_n217), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n222), .ZN(new_n236));
  AND3_X1   g035(.A1(new_n207), .A2(new_n210), .A3(new_n208), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n210), .B1(new_n207), .B2(new_n208), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n231), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n236), .B1(new_n215), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G228gat), .ZN(new_n241));
  INV_X1    g040(.A(G233gat), .ZN(new_n242));
  OAI22_X1  g041(.A1(new_n232), .A2(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n239), .A2(new_n215), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n235), .A2(KEYINPUT69), .A3(new_n222), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT69), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n246), .B1(new_n223), .B2(new_n229), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n244), .A2(new_n245), .A3(new_n247), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n237), .A2(new_n238), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT29), .B1(new_n235), .B2(new_n222), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n249), .B1(new_n250), .B2(KEYINPUT3), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n241), .A2(new_n242), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n248), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n202), .B1(new_n243), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n243), .A2(new_n253), .A3(new_n202), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G78gat), .B(G106gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(KEYINPUT31), .B(G50gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT80), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n260), .B1(new_n254), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n255), .A2(new_n261), .A3(new_n256), .A4(new_n260), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT65), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n269));
  INV_X1    g068(.A(G169gat), .ZN(new_n270));
  INV_X1    g069(.A(G176gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT23), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n268), .A2(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G190gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(G183gat), .ZN(new_n276));
  INV_X1    g075(.A(G183gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n277), .A2(G190gat), .ZN(new_n278));
  OAI21_X1  g077(.A(KEYINPUT24), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n280), .A2(KEYINPUT24), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n273), .A2(G176gat), .ZN(new_n283));
  OR2_X1    g082(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n274), .A2(new_n279), .A3(new_n282), .A4(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT25), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n271), .A2(KEYINPUT23), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT25), .B1(new_n290), .B2(G169gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n292), .A2(new_n274), .A3(new_n279), .A4(new_n282), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT27), .B(G183gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(new_n275), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT28), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n295), .A2(KEYINPUT28), .A3(new_n275), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OR3_X1    g099(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n269), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n301), .B(new_n302), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n300), .A2(new_n280), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT29), .B1(new_n294), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G226gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n308), .A2(new_n242), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT71), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT24), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n277), .A2(G190gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n275), .A2(G183gat), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NOR3_X1   g113(.A1(new_n314), .A2(new_n291), .A3(new_n281), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n288), .A2(new_n287), .B1(new_n315), .B2(new_n274), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n305), .A2(new_n280), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n317), .B1(new_n298), .B2(new_n299), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n215), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT71), .ZN(new_n320));
  INV_X1    g119(.A(new_n309), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n310), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n309), .B1(new_n316), .B2(new_n318), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT72), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI211_X1 g125(.A(KEYINPUT72), .B(new_n309), .C1(new_n316), .C2(new_n318), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n323), .A2(new_n236), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT70), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n324), .A2(new_n329), .B1(new_n319), .B2(new_n321), .ZN(new_n330));
  OAI211_X1 g129(.A(KEYINPUT70), .B(new_n309), .C1(new_n316), .C2(new_n318), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n247), .A2(new_n245), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n328), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G8gat), .B(G36gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(G64gat), .B(G92gat), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n337), .B(new_n338), .Z(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n328), .A2(new_n335), .A3(new_n339), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(KEYINPUT30), .A3(new_n342), .ZN(new_n343));
  OR3_X1    g142(.A1(new_n336), .A2(KEYINPUT30), .A3(new_n340), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n212), .A2(KEYINPUT3), .A3(new_n213), .ZN(new_n346));
  XOR2_X1   g145(.A(G127gat), .B(G134gat), .Z(new_n347));
  XNOR2_X1  g146(.A(G113gat), .B(G120gat), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n347), .B1(KEYINPUT1), .B2(new_n348), .ZN(new_n349));
  XOR2_X1   g148(.A(G113gat), .B(G120gat), .Z(new_n350));
  INV_X1    g149(.A(KEYINPUT1), .ZN(new_n351));
  XNOR2_X1  g150(.A(G127gat), .B(G134gat), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n239), .A2(new_n346), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT4), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n356), .B1(new_n249), .B2(new_n354), .ZN(new_n357));
  AND2_X1   g156(.A1(new_n349), .A2(new_n353), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n214), .A2(new_n358), .A3(KEYINPUT4), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n355), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G225gat), .A2(G233gat), .ZN(new_n361));
  OR2_X1    g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n249), .B(new_n354), .ZN(new_n363));
  INV_X1    g162(.A(new_n361), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT39), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI211_X1 g166(.A(KEYINPUT81), .B(KEYINPUT39), .C1(new_n363), .C2(new_n364), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n362), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  XOR2_X1   g168(.A(KEYINPUT77), .B(KEYINPUT0), .Z(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(KEYINPUT78), .ZN(new_n371));
  XNOR2_X1  g170(.A(G1gat), .B(G29gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G57gat), .B(G85gat), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n373), .B(new_n374), .Z(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(new_n362), .B2(KEYINPUT39), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT40), .ZN(new_n377));
  OR3_X1    g176(.A1(new_n369), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n375), .ZN(new_n379));
  NOR3_X1   g178(.A1(new_n249), .A2(new_n356), .A3(new_n354), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT4), .B1(new_n214), .B2(new_n358), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT75), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n382), .A2(new_n383), .A3(new_n361), .A4(new_n355), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n355), .A2(new_n357), .A3(new_n361), .A4(new_n359), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT75), .ZN(new_n386));
  XOR2_X1   g185(.A(KEYINPUT76), .B(KEYINPUT5), .Z(new_n387));
  AOI21_X1  g186(.A(new_n387), .B1(new_n363), .B2(new_n364), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n384), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n360), .A2(KEYINPUT79), .A3(new_n361), .A4(new_n387), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT79), .ZN(new_n391));
  INV_X1    g190(.A(new_n387), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n391), .B1(new_n385), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n379), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT82), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI211_X1 g196(.A(KEYINPUT82), .B(new_n379), .C1(new_n389), .C2(new_n394), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n377), .B1(new_n369), .B2(new_n376), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n378), .A2(new_n397), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n265), .B1(new_n345), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n386), .A3(new_n388), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(new_n393), .A3(new_n390), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(KEYINPUT6), .A3(new_n379), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n389), .A2(new_n394), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT6), .B1(new_n406), .B2(new_n375), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(new_n397), .A3(new_n398), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT83), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT83), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n407), .A2(new_n397), .A3(new_n410), .A4(new_n398), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n405), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n336), .A2(KEYINPUT37), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n340), .B1(new_n336), .B2(KEYINPUT37), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT38), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n340), .A2(KEYINPUT37), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n341), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n319), .A2(new_n321), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n324), .A2(new_n329), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n418), .A2(new_n419), .A3(new_n331), .A4(new_n333), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT84), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT84), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n330), .A2(new_n422), .A3(new_n331), .A4(new_n333), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n326), .A2(new_n327), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n424), .B1(new_n310), .B2(new_n322), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n421), .B(new_n423), .C1(new_n425), .C2(new_n236), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT38), .B1(new_n426), .B2(KEYINPUT37), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n417), .A2(new_n427), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n415), .A2(new_n428), .A3(new_n342), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n401), .B1(new_n412), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n407), .A2(new_n395), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n343), .A2(new_n344), .B1(new_n431), .B2(new_n404), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n432), .A2(new_n265), .ZN(new_n433));
  XNOR2_X1  g232(.A(G15gat), .B(G43gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(G71gat), .B(G99gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(G227gat), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n438), .A2(new_n242), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n354), .B1(new_n316), .B2(new_n318), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n294), .A2(new_n358), .A3(new_n306), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n437), .B1(new_n443), .B2(KEYINPUT33), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT32), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n441), .A2(new_n442), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n445), .B1(new_n446), .B2(new_n439), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT66), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n316), .A2(new_n318), .A3(new_n354), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n358), .B1(new_n294), .B2(new_n306), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n439), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT32), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT33), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT66), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n452), .A2(new_n454), .A3(new_n455), .A4(new_n437), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n448), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n436), .A2(new_n453), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n451), .A2(KEYINPUT32), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT34), .B1(new_n446), .B2(new_n439), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT34), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n441), .A2(new_n442), .A3(new_n463), .A4(new_n440), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT67), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n460), .A2(new_n462), .A3(new_n464), .ZN(new_n468));
  AOI211_X1 g267(.A(new_n467), .B(new_n468), .C1(new_n448), .C2(new_n456), .ZN(new_n469));
  INV_X1    g268(.A(new_n468), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT67), .B1(new_n457), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n466), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT36), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n436), .B1(new_n451), .B2(new_n453), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n455), .B1(new_n474), .B2(new_n452), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n444), .A2(KEYINPUT66), .A3(new_n447), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n470), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n467), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n457), .A2(KEYINPUT67), .A3(new_n470), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT36), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(new_n466), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n473), .A2(new_n482), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n430), .A2(new_n433), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n472), .A2(KEYINPUT85), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT85), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n480), .A2(new_n486), .A3(new_n466), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT35), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n345), .A2(new_n489), .A3(new_n265), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n412), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT86), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n469), .A2(new_n471), .ZN(new_n493));
  INV_X1    g292(.A(new_n465), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n448), .A2(new_n456), .B1(new_n447), .B2(new_n459), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n265), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n492), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n461), .A2(new_n465), .B1(new_n264), .B2(new_n263), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n480), .A2(new_n498), .A3(KEYINPUT86), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n497), .A2(new_n432), .A3(new_n499), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n488), .A2(new_n491), .B1(new_n500), .B2(KEYINPUT35), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT87), .B1(new_n484), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n412), .A2(new_n429), .ZN(new_n503));
  INV_X1    g302(.A(new_n401), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n433), .ZN(new_n506));
  INV_X1    g305(.A(new_n483), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n500), .A2(KEYINPUT35), .ZN(new_n509));
  INV_X1    g308(.A(new_n398), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT82), .B1(new_n403), .B2(new_n379), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n410), .B1(new_n512), .B2(new_n407), .ZN(new_n513));
  INV_X1    g312(.A(new_n411), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n404), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n345), .A2(new_n489), .A3(new_n265), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n515), .A2(new_n516), .A3(new_n485), .A4(new_n487), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n509), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT87), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n508), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(G15gat), .B(G22gat), .Z(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G1gat), .ZN(new_n522));
  INV_X1    g321(.A(G1gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT16), .ZN(new_n524));
  OAI221_X1 g323(.A(new_n522), .B1(KEYINPUT90), .B2(G8gat), .C1(new_n521), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n526));
  XOR2_X1   g325(.A(new_n525), .B(new_n526), .Z(new_n527));
  INV_X1    g326(.A(KEYINPUT15), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT14), .B(G29gat), .ZN(new_n529));
  INV_X1    g328(.A(G36gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G29gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n532), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  XOR2_X1   g333(.A(G43gat), .B(G50gat), .Z(new_n535));
  INV_X1    g334(.A(KEYINPUT89), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n531), .A2(new_n535), .A3(new_n533), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n528), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g339(.A(KEYINPUT15), .B1(new_n534), .B2(new_n537), .ZN(new_n541));
  NOR3_X1   g340(.A1(new_n527), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n540), .A2(new_n541), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT17), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n542), .B1(new_n527), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G229gat), .A2(G233gat), .ZN(new_n546));
  AOI21_X1  g345(.A(KEYINPUT18), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n527), .B(new_n543), .Z(new_n548));
  XNOR2_X1  g347(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(new_n546), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n547), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n545), .A2(KEYINPUT18), .A3(new_n546), .ZN(new_n552));
  AND2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G113gat), .B(G141gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(G197gat), .ZN(new_n555));
  XOR2_X1   g354(.A(KEYINPUT11), .B(G169gat), .Z(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(KEYINPUT88), .B(KEYINPUT12), .Z(new_n558));
  XNOR2_X1  g357(.A(new_n557), .B(new_n558), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n553), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n551), .A2(new_n559), .A3(new_n552), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT92), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n551), .A2(KEYINPUT92), .A3(new_n559), .A4(new_n552), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G85gat), .A2(G92gat), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n567), .B(KEYINPUT7), .Z(new_n568));
  XNOR2_X1  g367(.A(G99gat), .B(G106gat), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT95), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n568), .B1(new_n571), .B2(KEYINPUT96), .ZN(new_n572));
  NAND2_X1  g371(.A1(G99gat), .A2(G106gat), .ZN(new_n573));
  INV_X1    g372(.A(G85gat), .ZN(new_n574));
  INV_X1    g373(.A(G92gat), .ZN(new_n575));
  AOI22_X1  g374(.A1(KEYINPUT8), .A2(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n576), .B(KEYINPUT94), .Z(new_n577));
  NAND2_X1  g376(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n571), .A2(KEYINPUT96), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n572), .B(new_n577), .C1(KEYINPUT96), .C2(new_n571), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT97), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(new_n543), .ZN(new_n584));
  NAND3_X1  g383(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n543), .B(KEYINPUT17), .Z(new_n586));
  OAI211_X1 g385(.A(new_n584), .B(new_n585), .C1(new_n586), .C2(new_n583), .ZN(new_n587));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G134gat), .B(G162gat), .ZN(new_n590));
  AOI21_X1  g389(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n589), .A2(new_n592), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT21), .ZN(new_n597));
  XNOR2_X1  g396(.A(G57gat), .B(G64gat), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G71gat), .B(G78gat), .Z(new_n601));
  OR2_X1    g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n527), .B1(new_n597), .B2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT93), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n607));
  INV_X1    g406(.A(G155gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n606), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n604), .A2(new_n597), .ZN(new_n611));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G127gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  OR2_X1    g415(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n610), .A2(new_n616), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n604), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n582), .B1(KEYINPUT98), .B2(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n620), .A2(KEYINPUT98), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT99), .B(KEYINPUT10), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n583), .A2(KEYINPUT10), .A3(new_n620), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT100), .ZN(new_n629));
  NAND2_X1  g428(.A1(G230gat), .A2(G233gat), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n631), .B1(new_n627), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n623), .A2(new_n630), .ZN(new_n635));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(G176gat), .B(G204gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  AND2_X1   g437(.A1(new_n635), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n635), .B1(new_n628), .B2(new_n631), .ZN(new_n641));
  INV_X1    g440(.A(new_n638), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n596), .A2(new_n619), .A3(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n502), .A2(new_n520), .A3(new_n566), .A4(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n431), .A2(new_n404), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g453(.A(new_n345), .B1(new_n648), .B2(new_n649), .ZN(new_n655));
  INV_X1    g454(.A(G8gat), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(KEYINPUT16), .B(G8gat), .Z(new_n658));
  NAND3_X1  g457(.A1(new_n655), .A2(KEYINPUT42), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(KEYINPUT42), .B1(new_n655), .B2(new_n658), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n657), .B(new_n659), .C1(new_n660), .C2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n661), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(KEYINPUT103), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n657), .A2(new_n659), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n660), .A2(new_n661), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n666), .A2(new_n667), .A3(new_n668), .A4(new_n663), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n665), .A2(new_n669), .ZN(G1325gat));
  AOI21_X1  g469(.A(G15gat), .B1(new_n650), .B2(new_n488), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT104), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n483), .A2(G15gat), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n672), .B1(new_n650), .B2(new_n673), .ZN(G1326gat));
  INV_X1    g473(.A(new_n265), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n650), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT43), .B(G22gat), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1327gat));
  AND2_X1   g477(.A1(new_n502), .A2(new_n520), .ZN(new_n679));
  INV_X1    g478(.A(new_n644), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n619), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(new_n595), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n679), .A2(new_n566), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n683), .A2(new_n532), .A3(new_n652), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT45), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n686), .B1(new_n432), .B2(new_n265), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n651), .A2(new_n345), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n688), .A2(KEYINPUT107), .A3(new_n675), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n690), .A2(new_n430), .A3(new_n483), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT108), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n518), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n509), .A2(KEYINPUT108), .A3(new_n517), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n691), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT109), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n595), .B(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT110), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n505), .A2(new_n507), .A3(new_n687), .A4(new_n689), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n509), .A2(KEYINPUT108), .A3(new_n517), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT108), .B1(new_n509), .B2(new_n517), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n704), .A2(new_n705), .A3(new_n698), .A4(new_n697), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n700), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n502), .A2(new_n520), .A3(new_n596), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n708), .A2(new_n709), .A3(KEYINPUT44), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n709), .B1(new_n708), .B2(KEYINPUT44), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n707), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n566), .A2(KEYINPUT105), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT105), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n560), .A2(new_n565), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n681), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n712), .A2(new_n652), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G29gat), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n685), .A2(new_n719), .ZN(G1328gat));
  INV_X1    g519(.A(new_n345), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n712), .A2(new_n721), .A3(new_n717), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n530), .B1(new_n722), .B2(KEYINPUT112), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(KEYINPUT112), .B2(new_n722), .ZN(new_n724));
  AOI21_X1  g523(.A(G36gat), .B1(KEYINPUT111), .B2(KEYINPUT46), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n683), .A2(new_n721), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(KEYINPUT111), .A2(KEYINPUT46), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n724), .A2(new_n728), .ZN(G1329gat));
  AOI21_X1  g528(.A(G43gat), .B1(new_n683), .B2(new_n488), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n730), .B1(KEYINPUT113), .B2(KEYINPUT47), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n712), .A2(G43gat), .A3(new_n483), .A4(new_n717), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(KEYINPUT113), .A2(KEYINPUT47), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n733), .B(new_n734), .Z(G1330gat));
  NAND3_X1  g534(.A1(new_n712), .A2(new_n675), .A3(new_n717), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT115), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n712), .A2(KEYINPUT115), .A3(new_n675), .A4(new_n717), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n738), .A2(G50gat), .A3(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n679), .A2(new_n566), .A3(new_n682), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n741), .A2(G50gat), .A3(new_n265), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n740), .A2(KEYINPUT48), .A3(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT114), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n736), .A2(G50gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n743), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT48), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n742), .B1(new_n736), .B2(G50gat), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n750), .A2(KEYINPUT114), .A3(KEYINPUT48), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n744), .B1(new_n749), .B2(new_n751), .ZN(G1331gat));
  INV_X1    g551(.A(new_n619), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n595), .A2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n716), .ZN(new_n755));
  NOR4_X1   g554(.A1(new_n695), .A2(new_n754), .A3(new_n680), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n651), .B(KEYINPUT116), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g559(.A1(new_n756), .A2(new_n721), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n762));
  XOR2_X1   g561(.A(KEYINPUT49), .B(G64gat), .Z(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n761), .B2(new_n763), .ZN(G1333gat));
  NAND2_X1  g563(.A1(new_n756), .A2(new_n483), .ZN(new_n765));
  INV_X1    g564(.A(new_n488), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n766), .A2(G71gat), .ZN(new_n767));
  AOI22_X1  g566(.A1(new_n765), .A2(G71gat), .B1(new_n756), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g568(.A1(new_n756), .A2(new_n675), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n753), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n772), .A2(new_n596), .A3(new_n704), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT51), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n772), .A2(KEYINPUT51), .A3(new_n704), .A4(new_n596), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n680), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n777), .A2(new_n574), .A3(new_n652), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n712), .A2(new_n644), .A3(new_n772), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n779), .A2(new_n652), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n778), .B1(new_n780), .B2(new_n574), .ZN(G1336gat));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n345), .A2(G92gat), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT117), .B1(new_n777), .B2(new_n783), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n779), .A2(new_n721), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n782), .B(new_n784), .C1(new_n785), .C2(new_n575), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n575), .B1(new_n779), .B2(new_n721), .ZN(new_n787));
  INV_X1    g586(.A(new_n784), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT52), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(new_n789), .ZN(G1337gat));
  NAND2_X1  g589(.A1(new_n779), .A2(new_n483), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G99gat), .ZN(new_n792));
  INV_X1    g591(.A(new_n777), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n766), .A2(G99gat), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(G1338gat));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n793), .A2(G106gat), .A3(new_n265), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n779), .A2(new_n675), .ZN(new_n799));
  XNOR2_X1  g598(.A(KEYINPUT118), .B(G106gat), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n796), .B(new_n798), .C1(new_n799), .C2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n801), .B1(new_n779), .B2(new_n675), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT53), .B1(new_n803), .B2(new_n797), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(G1339gat));
  XNOR2_X1  g604(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n627), .A2(new_n630), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n642), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT54), .B1(new_n627), .B2(new_n630), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n808), .B1(new_n634), .B2(new_n810), .ZN(new_n811));
  AOI22_X1  g610(.A1(new_n811), .A2(KEYINPUT55), .B1(new_n634), .B2(new_n639), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n809), .B1(new_n629), .B2(new_n633), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n814), .B2(new_n808), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n713), .A2(new_n812), .A3(new_n815), .A4(new_n715), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n545), .A2(new_n546), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n548), .A2(new_n550), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n557), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(KEYINPUT120), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n820), .B1(new_n563), .B2(new_n564), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n644), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n697), .B1(new_n816), .B2(new_n822), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n595), .B(KEYINPUT109), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n812), .A2(new_n815), .A3(new_n821), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n619), .B1(new_n823), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n645), .A2(new_n716), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n675), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n829), .A2(new_n652), .A3(new_n345), .A4(new_n488), .ZN(new_n830));
  INV_X1    g629(.A(G113gat), .ZN(new_n831));
  INV_X1    g630(.A(new_n566), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n757), .B1(new_n827), .B2(new_n828), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n497), .A2(new_n499), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(new_n721), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n755), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n833), .B1(new_n838), .B2(new_n831), .ZN(G1340gat));
  INV_X1    g638(.A(G120gat), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n830), .A2(new_n840), .A3(new_n680), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n837), .A2(new_n644), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n841), .B1(new_n842), .B2(new_n840), .ZN(G1341gat));
  INV_X1    g642(.A(G127gat), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n837), .A2(new_n844), .A3(new_n753), .ZN(new_n845));
  OAI21_X1  g644(.A(G127gat), .B1(new_n830), .B2(new_n619), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1342gat));
  INV_X1    g646(.A(G134gat), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n595), .A2(new_n721), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n834), .A2(new_n848), .A3(new_n835), .A4(new_n849), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n851));
  OAI21_X1  g650(.A(G134gat), .B1(new_n830), .B2(new_n595), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(KEYINPUT56), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(G1343gat));
  NAND2_X1  g653(.A1(new_n507), .A2(new_n675), .ZN(new_n855));
  XOR2_X1   g654(.A(new_n855), .B(KEYINPUT122), .Z(new_n856));
  NAND2_X1  g655(.A1(new_n834), .A2(new_n856), .ZN(new_n857));
  NOR4_X1   g656(.A1(new_n857), .A2(G141gat), .A3(new_n721), .A4(new_n832), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n815), .A2(KEYINPUT121), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n860), .B(new_n813), .C1(new_n814), .C2(new_n808), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n812), .A2(new_n859), .A3(new_n566), .A4(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n596), .B1(new_n862), .B2(new_n822), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n619), .B1(new_n863), .B2(new_n826), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n265), .B1(new_n864), .B2(new_n828), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT57), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI211_X1 g666(.A(KEYINPUT57), .B(new_n265), .C1(new_n827), .C2(new_n828), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n483), .A2(new_n651), .A3(new_n721), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n867), .A2(new_n869), .A3(new_n755), .A4(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n858), .B1(new_n871), .B2(G141gat), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT58), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n870), .B1(new_n865), .B2(new_n866), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n874), .A2(new_n868), .A3(new_n832), .ZN(new_n875));
  INV_X1    g674(.A(G141gat), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n857), .A2(KEYINPUT123), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n832), .A2(G141gat), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n834), .A2(new_n880), .A3(new_n856), .ZN(new_n881));
  AND4_X1   g680(.A1(new_n345), .A2(new_n878), .A3(new_n879), .A4(new_n881), .ZN(new_n882));
  OAI22_X1  g681(.A1(new_n872), .A2(new_n873), .B1(new_n877), .B2(new_n882), .ZN(G1344gat));
  NOR2_X1   g682(.A1(new_n680), .A2(G148gat), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n878), .A2(new_n345), .A3(new_n881), .A4(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n265), .B1(new_n827), .B2(new_n828), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n887), .A2(new_n866), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n265), .A2(KEYINPUT57), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n862), .A2(new_n822), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n595), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n825), .A2(new_n595), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n753), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n754), .A2(new_n566), .A3(new_n644), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n889), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n888), .A2(new_n644), .A3(new_n870), .A4(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n886), .B1(new_n896), .B2(G148gat), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n886), .A2(G148gat), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n874), .A2(new_n868), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(new_n644), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n885), .B1(new_n897), .B2(new_n900), .ZN(G1345gat));
  NAND4_X1  g700(.A1(new_n878), .A2(new_n345), .A3(new_n753), .A4(new_n881), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n753), .A2(G155gat), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT124), .ZN(new_n904));
  AOI22_X1  g703(.A1(new_n902), .A2(new_n608), .B1(new_n899), .B2(new_n904), .ZN(G1346gat));
  INV_X1    g704(.A(G162gat), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n878), .A2(new_n906), .A3(new_n849), .A4(new_n881), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n874), .A2(new_n868), .A3(new_n824), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(new_n906), .ZN(G1347gat));
  NAND2_X1  g708(.A1(new_n757), .A2(new_n721), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n766), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT125), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n829), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(G169gat), .B1(new_n913), .B2(new_n832), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n652), .B1(new_n827), .B2(new_n828), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n835), .A2(new_n721), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n755), .A2(new_n284), .A3(new_n285), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n914), .B1(new_n917), .B2(new_n918), .ZN(G1348gat));
  OAI21_X1  g718(.A(G176gat), .B1(new_n913), .B2(new_n680), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n644), .A2(new_n271), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n917), .B2(new_n921), .ZN(G1349gat));
  OAI21_X1  g721(.A(G183gat), .B1(new_n913), .B2(new_n619), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n753), .A2(new_n295), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n917), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g725(.A(G190gat), .B1(new_n913), .B2(new_n595), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n927), .A2(KEYINPUT61), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n927), .A2(KEYINPUT61), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n697), .A2(new_n275), .ZN(new_n930));
  OAI22_X1  g729(.A1(new_n928), .A2(new_n929), .B1(new_n917), .B2(new_n930), .ZN(G1351gat));
  NOR2_X1   g730(.A1(new_n910), .A2(new_n483), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n895), .B(new_n932), .C1(new_n887), .C2(new_n866), .ZN(new_n933));
  OAI21_X1  g732(.A(G197gat), .B1(new_n933), .B2(new_n832), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n915), .A2(new_n721), .A3(new_n675), .A4(new_n507), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n716), .A2(G197gat), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(KEYINPUT126), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n934), .A2(new_n940), .A3(new_n937), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n941), .ZN(G1352gat));
  NOR3_X1   g741(.A1(new_n935), .A2(G204gat), .A3(new_n680), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT62), .ZN(new_n944));
  OAI21_X1  g743(.A(G204gat), .B1(new_n933), .B2(new_n680), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1353gat));
  NAND2_X1  g745(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n947));
  OAI21_X1  g746(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n948));
  INV_X1    g747(.A(new_n933), .ZN(new_n949));
  AOI211_X1 g748(.A(new_n947), .B(new_n948), .C1(new_n949), .C2(new_n753), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n888), .A2(new_n753), .A3(new_n895), .A4(new_n932), .ZN(new_n951));
  INV_X1    g750(.A(new_n948), .ZN(new_n952));
  AOI22_X1  g751(.A1(new_n951), .A2(new_n952), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n753), .A2(new_n218), .ZN(new_n954));
  OAI22_X1  g753(.A1(new_n950), .A2(new_n953), .B1(new_n935), .B2(new_n954), .ZN(G1354gat));
  NOR2_X1   g754(.A1(new_n935), .A2(new_n824), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n956), .A2(G218gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n595), .B1(new_n219), .B2(new_n220), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n949), .B2(new_n958), .ZN(G1355gat));
endmodule


