//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 0 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1117, new_n1118,
    new_n1119;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT67), .Z(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT1), .ZN(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  AND2_X1   g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n457), .A2(KEYINPUT68), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(KEYINPUT68), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n456), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT69), .Z(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(KEYINPUT70), .A2(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT3), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(G137), .A3(new_n464), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n471), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n469), .B1(new_n476), .B2(new_n462), .ZN(G160));
  NAND2_X1  g052(.A1(new_n472), .A2(new_n464), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(new_n462), .B2(G112), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT71), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n472), .A2(new_n464), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G2105), .ZN(new_n485));
  NOR3_X1   g060(.A1(new_n478), .A2(KEYINPUT71), .A3(new_n462), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G124), .ZN(new_n488));
  OAI221_X1 g063(.A(new_n480), .B1(new_n481), .B2(new_n482), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT72), .ZN(G162));
  NAND3_X1  g065(.A1(new_n462), .A2(KEYINPUT4), .A3(G138), .ZN(new_n491));
  NAND2_X1  g066(.A1(G126), .A2(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n472), .A2(new_n493), .A3(new_n464), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(new_n464), .A3(new_n466), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT73), .B1(new_n462), .B2(G114), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT73), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n501), .A2(new_n502), .A3(G2105), .ZN(new_n503));
  OR2_X1    g078(.A1(G102), .A2(G2105), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n500), .A2(new_n503), .A3(G2104), .A4(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n494), .A2(new_n499), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(KEYINPUT74), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT74), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(KEYINPUT5), .A3(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G62), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT76), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n508), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT6), .B(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n514), .A2(new_n519), .ZN(new_n520));
  XOR2_X1   g095(.A(KEYINPUT75), .B(G88), .Z(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n520), .A2(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n518), .A2(new_n524), .ZN(G166));
  INV_X1    g100(.A(new_n520), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G89), .ZN(new_n527));
  INV_X1    g102(.A(new_n522), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n532));
  NAND4_X1  g107(.A1(new_n527), .A2(new_n529), .A3(new_n531), .A4(new_n532), .ZN(G286));
  INV_X1    g108(.A(G286), .ZN(G168));
  AOI22_X1  g109(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n508), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(KEYINPUT77), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n526), .A2(G90), .B1(new_n528), .B2(G52), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(KEYINPUT77), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(G301));
  INV_X1    g115(.A(G301), .ZN(G171));
  AOI22_X1  g116(.A1(new_n526), .A2(G81), .B1(new_n528), .B2(G43), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n514), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n508), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(KEYINPUT78), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT78), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n544), .A2(new_n542), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(new_n528), .A2(G53), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(KEYINPUT79), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n556), .B(new_n558), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n526), .A2(KEYINPUT80), .A3(G91), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT80), .ZN(new_n561));
  INV_X1    g136(.A(G91), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n520), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n514), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n565));
  OAI211_X1 g140(.A(new_n559), .B(new_n564), .C1(new_n508), .C2(new_n565), .ZN(G299));
  INV_X1    g141(.A(G166), .ZN(G303));
  NAND2_X1  g142(.A1(new_n526), .A2(G87), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n528), .A2(G49), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  AOI22_X1  g146(.A1(new_n526), .A2(G86), .B1(new_n528), .B2(G48), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n514), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n573));
  OR2_X1    g148(.A1(new_n573), .A2(new_n508), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(G305));
  AOI22_X1  g150(.A1(new_n526), .A2(G85), .B1(new_n528), .B2(G47), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT81), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n508), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT82), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n580), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n526), .A2(G92), .ZN(new_n585));
  XOR2_X1   g160(.A(KEYINPUT83), .B(KEYINPUT10), .Z(new_n586));
  XNOR2_X1  g161(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n514), .A2(G66), .ZN(new_n588));
  INV_X1    g163(.A(G79), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n589), .B2(new_n509), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(G54), .B2(new_n528), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n584), .B1(new_n593), .B2(G868), .ZN(G284));
  OAI21_X1  g169(.A(new_n584), .B1(new_n593), .B2(G868), .ZN(G321));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(G299), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(new_n596), .B2(G168), .ZN(G297));
  OAI21_X1  g173(.A(new_n597), .B1(new_n596), .B2(G168), .ZN(G280));
  INV_X1    g174(.A(G860), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n592), .B1(G559), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT84), .ZN(G148));
  NOR2_X1   g177(.A1(new_n549), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n593), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT85), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n603), .B1(new_n607), .B2(G868), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT86), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n474), .A2(new_n462), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n464), .A2(new_n466), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g188(.A(new_n613), .B(KEYINPUT12), .Z(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2100), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT87), .B(KEYINPUT13), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n487), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n618), .A2(G123), .B1(G135), .B2(new_n479), .ZN(new_n619));
  OR2_X1    g194(.A1(G99), .A2(G2105), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n620), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G2096), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n617), .A2(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2430), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2435), .ZN(new_n627));
  XOR2_X1   g202(.A(G2427), .B(G2438), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(KEYINPUT14), .ZN(new_n630));
  XOR2_X1   g205(.A(G2451), .B(G2454), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT16), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n630), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G1341), .B(G1348), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n635), .B(new_n636), .Z(new_n637));
  AND2_X1   g212(.A1(new_n637), .A2(G14), .ZN(G401));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2067), .B(G2678), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2072), .B(G2078), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT88), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(KEYINPUT17), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n645), .B1(new_n641), .B2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT89), .Z(new_n649));
  NAND3_X1  g224(.A1(new_n642), .A2(new_n643), .A3(new_n639), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT18), .Z(new_n651));
  NAND3_X1  g226(.A1(new_n647), .A2(new_n639), .A3(new_n641), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n649), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(new_n623), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2100), .ZN(G227));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  XOR2_X1   g232(.A(G1956), .B(G2474), .Z(new_n658));
  XOR2_X1   g233(.A(G1961), .B(G1966), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n658), .A2(new_n659), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n665), .A2(new_n657), .A3(new_n660), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n663), .B(new_n666), .C1(new_n657), .C2(new_n665), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT21), .B(G1986), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G1991), .B(G1996), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT22), .B(G1981), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n671), .B(new_n672), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G229));
  NAND2_X1  g249(.A1(new_n593), .A2(G16), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(G4), .B2(G16), .ZN(new_n676));
  INV_X1    g251(.A(G1348), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(G29), .A2(G32), .ZN(new_n679));
  AND2_X1   g254(.A1(new_n618), .A2(G129), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n479), .A2(G141), .ZN(new_n681));
  NAND3_X1  g256(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT26), .Z(new_n683));
  INV_X1    g258(.A(G105), .ZN(new_n684));
  OAI211_X1 g259(.A(new_n681), .B(new_n683), .C1(new_n684), .C2(new_n611), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n679), .B1(new_n686), .B2(G29), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT27), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT97), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n689), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n619), .A2(G29), .A3(new_n621), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n693), .A2(KEYINPUT98), .ZN(new_n694));
  NAND4_X1  g269(.A1(new_n678), .A2(new_n690), .A3(new_n691), .A4(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(KEYINPUT98), .B2(new_n693), .ZN(new_n696));
  INV_X1    g271(.A(G16), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G19), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(new_n549), .B2(new_n697), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT94), .B(G1341), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n479), .A2(G139), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT25), .Z(new_n704));
  INV_X1    g279(.A(new_n612), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n705), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n702), .B(new_n704), .C1(new_n462), .C2(new_n706), .ZN(new_n707));
  MUX2_X1   g282(.A(G33), .B(new_n707), .S(G29), .Z(new_n708));
  XOR2_X1   g283(.A(KEYINPUT95), .B(G2072), .Z(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(G29), .A2(G35), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G162), .B2(G29), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT29), .B(G2090), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND4_X1  g289(.A1(new_n696), .A2(new_n701), .A3(new_n710), .A4(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT28), .ZN(new_n716));
  INV_X1    g291(.A(G26), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n717), .B2(G29), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(G29), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n618), .A2(G128), .B1(G140), .B2(new_n479), .ZN(new_n720));
  NOR2_X1   g295(.A1(G104), .A2(G2105), .ZN(new_n721));
  OAI21_X1  g296(.A(G2104), .B1(new_n462), .B2(G116), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n719), .B1(new_n723), .B2(G29), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n718), .B1(new_n724), .B2(new_n716), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n725), .A2(G2067), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(G2067), .ZN(new_n727));
  INV_X1    g302(.A(G1961), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT99), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G5), .B2(G16), .ZN(new_n730));
  OR3_X1    g305(.A1(new_n729), .A2(G5), .A3(G16), .ZN(new_n731));
  OAI211_X1 g306(.A(new_n730), .B(new_n731), .C1(G301), .C2(new_n697), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n727), .B1(new_n728), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(G299), .A2(G16), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n697), .A2(KEYINPUT23), .A3(G20), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT23), .ZN(new_n736));
  INV_X1    g311(.A(G20), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(G16), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n734), .A2(new_n735), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1956), .ZN(new_n740));
  NAND2_X1  g315(.A1(G168), .A2(G16), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G16), .B2(G21), .ZN(new_n742));
  INV_X1    g317(.A(G1966), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(G164), .A2(G29), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G27), .B2(G29), .ZN(new_n746));
  INV_X1    g321(.A(G2078), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n747), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT30), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n750), .A2(G28), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n750), .A2(G28), .ZN(new_n752));
  OR3_X1    g327(.A1(new_n751), .A2(new_n752), .A3(G29), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n744), .A2(new_n748), .A3(new_n749), .A4(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n740), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT31), .B(G11), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n742), .A2(new_n743), .ZN(new_n757));
  INV_X1    g332(.A(G2084), .ZN(new_n758));
  NOR2_X1   g333(.A1(KEYINPUT24), .A2(G34), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(KEYINPUT24), .A2(G34), .ZN(new_n761));
  AOI21_X1  g336(.A(G29), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI22_X1  g337(.A1(G160), .A2(G29), .B1(KEYINPUT96), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(KEYINPUT96), .B2(new_n762), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n676), .A2(new_n677), .B1(new_n758), .B2(new_n764), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n755), .A2(new_n756), .A3(new_n757), .A4(new_n765), .ZN(new_n766));
  NOR4_X1   g341(.A1(new_n715), .A2(new_n726), .A3(new_n733), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n732), .A2(new_n728), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n767), .B(new_n768), .C1(new_n758), .C2(new_n764), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT100), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n697), .A2(G22), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G166), .B2(new_n697), .ZN(new_n773));
  INV_X1    g348(.A(G1971), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G16), .A2(G23), .ZN(new_n776));
  INV_X1    g351(.A(G288), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(G16), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT33), .B(G1976), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n697), .A2(G6), .ZN(new_n781));
  INV_X1    g356(.A(G305), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(new_n697), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT32), .B(G1981), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n775), .A2(new_n780), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n479), .A2(G131), .ZN(new_n787));
  OR2_X1    g362(.A1(G95), .A2(G2105), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n788), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n789));
  INV_X1    g364(.A(G119), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n787), .B(new_n789), .C1(new_n487), .C2(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT91), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT92), .ZN(new_n793));
  MUX2_X1   g368(.A(G25), .B(new_n793), .S(G29), .Z(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT35), .B(G1991), .ZN(new_n795));
  OAI221_X1 g370(.A(KEYINPUT93), .B1(KEYINPUT34), .B2(new_n786), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n795), .B2(new_n794), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n786), .A2(KEYINPUT34), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n697), .A2(G24), .ZN(new_n799));
  INV_X1    g374(.A(G290), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n697), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(G1986), .Z(new_n802));
  NAND3_X1  g377(.A1(new_n797), .A2(new_n798), .A3(new_n802), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT36), .Z(new_n804));
  NOR2_X1   g379(.A1(new_n771), .A2(new_n804), .ZN(G311));
  XNOR2_X1  g380(.A(new_n769), .B(KEYINPUT100), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n803), .B(KEYINPUT36), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(new_n807), .ZN(G150));
  AOI22_X1  g383(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT101), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n810), .A2(G651), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n526), .A2(G93), .B1(new_n528), .B2(G55), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G860), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT104), .B(KEYINPUT37), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n813), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(new_n545), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n549), .A2(new_n813), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT102), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT102), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n818), .A2(new_n822), .A3(new_n819), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n592), .A2(new_n604), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT38), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n824), .B(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT39), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT103), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n600), .B1(new_n827), .B2(new_n828), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n816), .B1(new_n830), .B2(new_n831), .ZN(G145));
  AOI22_X1  g407(.A1(new_n618), .A2(G130), .B1(G142), .B2(new_n479), .ZN(new_n833));
  NOR2_X1   g408(.A1(G106), .A2(G2105), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(G162), .B(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n622), .B(G160), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n792), .B(new_n686), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n707), .B(G164), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n839), .B(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n723), .B(new_n614), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT105), .B(G37), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g423(.A1(new_n824), .A2(KEYINPUT106), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n824), .A2(KEYINPUT106), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n607), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n593), .B(G299), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT41), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n824), .A2(KEYINPUT106), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n855), .A2(new_n606), .A3(new_n849), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n852), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  NOR3_X1   g432(.A1(new_n850), .A2(new_n851), .A3(new_n607), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n606), .B1(new_n855), .B2(new_n849), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n857), .B1(new_n860), .B2(new_n853), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n861), .A2(KEYINPUT42), .ZN(new_n862));
  XNOR2_X1  g437(.A(G305), .B(KEYINPUT107), .ZN(new_n863));
  XNOR2_X1  g438(.A(G290), .B(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(G166), .B(new_n777), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n865), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n800), .A2(new_n863), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n581), .A2(new_n582), .A3(new_n863), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n861), .A2(KEYINPUT42), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n862), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n872), .B1(new_n862), .B2(new_n873), .ZN(new_n875));
  OAI21_X1  g450(.A(G868), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(G868), .B2(new_n817), .ZN(G295));
  OAI21_X1  g452(.A(new_n876), .B1(G868), .B2(new_n817), .ZN(G331));
  XNOR2_X1  g453(.A(G301), .B(G286), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n824), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT109), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n821), .A2(new_n823), .A3(new_n879), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n854), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n883), .A2(new_n882), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n881), .A2(new_n853), .A3(new_n883), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n872), .ZN(new_n890));
  INV_X1    g465(.A(G37), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n871), .A2(new_n887), .A3(new_n888), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT110), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n854), .B1(new_n883), .B2(new_n881), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n884), .A2(new_n886), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n898), .B1(new_n899), .B2(new_n853), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n892), .B(new_n846), .C1(new_n900), .C2(new_n871), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n901), .A2(new_n894), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n893), .A2(KEYINPUT110), .A3(new_n894), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n897), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT44), .B1(new_n893), .B2(new_n894), .ZN(new_n907));
  AND2_X1   g482(.A1(new_n901), .A2(KEYINPUT43), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n909), .A2(KEYINPUT111), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT111), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n907), .A2(new_n908), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n906), .B1(new_n910), .B2(new_n912), .ZN(G397));
  XOR2_X1   g488(.A(KEYINPUT112), .B(G1384), .Z(new_n914));
  AND2_X1   g489(.A1(new_n506), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(KEYINPUT113), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT45), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(G160), .A2(G40), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT114), .ZN(new_n920));
  AOI21_X1  g495(.A(G2105), .B1(new_n473), .B2(new_n475), .ZN(new_n921));
  INV_X1    g496(.A(G40), .ZN(new_n922));
  NOR4_X1   g497(.A1(new_n921), .A2(KEYINPUT114), .A3(new_n922), .A4(new_n469), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n918), .A2(new_n925), .ZN(new_n926));
  XOR2_X1   g501(.A(new_n686), .B(G1996), .Z(new_n927));
  XNOR2_X1  g502(.A(new_n723), .B(G2067), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n795), .ZN(new_n930));
  OR2_X1    g505(.A1(new_n792), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n792), .A2(new_n930), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n932), .A3(new_n926), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(G290), .B(G1986), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n934), .B1(new_n926), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT121), .ZN(new_n937));
  INV_X1    g512(.A(G1384), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n506), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT50), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n506), .A2(KEYINPUT117), .A3(new_n938), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT117), .B1(new_n506), .B2(new_n938), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n941), .B1(new_n944), .B2(new_n940), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n937), .B1(new_n945), .B2(new_n925), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT117), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n939), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n506), .A2(KEYINPUT117), .A3(new_n938), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n940), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n941), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT114), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n953), .B1(G160), .B2(G40), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n954), .A2(new_n923), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n952), .A2(KEYINPUT121), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n946), .A2(new_n677), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT122), .ZN(new_n958));
  INV_X1    g533(.A(new_n944), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n960), .A2(G2067), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n957), .A2(new_n958), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n958), .B1(new_n957), .B2(new_n962), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT60), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n952), .A2(KEYINPUT121), .A3(new_n955), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT121), .B1(new_n952), .B2(new_n955), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n969), .A2(new_n970), .A3(G1348), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT122), .B1(new_n971), .B2(new_n961), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n957), .A2(new_n958), .A3(new_n962), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(new_n966), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT124), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n974), .A2(new_n975), .A3(new_n593), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n975), .B1(new_n974), .B2(new_n593), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n968), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(KEYINPUT58), .B(G1341), .Z(new_n979));
  NAND2_X1  g554(.A1(new_n960), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n915), .A2(KEYINPUT45), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT115), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n939), .A2(new_n917), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(new_n955), .A3(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n980), .B1(new_n984), .B2(G1996), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n549), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT123), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n987), .A2(KEYINPUT59), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n986), .B(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n987), .A2(KEYINPUT59), .ZN(new_n990));
  INV_X1    g565(.A(new_n939), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n940), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n955), .B(new_n992), .C1(new_n959), .C2(new_n940), .ZN(new_n993));
  INV_X1    g568(.A(G1956), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  XOR2_X1   g570(.A(KEYINPUT56), .B(G2072), .Z(new_n996));
  OAI21_X1  g571(.A(new_n995), .B1(new_n984), .B2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(G299), .B(KEYINPUT57), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n997), .A2(new_n998), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT61), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1001), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT61), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n1004), .A3(new_n999), .ZN(new_n1005));
  AOI22_X1  g580(.A1(new_n989), .A2(new_n990), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n963), .A2(new_n964), .A3(KEYINPUT60), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT124), .B1(new_n1007), .B2(new_n592), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n974), .A2(new_n975), .A3(new_n593), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(new_n967), .A3(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n978), .A2(new_n1006), .A3(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1001), .A2(new_n592), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1000), .B1(new_n1012), .B2(new_n965), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n1011), .A2(KEYINPUT125), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT125), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1015));
  XNOR2_X1  g590(.A(G305), .B(G1981), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT49), .ZN(new_n1017));
  OR2_X1    g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g593(.A(KEYINPUT119), .B(G8), .Z(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(new_n955), .B2(new_n959), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1018), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT120), .ZN(new_n1024));
  INV_X1    g599(.A(G1976), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1021), .B1(new_n1025), .B2(G288), .ZN(new_n1026));
  AOI211_X1 g601(.A(KEYINPUT52), .B(new_n1026), .C1(new_n1025), .C2(G288), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1026), .A2(KEYINPUT52), .ZN(new_n1028));
  OR3_X1    g603(.A1(new_n1024), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n984), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n982), .A2(KEYINPUT116), .A3(new_n955), .A4(new_n983), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(new_n747), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n991), .A2(KEYINPUT45), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n955), .B(new_n1036), .C1(new_n959), .C2(KEYINPUT45), .ZN(new_n1037));
  OR3_X1    g612(.A1(new_n1037), .A2(new_n1034), .A3(G2078), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n946), .A2(new_n728), .A3(new_n956), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1035), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(G171), .ZN(new_n1041));
  INV_X1    g616(.A(new_n919), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1034), .A2(G2078), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n918), .A2(new_n982), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1035), .A2(new_n1039), .A3(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1041), .B1(G171), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1029), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G8), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n774), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n945), .A2(new_n925), .ZN(new_n1052));
  INV_X1    g627(.A(G2090), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1049), .B1(new_n1051), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(G166), .A2(new_n1049), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1056), .B(KEYINPUT55), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1058), .B(KEYINPUT118), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1045), .A2(G171), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT127), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OR2_X1    g637(.A1(new_n1040), .A2(G171), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1045), .A2(KEYINPUT127), .A3(G171), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1062), .A2(new_n1063), .A3(KEYINPUT54), .A4(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1052), .A2(new_n758), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1037), .A2(new_n743), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n1019), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT51), .ZN(new_n1070));
  NAND2_X1  g645(.A1(G286), .A2(new_n1019), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1049), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1073));
  XOR2_X1   g648(.A(new_n1071), .B(KEYINPUT126), .Z(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT51), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1071), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1072), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1051), .B1(G2090), .B2(new_n993), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n1019), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1057), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1077), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1048), .A2(new_n1059), .A3(new_n1065), .A4(new_n1081), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1014), .A2(new_n1015), .A3(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1069), .A2(G286), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1084), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1029), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n777), .A2(new_n1025), .ZN(new_n1087));
  OAI22_X1  g662(.A1(new_n1024), .A2(new_n1087), .B1(G1981), .B2(G305), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1086), .A2(KEYINPUT63), .B1(new_n1021), .B2(new_n1088), .ZN(new_n1089));
  XOR2_X1   g664(.A(new_n1058), .B(KEYINPUT118), .Z(new_n1090));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1077), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1072), .B(KEYINPUT62), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1084), .ZN(new_n1095));
  OAI22_X1  g670(.A1(new_n1094), .A2(new_n1041), .B1(KEYINPUT63), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1090), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1089), .B1(new_n1098), .B2(new_n1029), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n936), .B1(new_n1083), .B2(new_n1099), .ZN(new_n1100));
  NOR4_X1   g675(.A1(G290), .A2(G1986), .A3(new_n925), .A4(new_n918), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1101), .A2(KEYINPUT48), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1101), .A2(KEYINPUT48), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n1102), .A2(new_n934), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n686), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n926), .B1(new_n928), .B2(new_n1105), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n918), .A2(G1996), .A3(new_n925), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1107), .A2(KEYINPUT46), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(KEYINPUT46), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1106), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  XOR2_X1   g685(.A(new_n1110), .B(KEYINPUT47), .Z(new_n1111));
  NAND2_X1  g686(.A1(new_n929), .A2(new_n930), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n1112), .A2(new_n793), .B1(G2067), .B2(new_n723), .ZN(new_n1113));
  AOI211_X1 g688(.A(new_n1104), .B(new_n1111), .C1(new_n926), .C2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1100), .A2(new_n1114), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g690(.A(G319), .ZN(new_n1117));
  AOI21_X1  g691(.A(new_n1117), .B1(new_n845), .B2(new_n846), .ZN(new_n1118));
  NOR2_X1   g692(.A1(G227), .A2(G401), .ZN(new_n1119));
  NAND4_X1  g693(.A1(new_n904), .A2(new_n1118), .A3(new_n673), .A4(new_n1119), .ZN(G225));
  INV_X1    g694(.A(G225), .ZN(G308));
endmodule


