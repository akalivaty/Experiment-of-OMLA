//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n584, new_n585, new_n586, new_n588, new_n589,
    new_n590, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n622, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1199;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT67), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT68), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(new_n454), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(G2106), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n455), .A2(new_n449), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G101), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT69), .B1(new_n472), .B2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(new_n463), .A3(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n471), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NOR3_X1   g051(.A1(new_n468), .A2(new_n470), .A3(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(new_n464), .A2(new_n465), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT70), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G136), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n479), .A2(new_n463), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n463), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n481), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT71), .Z(G162));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n488), .A2(new_n490), .A3(G2104), .ZN(new_n491));
  AND2_X1   g066(.A1(G126), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n464), .B2(new_n465), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n497));
  NAND2_X1  g072(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G138), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n496), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OR2_X1    g075(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n498), .A2(G138), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n503), .A2(new_n504), .A3(new_n463), .A4(new_n495), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n494), .B1(new_n500), .B2(new_n505), .ZN(G164));
  INV_X1    g081(.A(KEYINPUT73), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n507), .B1(new_n508), .B2(G651), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(KEYINPUT73), .A3(KEYINPUT6), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n513), .B1(new_n510), .B2(KEYINPUT6), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n508), .A2(KEYINPUT74), .A3(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT5), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n519), .B2(KEYINPUT75), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT75), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(KEYINPUT5), .A3(G543), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G88), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n517), .A2(new_n518), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G50), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n520), .A2(new_n522), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n528), .A2(G62), .ZN(new_n529));
  AND2_X1   g104(.A1(G75), .A2(G543), .ZN(new_n530));
  OAI211_X1 g105(.A(KEYINPUT76), .B(G651), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT76), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n528), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n533), .B2(new_n510), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n525), .A2(new_n527), .A3(new_n531), .A4(new_n534), .ZN(G303));
  INV_X1    g110(.A(G303), .ZN(G166));
  AND2_X1   g111(.A1(new_n512), .A2(new_n516), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n537), .A2(G89), .A3(new_n528), .ZN(new_n538));
  XNOR2_X1  g113(.A(KEYINPUT77), .B(KEYINPUT7), .ZN(new_n539));
  AND3_X1   g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n540), .ZN(new_n542));
  AND2_X1   g117(.A1(G63), .A2(G651), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n541), .A2(new_n542), .B1(new_n528), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n537), .A2(G51), .A3(G543), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n538), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(G168));
  AND2_X1   g122(.A1(new_n528), .A2(G64), .ZN(new_n548));
  AND2_X1   g123(.A1(G77), .A2(G543), .ZN(new_n549));
  OAI21_X1  g124(.A(G651), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g125(.A(KEYINPUT78), .B(G90), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n537), .A2(new_n528), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n537), .A2(G52), .A3(G543), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(G171));
  NAND2_X1  g130(.A1(G68), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G56), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n523), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G651), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n537), .A2(G43), .A3(G543), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n537), .A2(G81), .A3(new_n528), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  NAND2_X1  g142(.A1(new_n537), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G53), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT9), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n526), .A2(new_n571), .A3(G53), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT79), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n523), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n528), .A2(KEYINPUT79), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(G78), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n518), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n524), .A2(G91), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n573), .A2(new_n581), .A3(new_n582), .ZN(G299));
  NAND2_X1  g158(.A1(new_n554), .A2(KEYINPUT80), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT80), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n550), .A2(new_n552), .A3(new_n553), .A4(new_n585), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n584), .A2(new_n586), .ZN(G301));
  NAND2_X1  g162(.A1(new_n546), .A2(KEYINPUT81), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT81), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n538), .A2(new_n544), .A3(new_n545), .A4(new_n589), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n588), .A2(new_n590), .ZN(G286));
  NAND4_X1  g166(.A1(new_n528), .A2(new_n512), .A3(new_n516), .A4(G87), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n512), .A2(new_n516), .A3(G49), .A4(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(G651), .B1(new_n528), .B2(G74), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(G288));
  INV_X1    g170(.A(G61), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n596), .B1(new_n520), .B2(new_n522), .ZN(new_n597));
  AND2_X1   g172(.A1(G73), .A2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND4_X1  g174(.A1(new_n528), .A2(new_n512), .A3(new_n516), .A4(G86), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n512), .A2(new_n516), .A3(G48), .A4(G543), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(G305));
  NAND2_X1  g177(.A1(new_n526), .A2(G47), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n524), .A2(G85), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  OAI211_X1 g180(.A(new_n603), .B(new_n604), .C1(new_n510), .C2(new_n605), .ZN(G290));
  NAND3_X1  g181(.A1(new_n537), .A2(G92), .A3(new_n528), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n524), .A2(KEYINPUT10), .A3(G92), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n609), .A2(new_n610), .B1(G54), .B2(new_n526), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n528), .B(new_n575), .ZN(new_n612));
  INV_X1    g187(.A(G66), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g189(.A1(G79), .A2(G543), .ZN(new_n615));
  OAI21_X1  g190(.A(G651), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  MUX2_X1   g192(.A(new_n617), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g193(.A(new_n617), .B(G301), .S(G868), .Z(G321));
  MUX2_X1   g194(.A(G299), .B(G286), .S(G868), .Z(G297));
  XNOR2_X1  g195(.A(G297), .B(KEYINPUT82), .ZN(G280));
  INV_X1    g196(.A(new_n617), .ZN(new_n622));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n562), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  INV_X1    g204(.A(G111), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G2105), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(new_n480), .B2(G135), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT85), .ZN(new_n633));
  AND3_X1   g208(.A1(new_n482), .A2(new_n633), .A3(G123), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n633), .B1(new_n482), .B2(G123), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(KEYINPUT86), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(KEYINPUT86), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n473), .A2(new_n475), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(new_n503), .ZN(new_n642));
  XOR2_X1   g217(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(KEYINPUT13), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT84), .ZN(new_n646));
  AOI22_X1  g221(.A1(new_n644), .A2(new_n645), .B1(new_n646), .B2(G2100), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n645), .B2(new_n644), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n646), .A2(G2100), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n640), .A2(new_n650), .ZN(G156));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT87), .B(G2438), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n652), .B(new_n653), .Z(new_n654));
  XNOR2_X1  g229(.A(G2427), .B(G2430), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(KEYINPUT14), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2451), .B(G2454), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT16), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1341), .B(G1348), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n658), .B(new_n662), .Z(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  AND3_X1   g241(.A1(new_n665), .A2(G14), .A3(new_n666), .ZN(G401));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(G2072), .A2(G2078), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n442), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g248(.A1(new_n669), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT18), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n671), .A2(KEYINPUT88), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(KEYINPUT88), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n676), .A2(new_n677), .A3(new_n673), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n671), .B(KEYINPUT17), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n678), .B(new_n669), .C1(new_n679), .C2(new_n673), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n679), .A2(new_n673), .A3(new_n668), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n675), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G2096), .B(G2100), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G227));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT90), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1971), .B(G1976), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT20), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n690), .A2(new_n691), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT89), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  OR3_X1    g273(.A1(new_n689), .A2(new_n692), .A3(new_n695), .ZN(new_n699));
  AND3_X1   g274(.A1(new_n694), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G1981), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G1986), .ZN(new_n702));
  INV_X1    g277(.A(G1981), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n700), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G1986), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n687), .B1(new_n702), .B2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1991), .B(G1996), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n702), .A2(new_n706), .A3(new_n687), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n709), .ZN(new_n712));
  INV_X1    g287(.A(new_n710), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n707), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n711), .A2(new_n714), .ZN(G229));
  XNOR2_X1  g290(.A(KEYINPUT91), .B(G29), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(G162), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G35), .B2(new_n717), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(KEYINPUT29), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n719), .A2(KEYINPUT29), .ZN(new_n722));
  OAI21_X1  g297(.A(G2090), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n722), .ZN(new_n724));
  INV_X1    g299(.A(G2090), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n724), .A2(new_n725), .A3(new_n720), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G32), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n480), .A2(G141), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n482), .A2(G129), .ZN(new_n731));
  NAND3_X1  g306(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT26), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n641), .A2(G105), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n730), .A2(new_n731), .A3(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n729), .B1(new_n738), .B2(new_n728), .ZN(new_n739));
  XNOR2_X1  g314(.A(KEYINPUT27), .B(G1996), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT99), .ZN(new_n741));
  INV_X1    g316(.A(G16), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G5), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G171), .B2(new_n742), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n739), .A2(new_n741), .B1(G1961), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n742), .A2(G21), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G168), .B2(new_n742), .ZN(new_n747));
  OAI221_X1 g322(.A(new_n745), .B1(G1961), .B2(new_n744), .C1(G1966), .C2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n717), .A2(G27), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G164), .B2(new_n717), .ZN(new_n750));
  XOR2_X1   g325(.A(KEYINPUT100), .B(G2078), .Z(new_n751));
  XOR2_X1   g326(.A(new_n750), .B(new_n751), .Z(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G1966), .B2(new_n747), .ZN(new_n753));
  INV_X1    g328(.A(G28), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(KEYINPUT30), .ZN(new_n755));
  AOI21_X1  g330(.A(G29), .B1(new_n754), .B2(KEYINPUT30), .ZN(new_n756));
  OR2_X1    g331(.A1(KEYINPUT31), .A2(G11), .ZN(new_n757));
  NAND2_X1  g332(.A1(KEYINPUT31), .A2(G11), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n755), .A2(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT98), .B(KEYINPUT24), .Z(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(G34), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(G34), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n761), .A2(new_n716), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G160), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(new_n728), .ZN(new_n765));
  INV_X1    g340(.A(G2084), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n759), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(new_n766), .B2(new_n765), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n753), .B(new_n768), .C1(new_n741), .C2(new_n739), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n742), .A2(G4), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n622), .B2(new_n742), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G1348), .ZN(new_n772));
  NOR3_X1   g347(.A1(new_n748), .A2(new_n769), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n728), .A2(G33), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT25), .Z(new_n776));
  AOI22_X1  g351(.A1(new_n503), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n776), .B1(new_n463), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n480), .B2(G139), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(KEYINPUT96), .Z(new_n780));
  OAI21_X1  g355(.A(new_n774), .B1(new_n780), .B2(new_n728), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n781), .A2(G2072), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT97), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n781), .A2(G2072), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n637), .A2(new_n638), .A3(new_n717), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n742), .A2(G19), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n562), .B2(new_n742), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(G1341), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n716), .A2(G26), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT28), .Z(new_n790));
  NAND2_X1  g365(.A1(new_n480), .A2(G140), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n482), .A2(G128), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n463), .A2(G116), .ZN(new_n793));
  OAI21_X1  g368(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n791), .B(new_n792), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n790), .B1(new_n795), .B2(G29), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G2067), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n784), .A2(new_n785), .A3(new_n788), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n742), .A2(G20), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT101), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT23), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G299), .B2(G16), .ZN(new_n802));
  INV_X1    g377(.A(G1956), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n798), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n727), .A2(new_n773), .A3(new_n783), .A4(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G6), .B(G305), .S(G16), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT32), .ZN(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT94), .ZN(new_n810));
  XNOR2_X1  g385(.A(G288), .B(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n811), .A2(new_n742), .ZN(new_n812));
  NOR2_X1   g387(.A1(G16), .A2(G23), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT93), .Z(new_n814));
  NOR2_X1   g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT33), .B(G1976), .Z(new_n816));
  AOI22_X1  g391(.A1(new_n809), .A2(new_n703), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n815), .B2(new_n816), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n742), .A2(G22), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT95), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(G166), .B2(new_n742), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(G1971), .Z(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n809), .B2(new_n703), .ZN(new_n823));
  OR3_X1    g398(.A1(new_n818), .A2(new_n823), .A3(KEYINPUT34), .ZN(new_n824));
  OAI21_X1  g399(.A(KEYINPUT34), .B1(new_n818), .B2(new_n823), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n480), .A2(G131), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n482), .A2(G119), .ZN(new_n827));
  OR2_X1    g402(.A1(G95), .A2(G2105), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n828), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT92), .Z(new_n830));
  NAND3_X1  g405(.A1(new_n826), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  MUX2_X1   g406(.A(G25), .B(new_n831), .S(new_n717), .Z(new_n832));
  XOR2_X1   g407(.A(KEYINPUT35), .B(G1991), .Z(new_n833));
  INV_X1    g408(.A(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n832), .B(new_n834), .ZN(new_n835));
  MUX2_X1   g410(.A(G24), .B(G290), .S(G16), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(G1986), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n824), .A2(new_n825), .A3(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n839), .A2(KEYINPUT36), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(KEYINPUT36), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n806), .B1(new_n840), .B2(new_n841), .ZN(G311));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n841), .ZN(new_n843));
  INV_X1    g418(.A(new_n806), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(G150));
  XNOR2_X1  g420(.A(KEYINPUT103), .B(G860), .ZN(new_n846));
  INV_X1    g421(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n622), .A2(G559), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT38), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n850));
  NAND2_X1  g425(.A1(G80), .A2(G543), .ZN(new_n851));
  INV_X1    g426(.A(G67), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n851), .B1(new_n523), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(G651), .ZN(new_n854));
  XNOR2_X1  g429(.A(KEYINPUT102), .B(G93), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n537), .A2(new_n528), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n537), .A2(G55), .A3(G543), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n850), .B(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n849), .B(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n847), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(new_n861), .B2(new_n860), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n858), .A2(new_n847), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT37), .Z(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(G145));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n480), .A2(G142), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n482), .A2(G130), .ZN(new_n869));
  NOR3_X1   g444(.A1(new_n463), .A2(KEYINPUT105), .A3(G118), .ZN(new_n870));
  OAI21_X1  g445(.A(KEYINPUT105), .B1(new_n463), .B2(G118), .ZN(new_n871));
  OAI211_X1 g446(.A(new_n871), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n868), .B(new_n869), .C1(new_n870), .C2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n644), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n831), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n779), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n878));
  AOI211_X1 g453(.A(new_n878), .B(new_n494), .C1(new_n500), .C2(new_n505), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n500), .A2(new_n505), .ZN(new_n880));
  INV_X1    g455(.A(new_n494), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT104), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n795), .B(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n737), .ZN(new_n885));
  AOI21_X1  g460(.A(G2105), .B1(new_n501), .B2(new_n502), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n495), .B1(new_n886), .B2(new_n504), .ZN(new_n887));
  NOR3_X1   g462(.A1(new_n497), .A2(new_n496), .A3(new_n499), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n881), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n878), .ZN(new_n890));
  NAND2_X1  g465(.A1(G164), .A2(KEYINPUT104), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n795), .B(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n738), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n877), .B1(new_n885), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n885), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n876), .B(new_n896), .C1(new_n780), .C2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n639), .A2(G160), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n637), .A2(new_n764), .A3(new_n638), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n899), .A2(G162), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(G162), .B1(new_n899), .B2(new_n900), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n884), .A2(new_n737), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n893), .A2(new_n738), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n904), .A2(new_n905), .A3(new_n780), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n875), .B1(new_n906), .B2(new_n895), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n898), .A2(new_n903), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(G37), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n903), .B1(new_n898), .B2(new_n907), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n867), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n911), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n913), .A2(KEYINPUT40), .A3(new_n909), .A4(new_n908), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n912), .A2(new_n914), .ZN(G395));
  XNOR2_X1  g490(.A(new_n625), .B(new_n859), .ZN(new_n916));
  OAI22_X1  g491(.A1(new_n612), .A2(new_n574), .B1(new_n579), .B2(new_n518), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n917), .A2(G651), .B1(G91), .B2(new_n524), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n918), .A2(new_n573), .B1(new_n611), .B2(new_n616), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n617), .A2(G299), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(KEYINPUT41), .B1(new_n920), .B2(new_n919), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n617), .A2(G299), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT41), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n918), .A2(new_n573), .A3(new_n611), .A4(new_n616), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n922), .A2(new_n923), .A3(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n920), .A2(new_n919), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(KEYINPUT106), .A3(new_n925), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n921), .B1(new_n931), .B2(new_n916), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT42), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n811), .B(G303), .ZN(new_n934));
  XOR2_X1   g509(.A(G290), .B(G305), .Z(new_n935));
  XNOR2_X1  g510(.A(new_n934), .B(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT42), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n937), .B(new_n921), .C1(new_n931), .C2(new_n916), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n933), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n936), .B1(new_n933), .B2(new_n938), .ZN(new_n940));
  OAI21_X1  g515(.A(G868), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G868), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n858), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(G295));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n943), .ZN(G331));
  NAND3_X1  g520(.A1(new_n584), .A2(G168), .A3(new_n586), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n588), .A2(G171), .A3(new_n590), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n562), .B(new_n858), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n859), .A2(new_n946), .A3(new_n947), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n928), .A2(new_n952), .A3(new_n930), .ZN(new_n953));
  INV_X1    g528(.A(new_n936), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n950), .A2(new_n924), .A3(new_n951), .A4(new_n926), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n956), .A2(new_n909), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n953), .A2(new_n955), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(new_n936), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(KEYINPUT43), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n929), .A2(new_n962), .A3(new_n950), .A4(new_n951), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n955), .A2(KEYINPUT107), .ZN(new_n964));
  AOI22_X1  g539(.A1(new_n922), .A2(new_n927), .B1(new_n950), .B2(new_n951), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n936), .B(new_n963), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n956), .A2(new_n966), .A3(new_n909), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n960), .A2(new_n961), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT43), .B1(new_n958), .B2(new_n936), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n961), .B1(new_n957), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n973));
  AOI21_X1  g548(.A(KEYINPUT108), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n959), .A2(new_n968), .A3(new_n909), .A4(new_n956), .ZN(new_n975));
  AND4_X1   g550(.A1(KEYINPUT108), .A2(new_n973), .A3(new_n975), .A4(KEYINPUT44), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n970), .B1(new_n974), .B2(new_n976), .ZN(G397));
  OAI21_X1  g552(.A(KEYINPUT109), .B1(new_n892), .B2(G1384), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n979));
  INV_X1    g554(.A(G1384), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n883), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  INV_X1    g557(.A(G125), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n983), .B1(new_n501), .B2(new_n502), .ZN(new_n984));
  INV_X1    g559(.A(new_n467), .ZN(new_n985));
  OAI21_X1  g560(.A(G2105), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n476), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n986), .A2(G40), .A3(new_n987), .A4(new_n469), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n978), .A2(new_n981), .A3(new_n982), .A4(new_n989), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n990), .A2(G1986), .A3(G290), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT48), .ZN(new_n992));
  XOR2_X1   g567(.A(new_n795), .B(G2067), .Z(new_n993));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n994));
  OR3_X1    g569(.A1(new_n993), .A2(new_n994), .A3(new_n990), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n994), .B1(new_n993), .B2(new_n990), .ZN(new_n996));
  INV_X1    g571(.A(new_n990), .ZN(new_n997));
  XNOR2_X1  g572(.A(new_n737), .B(G1996), .ZN(new_n998));
  AOI22_X1  g573(.A1(new_n995), .A2(new_n996), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n831), .A2(new_n834), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n831), .A2(new_n834), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n997), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT127), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n999), .A2(KEYINPUT127), .A3(new_n1002), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n992), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n795), .A2(G2067), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1008), .B1(new_n999), .B2(new_n1001), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n990), .B1(new_n993), .B2(new_n738), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT46), .B1(new_n990), .B2(G1996), .ZN(new_n1011));
  OR3_X1    g586(.A1(new_n990), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  OAI22_X1  g591(.A1(new_n1009), .A2(new_n990), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1007), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(G303), .A2(G8), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1019), .B(KEYINPUT55), .ZN(new_n1020));
  NOR2_X1   g595(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n988), .B1(new_n889), .B2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(G2090), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT111), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n889), .A2(new_n980), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1026), .B1(new_n1027), .B2(new_n982), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1026), .B(new_n982), .C1(G164), .C2(G1384), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n989), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n982), .A2(G1384), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT112), .B1(new_n883), .B2(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n890), .A2(KEYINPUT112), .A3(new_n891), .A4(new_n1032), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1031), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT113), .B(G1971), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1025), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g613(.A(KEYINPUT114), .B(G8), .Z(new_n1039));
  OAI21_X1  g614(.A(new_n1020), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1020), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1037), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n890), .A2(new_n891), .A3(new_n1032), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT112), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n1034), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1042), .B1(new_n1046), .B2(new_n1031), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1041), .B(G8), .C1(new_n1047), .C2(new_n1025), .ZN(new_n1048));
  XNOR2_X1  g623(.A(G305), .B(new_n703), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(KEYINPUT49), .ZN(new_n1050));
  XNOR2_X1  g625(.A(G305), .B(G1981), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT49), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(G164), .A2(G1384), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1039), .B1(new_n1054), .B2(new_n989), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1050), .A2(new_n1053), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT116), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1050), .A2(new_n1053), .A3(KEYINPUT116), .A4(new_n1055), .ZN(new_n1059));
  INV_X1    g634(.A(G1976), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1055), .B1(new_n811), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT52), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(KEYINPUT115), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  OR2_X1    g639(.A1(new_n1061), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(KEYINPUT52), .A2(G1976), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1061), .A2(new_n1064), .B1(G288), .B2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1058), .A2(new_n1059), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1039), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1022), .A2(new_n766), .A3(new_n1023), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n988), .B1(new_n889), .B2(new_n1032), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n982), .B1(G164), .B2(G1384), .ZN(new_n1072));
  AOI21_X1  g647(.A(G1966), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1069), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1074), .A2(G286), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1040), .A2(new_n1048), .A3(new_n1068), .A4(new_n1075), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT117), .B(KEYINPUT63), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G8), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1020), .B1(new_n1038), .B2(new_n1079), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1075), .A2(KEYINPUT63), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1080), .A2(new_n1048), .A3(new_n1068), .A4(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1078), .A2(new_n1082), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1040), .A2(new_n1048), .A3(new_n1068), .ZN(new_n1084));
  INV_X1    g659(.A(G1966), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1072), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1032), .ZN(new_n1087));
  OAI211_X1 g662(.A(G160), .B(G40), .C1(G164), .C2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1085), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1022), .A2(new_n766), .A3(new_n1023), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1079), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(G168), .A2(new_n1039), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT51), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1039), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT51), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(G168), .B2(new_n1039), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT121), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1096), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1074), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1093), .A2(new_n1097), .A3(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1092), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(KEYINPUT62), .ZN(new_n1104));
  INV_X1    g679(.A(G2078), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1046), .A2(new_n1105), .A3(new_n1031), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(KEYINPUT122), .B(G1961), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1024), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1107), .A2(G2078), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1071), .A2(new_n1072), .A3(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(G301), .B1(new_n1108), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT62), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1101), .A2(new_n1116), .A3(new_n1102), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1084), .A2(new_n1104), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1119));
  OR2_X1    g694(.A1(G288), .A2(G1976), .ZN(new_n1120));
  OAI22_X1  g695(.A1(new_n1119), .A2(new_n1120), .B1(G1981), .B2(G305), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1048), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1121), .A2(new_n1055), .B1(new_n1122), .B2(new_n1068), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1083), .A2(new_n1118), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1084), .A2(new_n1103), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n1126));
  XNOR2_X1  g701(.A(G299), .B(KEYINPUT57), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1024), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1128), .A2(G1956), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1072), .A2(KEYINPUT111), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1131), .A2(new_n989), .A3(new_n1029), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1132), .B1(new_n1045), .B2(new_n1034), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT56), .B(G2072), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1126), .B1(new_n1130), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1129), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1127), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1054), .A2(new_n989), .ZN(new_n1140));
  OR3_X1    g715(.A1(new_n1140), .A2(KEYINPUT118), .A3(G2067), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT118), .B1(new_n1140), .B2(G2067), .ZN(new_n1142));
  INV_X1    g717(.A(G1348), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1024), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1141), .A2(KEYINPUT60), .A3(new_n1142), .A4(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(new_n622), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n1142), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT60), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1136), .A2(new_n1139), .B1(new_n1146), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1130), .A2(new_n1135), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1139), .A2(new_n1152), .ZN(new_n1153));
  XOR2_X1   g728(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  XOR2_X1   g730(.A(KEYINPUT119), .B(G1996), .Z(new_n1156));
  XOR2_X1   g731(.A(KEYINPUT58), .B(G1341), .Z(new_n1157));
  AOI22_X1  g732(.A1(new_n1133), .A2(new_n1156), .B1(new_n1140), .B2(new_n1157), .ZN(new_n1158));
  OR3_X1    g733(.A1(new_n1158), .A2(KEYINPUT59), .A3(new_n850), .ZN(new_n1159));
  OAI21_X1  g734(.A(KEYINPUT59), .B1(new_n1158), .B2(new_n850), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1151), .A2(new_n1155), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1139), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n617), .B1(new_n1147), .B2(new_n1142), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1152), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1125), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT53), .B1(new_n1133), .B2(new_n1105), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1114), .A2(G301), .ZN(new_n1168));
  OAI21_X1  g743(.A(KEYINPUT124), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1108), .A2(new_n1170), .A3(G301), .A4(new_n1114), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT54), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1111), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n978), .A2(new_n982), .A3(new_n981), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n989), .A2(new_n1112), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1176), .B1(new_n1045), .B2(new_n1034), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1174), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1108), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1173), .B1(new_n1179), .B2(G171), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1172), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT125), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1172), .A2(new_n1180), .A3(KEYINPUT125), .ZN(new_n1184));
  AND3_X1   g759(.A1(new_n1108), .A2(new_n1178), .A3(G301), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1173), .B1(new_n1185), .B2(new_n1115), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(KEYINPUT123), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT123), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1188), .B(new_n1173), .C1(new_n1185), .C2(new_n1115), .ZN(new_n1189));
  AOI22_X1  g764(.A1(new_n1183), .A2(new_n1184), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1124), .B1(new_n1166), .B2(new_n1190), .ZN(new_n1191));
  XNOR2_X1  g766(.A(G290), .B(new_n705), .ZN(new_n1192));
  OAI211_X1 g767(.A(new_n999), .B(new_n1002), .C1(new_n990), .C2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1018), .B1(new_n1191), .B2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g769(.A1(new_n960), .A2(new_n969), .ZN(new_n1196));
  NAND3_X1  g770(.A1(new_n913), .A2(new_n909), .A3(new_n908), .ZN(new_n1197));
  OR3_X1    g771(.A1(G401), .A2(new_n461), .A3(G227), .ZN(new_n1198));
  AOI21_X1  g772(.A(new_n1198), .B1(new_n711), .B2(new_n714), .ZN(new_n1199));
  AND3_X1   g773(.A1(new_n1196), .A2(new_n1197), .A3(new_n1199), .ZN(G308));
  NAND3_X1  g774(.A1(new_n1196), .A2(new_n1197), .A3(new_n1199), .ZN(G225));
endmodule


