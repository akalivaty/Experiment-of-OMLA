//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:42 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n456, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT64), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  AOI22_X1  g029(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(G319));
  NAND2_X1  g030(.A1(G113), .A2(G2104), .ZN(new_n456));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2104), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n456), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g038(.A(KEYINPUT65), .B(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g040(.A(KEYINPUT66), .B(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n458), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n470), .B1(new_n466), .B2(KEYINPUT3), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT65), .A2(G2105), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT65), .A2(G2105), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n471), .A2(G137), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n469), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n459), .A2(KEYINPUT66), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G2104), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n478), .A2(new_n480), .A3(KEYINPUT3), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(new_n458), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n482), .A2(new_n474), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OAI221_X1 g061(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n474), .C2(G112), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND4_X1  g064(.A1(new_n481), .A2(G138), .A3(new_n474), .A4(new_n458), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n464), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  AND3_X1   g068(.A1(new_n458), .A2(new_n460), .A3(new_n493), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n490), .A2(KEYINPUT4), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g070(.A1(G126), .A2(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n481), .A2(new_n458), .A3(new_n496), .ZN(new_n497));
  OR2_X1    g072(.A1(G102), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n498), .B(G2104), .C1(G114), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT67), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n497), .A2(new_n503), .A3(new_n500), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n495), .B1(new_n502), .B2(new_n504), .ZN(G164));
  NAND2_X1  g080(.A1(G75), .A2(G543), .ZN(new_n506));
  AND3_X1   g081(.A1(KEYINPUT68), .A2(KEYINPUT5), .A3(G543), .ZN(new_n507));
  AOI21_X1  g082(.A(G543), .B1(KEYINPUT68), .B2(KEYINPUT5), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G62), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n511), .A2(G651), .B1(G50), .B2(new_n516), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n507), .A2(new_n508), .B1(new_n512), .B2(new_n513), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT69), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT68), .A2(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(new_n515), .ZN(new_n522));
  NAND3_X1  g097(.A1(KEYINPUT68), .A2(KEYINPUT5), .A3(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT6), .B(G651), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n524), .A2(KEYINPUT69), .A3(new_n525), .ZN(new_n526));
  XOR2_X1   g101(.A(KEYINPUT70), .B(G88), .Z(new_n527));
  NAND3_X1  g102(.A1(new_n520), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n517), .A2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  AND2_X1   g105(.A1(new_n520), .A2(new_n526), .ZN(new_n531));
  XOR2_X1   g106(.A(KEYINPUT71), .B(G89), .Z(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT72), .ZN(new_n534));
  NAND3_X1  g109(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  AND2_X1   g112(.A1(G63), .A2(G651), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n516), .A2(G51), .B1(new_n524), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n534), .B1(new_n533), .B2(new_n536), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(G168));
  NAND2_X1  g117(.A1(new_n531), .A2(G90), .ZN(new_n543));
  INV_X1    g118(.A(G64), .ZN(new_n544));
  INV_X1    g119(.A(G77), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n509), .A2(new_n544), .B1(new_n545), .B2(new_n515), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI221_X1 g123(.A(KEYINPUT73), .B1(new_n545), .B2(new_n515), .C1(new_n509), .C2(new_n544), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n548), .A2(G651), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n516), .A2(G52), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n543), .A2(new_n550), .A3(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  NAND2_X1  g128(.A1(new_n531), .A2(G81), .ZN(new_n554));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G56), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n509), .B2(new_n556), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n557), .A2(G651), .B1(G43), .B2(new_n516), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  INV_X1    g141(.A(G78), .ZN(new_n567));
  OAI22_X1  g142(.A1(new_n509), .A2(new_n566), .B1(new_n567), .B2(new_n515), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT74), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT74), .ZN(new_n570));
  OAI221_X1 g145(.A(new_n570), .B1(new_n567), .B2(new_n515), .C1(new_n509), .C2(new_n566), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(G651), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n520), .A2(G91), .A3(new_n526), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n525), .A2(G53), .A3(G543), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT9), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n572), .A2(new_n573), .A3(new_n575), .ZN(G299));
  INV_X1    g151(.A(G168), .ZN(G286));
  INV_X1    g152(.A(G74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n509), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(G651), .A2(new_n579), .B1(new_n516), .B2(G49), .ZN(new_n580));
  INV_X1    g155(.A(G87), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n520), .A2(new_n526), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(G288));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n584));
  OAI21_X1  g159(.A(G61), .B1(new_n507), .B2(new_n508), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n584), .B1(new_n587), .B2(G651), .ZN(new_n588));
  INV_X1    g163(.A(G651), .ZN(new_n589));
  AOI211_X1 g164(.A(KEYINPUT75), .B(new_n589), .C1(new_n585), .C2(new_n586), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n516), .A2(G48), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n520), .A2(G86), .A3(new_n526), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT76), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n591), .A2(KEYINPUT76), .A3(new_n592), .A4(new_n593), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n524), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n589), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n600), .A2(KEYINPUT77), .B1(G47), .B2(new_n516), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n531), .A2(G85), .ZN(new_n602));
  OAI211_X1 g177(.A(new_n601), .B(new_n602), .C1(KEYINPUT77), .C2(new_n600), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n516), .A2(G54), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n524), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(new_n589), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n531), .A2(KEYINPUT10), .A3(G92), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n582), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n607), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n604), .B1(G868), .B2(new_n612), .ZN(G284));
  OAI21_X1  g188(.A(new_n604), .B1(G868), .B2(new_n612), .ZN(G321));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  NAND2_X1  g190(.A1(G299), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G168), .B2(new_n615), .ZN(G297));
  OAI21_X1  g192(.A(new_n616), .B1(G168), .B2(new_n615), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(G148));
  OAI21_X1  g195(.A(KEYINPUT78), .B1(new_n560), .B2(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n612), .A2(new_n619), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  MUX2_X1   g198(.A(KEYINPUT78), .B(new_n621), .S(new_n623), .Z(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g200(.A1(new_n467), .A2(new_n458), .A3(new_n460), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2100), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n483), .A2(G135), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT79), .ZN(new_n631));
  OAI221_X1 g206(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n474), .C2(G111), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n485), .A2(G123), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n634), .A2(G2096), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(G2096), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n629), .A2(new_n635), .A3(new_n636), .ZN(G156));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT81), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2427), .B(G2430), .Z(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n649), .B(new_n650), .Z(new_n651));
  OR2_X1    g226(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n648), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(G401));
  XNOR2_X1  g230(.A(G2072), .B(G2078), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT17), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NOR3_X1   g235(.A1(new_n657), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT82), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n657), .A2(new_n658), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n663), .B(new_n660), .C1(new_n656), .C2(new_n658), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n659), .A2(new_n656), .A3(new_n658), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT18), .Z(new_n666));
  NAND3_X1  g241(.A1(new_n662), .A2(new_n664), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2096), .B(G2100), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n669), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n676), .A2(KEYINPUT83), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(KEYINPUT83), .ZN(new_n678));
  XOR2_X1   g253(.A(G1971), .B(G1976), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n677), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n681), .A2(KEYINPUT84), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(KEYINPUT84), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT20), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n682), .A2(KEYINPUT20), .A3(new_n683), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n673), .A2(new_n674), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n680), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT85), .Z(new_n690));
  NOR3_X1   g265(.A1(new_n680), .A2(new_n676), .A3(new_n688), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n686), .A2(new_n687), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND4_X1  g271(.A1(new_n686), .A2(new_n687), .A3(new_n692), .A4(new_n694), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1991), .B(G1996), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n699), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n696), .A2(new_n701), .A3(new_n697), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1981), .B(G1986), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n703), .B(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(G229));
  NAND2_X1  g282(.A1(new_n485), .A2(G129), .ZN(new_n708));
  NAND3_X1  g283(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT26), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(KEYINPUT97), .B1(new_n467), .B2(G105), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n467), .A2(KEYINPUT97), .A3(G105), .ZN(new_n715));
  AOI22_X1  g290(.A1(new_n714), .A2(new_n715), .B1(G141), .B2(new_n483), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G29), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G32), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n721), .A2(KEYINPUT27), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(KEYINPUT27), .ZN(new_n723));
  INV_X1    g298(.A(G1996), .ZN(new_n724));
  OR3_X1    g299(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n719), .A2(G35), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G162), .B2(new_n719), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT29), .Z(new_n728));
  INV_X1    g303(.A(G2090), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n724), .B1(new_n722), .B2(new_n723), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n725), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G4), .A2(G16), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n612), .B2(G16), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n734), .B(G1348), .ZN(new_n735));
  INV_X1    g310(.A(G16), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G20), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT23), .Z(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G299), .B2(G16), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G1956), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n728), .B2(new_n729), .ZN(new_n741));
  NOR3_X1   g316(.A1(new_n732), .A2(new_n735), .A3(new_n741), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT93), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n719), .A2(G26), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n744), .B(new_n745), .Z(new_n746));
  NAND3_X1  g321(.A1(new_n471), .A2(G140), .A3(new_n499), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n471), .A2(G128), .A3(new_n464), .ZN(new_n748));
  OAI221_X1 g323(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n474), .C2(G116), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n746), .B1(new_n719), .B2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G2067), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n719), .A2(G27), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(G164), .B2(new_n719), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(G2078), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(G2078), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n754), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(G16), .A2(G19), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n560), .B2(G16), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(G1341), .Z(new_n762));
  INV_X1    g337(.A(G34), .ZN(new_n763));
  AOI21_X1  g338(.A(G29), .B1(new_n763), .B2(KEYINPUT24), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(KEYINPUT24), .B2(new_n763), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n476), .B2(new_n719), .ZN(new_n766));
  INV_X1    g341(.A(G2084), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G28), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n769), .A2(KEYINPUT30), .ZN(new_n770));
  AOI21_X1  g345(.A(G29), .B1(new_n769), .B2(KEYINPUT30), .ZN(new_n771));
  OR2_X1    g346(.A1(KEYINPUT31), .A2(G11), .ZN(new_n772));
  NAND2_X1  g347(.A1(KEYINPUT31), .A2(G11), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n770), .A2(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n634), .B2(new_n719), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n768), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n736), .A2(G5), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G171), .B2(new_n736), .ZN(new_n778));
  INV_X1    g353(.A(G1961), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n762), .A2(new_n776), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n719), .A2(G33), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n471), .A2(G139), .A3(new_n499), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT94), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT95), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT25), .ZN(new_n786));
  NAND2_X1  g361(.A1(G103), .A2(G2104), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n464), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n474), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n789));
  NAND2_X1  g364(.A1(G115), .A2(G2104), .ZN(new_n790));
  INV_X1    g365(.A(G127), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n461), .B2(new_n791), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n788), .A2(new_n789), .B1(new_n792), .B2(new_n464), .ZN(new_n793));
  AND3_X1   g368(.A1(new_n784), .A2(new_n785), .A3(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n785), .B1(new_n784), .B2(new_n793), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n782), .B1(new_n796), .B2(new_n719), .ZN(new_n797));
  AOI211_X1 g372(.A(new_n759), .B(new_n781), .C1(G2072), .C2(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT99), .B(G1966), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(KEYINPUT100), .ZN(new_n801));
  NAND2_X1  g376(.A1(G168), .A2(G16), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(KEYINPUT98), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n802), .B(KEYINPUT98), .C1(G16), .C2(G21), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n800), .A2(KEYINPUT100), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n797), .A2(G2072), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT96), .Z(new_n809));
  NAND4_X1  g384(.A1(new_n742), .A2(new_n798), .A3(new_n807), .A4(new_n809), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n596), .A2(G16), .A3(new_n597), .ZN(new_n811));
  OR2_X1    g386(.A1(G6), .A2(G16), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT32), .B(G1981), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n517), .A2(G16), .A3(new_n528), .ZN(new_n817));
  OR2_X1    g392(.A1(G16), .A2(G22), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT89), .B(G1971), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n817), .A2(new_n818), .A3(new_n820), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT90), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n826));
  XOR2_X1   g401(.A(KEYINPUT33), .B(G1976), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n531), .A2(G87), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n736), .B1(new_n828), .B2(new_n580), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n736), .A2(G23), .ZN(new_n830));
  NOR3_X1   g405(.A1(new_n829), .A2(KEYINPUT88), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n830), .B1(G288), .B2(G16), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT88), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n827), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(KEYINPUT88), .B1(new_n829), .B2(new_n830), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n832), .A2(new_n833), .ZN(new_n837));
  INV_X1    g412(.A(new_n827), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n816), .A2(new_n825), .A3(new_n826), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(KEYINPUT34), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT91), .ZN(new_n843));
  AND2_X1   g418(.A1(new_n825), .A2(new_n840), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT34), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n844), .A2(new_n845), .A3(new_n816), .A4(new_n826), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT35), .B(G1991), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n719), .A2(G25), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT86), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n483), .A2(G131), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n485), .A2(G119), .ZN(new_n851));
  OAI221_X1 g426(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n474), .C2(G107), .ZN(new_n852));
  NAND3_X1  g427(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(KEYINPUT87), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n854), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n847), .B(new_n849), .C1(new_n857), .C2(new_n719), .ZN(new_n858));
  NAND2_X1  g433(.A1(G290), .A2(G16), .ZN(new_n859));
  INV_X1    g434(.A(G24), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n859), .B1(G16), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(G1986), .ZN(new_n862));
  INV_X1    g437(.A(new_n847), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n719), .B1(new_n855), .B2(new_n856), .ZN(new_n864));
  INV_X1    g439(.A(new_n849), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(G1986), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n859), .B(new_n867), .C1(G16), .C2(new_n860), .ZN(new_n868));
  AND4_X1   g443(.A1(new_n858), .A2(new_n862), .A3(new_n866), .A4(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n843), .B1(new_n846), .B2(new_n869), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n869), .B(new_n843), .C1(new_n841), .C2(KEYINPUT34), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n842), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT36), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT36), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n875), .B(new_n842), .C1(new_n870), .C2(new_n872), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n810), .B1(new_n874), .B2(new_n876), .ZN(G311));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n876), .ZN(new_n878));
  INV_X1    g453(.A(new_n810), .ZN(new_n879));
  AOI21_X1  g454(.A(KEYINPUT101), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT101), .ZN(new_n881));
  AOI211_X1 g456(.A(new_n881), .B(new_n810), .C1(new_n874), .C2(new_n876), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n880), .A2(new_n882), .ZN(G150));
  NAND2_X1  g458(.A1(new_n516), .A2(G55), .ZN(new_n884));
  AOI22_X1  g459(.A1(new_n524), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n885));
  INV_X1    g460(.A(G93), .ZN(new_n886));
  OAI221_X1 g461(.A(new_n884), .B1(new_n589), .B2(new_n885), .C1(new_n582), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(G860), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT104), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT37), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n612), .A2(G559), .ZN(new_n891));
  XOR2_X1   g466(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  AND2_X1   g468(.A1(new_n559), .A2(new_n887), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n559), .A2(new_n887), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n893), .B(new_n897), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n898), .A2(KEYINPUT39), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n899), .B(KEYINPUT103), .Z(new_n900));
  INV_X1    g475(.A(G860), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n898), .B2(KEYINPUT39), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n890), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n903), .B(new_n904), .ZN(G145));
  NAND2_X1  g480(.A1(new_n483), .A2(G142), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n485), .A2(G130), .ZN(new_n907));
  OAI221_X1 g482(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n474), .C2(G118), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n627), .B(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n751), .B1(new_n495), .B2(new_n501), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n483), .A2(G141), .ZN(new_n913));
  INV_X1    g488(.A(new_n715), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n913), .B1(new_n914), .B2(new_n713), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n915), .A2(new_n711), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n492), .A2(new_n494), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n501), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n750), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n912), .A2(new_n916), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n916), .B1(new_n912), .B2(new_n921), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n796), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n912), .A2(new_n921), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n717), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n784), .A2(new_n793), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n912), .A2(new_n916), .A3(new_n921), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n924), .A2(new_n929), .A3(KEYINPUT106), .ZN(new_n930));
  INV_X1    g505(.A(new_n857), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n926), .A2(new_n932), .A3(new_n927), .A4(new_n928), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n931), .B1(new_n930), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n911), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n930), .A2(new_n933), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(new_n857), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n910), .A3(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n476), .B(new_n488), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(new_n634), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n936), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(G37), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n942), .B1(new_n936), .B2(new_n940), .ZN(new_n946));
  OAI21_X1  g521(.A(KEYINPUT107), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n936), .A2(new_n940), .ZN(new_n948));
  INV_X1    g523(.A(new_n942), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n950), .A2(new_n951), .A3(new_n944), .A4(new_n943), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n947), .A2(KEYINPUT40), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT40), .B1(new_n947), .B2(new_n952), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(G395));
  NAND2_X1  g530(.A1(new_n887), .A2(new_n615), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n612), .B(G299), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n957), .B(KEYINPUT41), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n896), .B(new_n622), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n960), .B1(new_n957), .B2(new_n959), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n961), .B(KEYINPUT42), .ZN(new_n962));
  INV_X1    g537(.A(G288), .ZN(new_n963));
  NAND2_X1  g538(.A1(G305), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n596), .A2(G288), .A3(new_n597), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(G290), .B(G303), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n964), .A2(new_n967), .A3(new_n965), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n962), .B(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n956), .B1(new_n973), .B2(new_n615), .ZN(G295));
  OAI21_X1  g549(.A(new_n956), .B1(new_n973), .B2(new_n615), .ZN(G331));
  INV_X1    g550(.A(new_n541), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n976), .A2(G171), .A3(new_n537), .A4(new_n539), .ZN(new_n977));
  OAI21_X1  g552(.A(G301), .B1(new_n540), .B2(new_n541), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n896), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n896), .A2(new_n978), .A3(new_n977), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT108), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n896), .A2(new_n978), .A3(new_n977), .A4(KEYINPUT108), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n979), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n984), .A2(new_n958), .ZN(new_n985));
  INV_X1    g560(.A(new_n957), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n979), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n980), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n971), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n971), .B(new_n988), .C1(new_n984), .C2(new_n958), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(new_n944), .ZN(new_n991));
  OR3_X1    g566(.A1(new_n989), .A2(new_n991), .A3(KEYINPUT43), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT43), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT109), .ZN(new_n994));
  INV_X1    g569(.A(new_n980), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n995), .A2(new_n979), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n994), .B1(new_n996), .B2(new_n958), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT41), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n957), .B(new_n998), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n999), .B(KEYINPUT109), .C1(new_n979), .C2(new_n995), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n982), .A2(new_n983), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n987), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n997), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n991), .B1(new_n972), .B2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n992), .B(KEYINPUT44), .C1(new_n993), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1003), .A2(new_n972), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1007), .A2(new_n993), .A3(new_n944), .A4(new_n990), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT43), .B1(new_n989), .B2(new_n991), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1006), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI211_X1 g587(.A(KEYINPUT110), .B(KEYINPUT44), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1005), .B1(new_n1012), .B2(new_n1013), .ZN(G397));
  AOI21_X1  g589(.A(G1384), .B1(new_n919), .B2(new_n920), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  XNOR2_X1  g592(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n1018));
  INV_X1    g593(.A(G1384), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(new_n495), .B2(new_n501), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT111), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1017), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n475), .A2(new_n465), .A3(G40), .A4(new_n468), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n750), .B(G2067), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1026), .B(KEYINPUT113), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1025), .B1(new_n1027), .B2(new_n916), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1028), .B(KEYINPUT125), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1024), .A2(new_n724), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1030), .B(KEYINPUT46), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1032), .B(KEYINPUT47), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n931), .A2(new_n863), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n916), .B(G1996), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n857), .A2(new_n847), .ZN(new_n1036));
  AND4_X1   g611(.A1(new_n1027), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1037), .A2(new_n1025), .ZN(new_n1038));
  NOR2_X1   g613(.A1(G290), .A2(G1986), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1025), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1038), .B1(KEYINPUT48), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1042), .B1(KEYINPUT48), .B2(new_n1041), .ZN(new_n1043));
  AND4_X1   g618(.A1(new_n847), .A2(new_n1027), .A3(new_n857), .A4(new_n1035), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n750), .A2(G2067), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1024), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AND3_X1   g621(.A1(new_n1033), .A2(new_n1043), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT118), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT50), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n497), .A2(new_n503), .A3(new_n500), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n503), .B1(new_n497), .B2(new_n500), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n493), .B1(new_n471), .B2(new_n492), .ZN(new_n1052));
  AND2_X1   g627(.A1(new_n492), .A2(new_n494), .ZN(new_n1053));
  OAI22_X1  g628(.A1(new_n1050), .A2(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1049), .B1(new_n1054), .B2(new_n1019), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1049), .B(new_n1019), .C1(new_n495), .C2(new_n501), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1023), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n767), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n1055), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT45), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1023), .B1(new_n1020), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1018), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1054), .A2(new_n1019), .A3(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n800), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(G8), .B(G168), .C1(new_n1060), .C2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT63), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NOR4_X1   g643(.A1(new_n1055), .A2(new_n1057), .A3(G2090), .A4(new_n1023), .ZN(new_n1069));
  XOR2_X1   g644(.A(KEYINPUT114), .B(G1971), .Z(new_n1070));
  OAI211_X1 g645(.A(KEYINPUT45), .B(new_n1019), .C1(new_n495), .C2(new_n501), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1071), .A2(new_n1058), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1018), .B1(G164), .B2(G1384), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1070), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g649(.A(G8), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT55), .ZN(new_n1076));
  INV_X1    g651(.A(G8), .ZN(new_n1077));
  NOR3_X1   g652(.A1(G166), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1075), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1068), .A2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n580), .B(G1976), .C1(new_n581), .C2(new_n582), .ZN(new_n1084));
  OAI211_X1 g659(.A(G8), .B(new_n1084), .C1(new_n1020), .C2(new_n1023), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT52), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT52), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n963), .B2(G1976), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1086), .B1(new_n1088), .B2(new_n1085), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n520), .A2(G86), .A3(new_n526), .ZN(new_n1090));
  INV_X1    g665(.A(G61), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n522), .B2(new_n523), .ZN(new_n1092));
  INV_X1    g667(.A(new_n586), .ZN(new_n1093));
  OAI21_X1  g668(.A(G651), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(new_n592), .ZN(new_n1095));
  OAI21_X1  g670(.A(G1981), .B1(new_n1090), .B2(new_n1095), .ZN(new_n1096));
  XOR2_X1   g671(.A(KEYINPUT115), .B(G1981), .Z(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n516), .B2(G48), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n593), .B(new_n1098), .C1(new_n588), .C2(new_n590), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT49), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1096), .A2(new_n1099), .A3(KEYINPUT49), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1077), .B1(new_n1015), .B2(new_n1058), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT116), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1102), .A2(KEYINPUT116), .A3(new_n1104), .A4(new_n1103), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1089), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g684(.A(G8), .B(new_n1080), .C1(new_n1069), .C2(new_n1074), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1048), .B1(new_n1083), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1089), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1113), .A2(new_n1110), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n799), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1118), .A2(new_n767), .A3(new_n1058), .A4(new_n1056), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1120), .A2(KEYINPUT63), .A3(G8), .A4(G168), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1118), .A2(new_n729), .A3(new_n1058), .A4(new_n1056), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1070), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1063), .B1(new_n1054), .B2(new_n1019), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1071), .A2(new_n1058), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1122), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1080), .B1(new_n1127), .B2(G8), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1121), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1115), .A2(new_n1129), .A3(KEYINPUT118), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1023), .B1(new_n1020), .B2(KEYINPUT50), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1054), .A2(new_n1049), .A3(new_n1019), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1131), .A2(new_n1132), .A3(new_n729), .ZN(new_n1133));
  OAI21_X1  g708(.A(G8), .B1(new_n1074), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n1081), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1066), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1135), .A2(new_n1109), .A3(new_n1110), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(new_n1067), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1112), .A2(new_n1130), .A3(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1113), .ZN(new_n1140));
  NOR3_X1   g715(.A1(new_n1140), .A2(new_n1110), .A3(new_n1089), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1099), .B(KEYINPUT117), .ZN(new_n1142));
  OR2_X1    g717(.A1(G288), .A2(G1976), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1142), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1141), .B1(new_n1104), .B2(new_n1144), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1139), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1147));
  INV_X1    g722(.A(G1956), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT57), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(KEYINPUT119), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n572), .A2(new_n573), .A3(new_n575), .A4(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1150), .A2(KEYINPUT119), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1152), .B(new_n1154), .ZN(new_n1155));
  XNOR2_X1  g730(.A(KEYINPUT56), .B(G2072), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1072), .A2(new_n1073), .A3(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1149), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n612), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n502), .A2(new_n504), .ZN(new_n1160));
  AOI21_X1  g735(.A(G1384), .B1(new_n1160), .B2(new_n919), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1058), .B(new_n1056), .C1(new_n1161), .C2(new_n1049), .ZN(new_n1162));
  INV_X1    g737(.A(G1348), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1015), .A2(new_n1058), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1165), .A2(G2067), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1159), .B1(new_n1164), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1155), .B1(new_n1149), .B2(new_n1157), .ZN(new_n1169));
  OAI211_X1 g744(.A(KEYINPUT120), .B(new_n1158), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1152), .B(new_n1153), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1156), .ZN(new_n1173));
  NOR3_X1   g748(.A1(new_n1124), .A2(new_n1125), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(G1956), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1172), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1166), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1176), .B1(new_n1159), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT120), .B1(new_n1178), .B2(new_n1158), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1171), .A2(new_n1179), .ZN(new_n1180));
  XOR2_X1   g755(.A(KEYINPUT58), .B(G1341), .Z(new_n1181));
  NAND2_X1  g756(.A1(new_n1165), .A2(new_n1181), .ZN(new_n1182));
  NOR3_X1   g757(.A1(new_n1124), .A2(new_n1125), .A3(G1996), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1182), .B1(new_n1183), .B2(KEYINPUT121), .ZN(new_n1184));
  AND4_X1   g759(.A1(KEYINPUT121), .A2(new_n1072), .A3(new_n1073), .A4(new_n724), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n560), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT59), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  OAI211_X1 g763(.A(KEYINPUT59), .B(new_n560), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n1190));
  AND3_X1   g765(.A1(new_n1158), .A2(new_n1176), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1190), .B1(new_n1158), .B2(new_n1176), .ZN(new_n1192));
  OAI211_X1 g767(.A(new_n1188), .B(new_n1189), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1193));
  AND2_X1   g768(.A1(new_n1177), .A2(KEYINPUT60), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n612), .B1(new_n1177), .B2(KEYINPUT60), .ZN(new_n1195));
  XNOR2_X1  g770(.A(new_n1194), .B(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1180), .B1(new_n1193), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT51), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1117), .A2(G168), .A3(new_n1119), .ZN(new_n1199));
  NAND2_X1  g774(.A1(KEYINPUT122), .A2(G8), .ZN(new_n1200));
  INV_X1    g775(.A(new_n1200), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1198), .B1(new_n1199), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g777(.A(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1199), .A2(new_n1198), .A3(new_n1201), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1120), .A2(G8), .A3(G286), .ZN(new_n1205));
  NAND3_X1  g780(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  INV_X1    g781(.A(KEYINPUT54), .ZN(new_n1207));
  INV_X1    g782(.A(G2078), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1072), .A2(new_n1073), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT53), .ZN(new_n1210));
  AOI22_X1  g785(.A1(new_n1209), .A2(new_n1210), .B1(new_n1162), .B2(new_n779), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1210), .A2(G2078), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1062), .A2(new_n1064), .A3(new_n1212), .ZN(new_n1213));
  AOI21_X1  g788(.A(G301), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g789(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1162), .A2(new_n779), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1022), .A2(new_n1072), .A3(new_n1212), .ZN(new_n1217));
  AND4_X1   g792(.A1(G301), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1207), .B1(new_n1214), .B2(new_n1218), .ZN(new_n1219));
  AND3_X1   g794(.A1(new_n1135), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1221), .A2(G171), .ZN(new_n1222));
  NAND3_X1  g797(.A1(new_n1211), .A2(G301), .A3(new_n1213), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1222), .A2(KEYINPUT54), .A3(new_n1223), .ZN(new_n1224));
  AND4_X1   g799(.A1(new_n1206), .A2(new_n1219), .A3(new_n1220), .A4(new_n1224), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1197), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g801(.A(KEYINPUT123), .ZN(new_n1227));
  INV_X1    g802(.A(new_n1204), .ZN(new_n1228));
  INV_X1    g803(.A(new_n1205), .ZN(new_n1229));
  NOR3_X1   g804(.A1(new_n1228), .A2(new_n1229), .A3(new_n1202), .ZN(new_n1230));
  INV_X1    g805(.A(KEYINPUT62), .ZN(new_n1231));
  OAI21_X1  g806(.A(new_n1227), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  NAND4_X1  g807(.A1(new_n1214), .A2(new_n1135), .A3(new_n1110), .A4(new_n1109), .ZN(new_n1233));
  AOI21_X1  g808(.A(new_n1233), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1234));
  NAND3_X1  g809(.A1(new_n1206), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n1235));
  NAND3_X1  g810(.A1(new_n1232), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  NAND3_X1  g811(.A1(new_n1146), .A2(new_n1226), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g812(.A(KEYINPUT124), .ZN(new_n1238));
  NAND2_X1  g813(.A1(G290), .A2(G1986), .ZN(new_n1239));
  NAND3_X1  g814(.A1(new_n1037), .A2(new_n1040), .A3(new_n1239), .ZN(new_n1240));
  NAND2_X1  g815(.A1(new_n1240), .A2(new_n1024), .ZN(new_n1241));
  AND3_X1   g816(.A1(new_n1237), .A2(new_n1238), .A3(new_n1241), .ZN(new_n1242));
  AOI21_X1  g817(.A(new_n1238), .B1(new_n1237), .B2(new_n1241), .ZN(new_n1243));
  OAI21_X1  g818(.A(new_n1047), .B1(new_n1242), .B2(new_n1243), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g819(.A1(new_n670), .A2(G319), .A3(new_n671), .ZN(new_n1246));
  INV_X1    g820(.A(KEYINPUT126), .ZN(new_n1247));
  OAI21_X1  g821(.A(new_n654), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g822(.A(new_n1248), .B1(new_n1247), .B2(new_n1246), .ZN(new_n1249));
  NAND3_X1  g823(.A1(new_n706), .A2(KEYINPUT127), .A3(new_n1249), .ZN(new_n1250));
  NOR2_X1   g824(.A1(new_n703), .A2(new_n705), .ZN(new_n1251));
  AOI21_X1  g825(.A(new_n704), .B1(new_n700), .B2(new_n702), .ZN(new_n1252));
  OAI21_X1  g826(.A(new_n1249), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g827(.A(KEYINPUT127), .ZN(new_n1254));
  NAND2_X1  g828(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g829(.A1(new_n1250), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g830(.A1(new_n947), .A2(new_n952), .ZN(new_n1257));
  AND3_X1   g831(.A1(new_n1256), .A2(new_n1257), .A3(new_n1010), .ZN(G308));
  NAND3_X1  g832(.A1(new_n1256), .A2(new_n1257), .A3(new_n1010), .ZN(G225));
endmodule


