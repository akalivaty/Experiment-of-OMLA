//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G128), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n190), .B(new_n192), .C1(KEYINPUT1), .C2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G125), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  XOR2_X1   g014(.A(KEYINPUT0), .B(G128), .Z(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(KEYINPUT64), .A3(new_n193), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n203));
  XNOR2_X1  g017(.A(G143), .B(G146), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT0), .B(G128), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n204), .A2(KEYINPUT0), .A3(G128), .ZN(new_n207));
  AND3_X1   g021(.A1(new_n202), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n200), .B1(new_n208), .B2(new_n199), .ZN(new_n209));
  INV_X1    g023(.A(G224), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G953), .ZN(new_n211));
  XNOR2_X1  g025(.A(new_n209), .B(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT3), .B1(new_n213), .B2(G107), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n215));
  INV_X1    g029(.A(G107), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(G104), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n213), .A2(G107), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n214), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT4), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G101), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(G116), .B(G119), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT2), .B(G113), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n223), .B(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n219), .A2(G101), .ZN(new_n227));
  AOI21_X1  g041(.A(G101), .B1(new_n213), .B2(G107), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n214), .A2(new_n228), .A3(new_n217), .ZN(new_n229));
  AND4_X1   g043(.A1(KEYINPUT79), .A2(new_n227), .A3(KEYINPUT4), .A4(new_n229), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n229), .A2(KEYINPUT4), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT79), .B1(new_n231), .B2(new_n227), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n226), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT84), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT80), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n235), .B1(new_n213), .B2(G107), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n216), .A2(KEYINPUT80), .A3(G104), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n218), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G101), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(new_n229), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT81), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(KEYINPUT81), .A3(new_n229), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n223), .A2(KEYINPUT5), .ZN(new_n245));
  INV_X1    g059(.A(G116), .ZN(new_n246));
  NOR3_X1   g060(.A1(new_n246), .A2(KEYINPUT5), .A3(G119), .ZN(new_n247));
  INV_X1    g061(.A(G113), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n224), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n245), .A2(new_n249), .B1(new_n250), .B2(new_n223), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n244), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT84), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n226), .B(new_n253), .C1(new_n230), .C2(new_n232), .ZN(new_n254));
  XNOR2_X1  g068(.A(G110), .B(G122), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n234), .A2(new_n252), .A3(new_n254), .A4(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n234), .A2(new_n252), .A3(new_n254), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n255), .B(KEYINPUT85), .ZN(new_n258));
  AOI22_X1  g072(.A1(KEYINPUT6), .A2(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n260));
  INV_X1    g074(.A(new_n258), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n250), .A2(new_n223), .ZN(new_n262));
  INV_X1    g076(.A(new_n223), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(new_n224), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(new_n221), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n227), .A2(KEYINPUT4), .A3(new_n229), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT79), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n231), .A2(KEYINPUT79), .A3(new_n227), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n266), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n271), .A2(new_n253), .B1(new_n244), .B2(new_n251), .ZN(new_n272));
  AOI211_X1 g086(.A(new_n260), .B(new_n261), .C1(new_n272), .C2(new_n234), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n212), .B1(new_n259), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT7), .B1(new_n210), .B2(G953), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n209), .B(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n255), .B(KEYINPUT8), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n239), .A2(KEYINPUT86), .A3(new_n229), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n277), .B1(new_n278), .B2(new_n251), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n279), .B1(new_n251), .B2(new_n278), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(G902), .B1(new_n281), .B2(new_n256), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n274), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(G210), .B1(G237), .B2(G902), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT87), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT87), .ZN(new_n287));
  AOI211_X1 g101(.A(new_n287), .B(new_n284), .C1(new_n274), .C2(new_n282), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n274), .A2(new_n282), .A3(new_n284), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT88), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT88), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n274), .A2(new_n292), .A3(new_n282), .A4(new_n284), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n188), .B1(new_n289), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G137), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G134), .ZN(new_n297));
  NAND2_X1  g111(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G134), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G137), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  OR2_X1    g116(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n297), .B1(new_n303), .B2(new_n298), .ZN(new_n304));
  OAI21_X1  g118(.A(G131), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n298), .ZN(new_n306));
  NOR2_X1   g120(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n307));
  OAI211_X1 g121(.A(G134), .B(new_n296), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G131), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n308), .A2(new_n309), .A3(new_n301), .A4(new_n299), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n208), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n198), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n297), .A2(KEYINPUT67), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n301), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n297), .A2(KEYINPUT67), .ZN(new_n316));
  OAI21_X1  g130(.A(G131), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n313), .A2(new_n317), .A3(new_n310), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT30), .ZN(new_n320));
  INV_X1    g134(.A(new_n318), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT66), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n312), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n208), .A2(new_n311), .A3(KEYINPUT66), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n321), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n320), .B(new_n265), .C1(new_n325), .C2(KEYINPUT30), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n327));
  INV_X1    g141(.A(G210), .ZN(new_n328));
  NOR3_X1   g142(.A1(new_n328), .A2(G237), .A3(G953), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n327), .B(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT26), .B(G101), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n330), .B(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n312), .A2(new_n225), .A3(new_n318), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n326), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT31), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(KEYINPUT28), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT28), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n312), .A2(new_n318), .A3(new_n337), .A4(new_n225), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n339), .B1(new_n225), .B2(new_n325), .ZN(new_n340));
  INV_X1    g154(.A(new_n332), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT31), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n326), .A2(new_n343), .A3(new_n332), .A4(new_n333), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n335), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT32), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n346), .A2(G472), .A3(G902), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT71), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT71), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n345), .A2(new_n350), .A3(new_n347), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n323), .A2(new_n324), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n318), .ZN(new_n354));
  AOI22_X1  g168(.A1(new_n354), .A2(new_n265), .B1(new_n336), .B2(new_n338), .ZN(new_n355));
  AOI21_X1  g169(.A(KEYINPUT29), .B1(new_n355), .B2(new_n332), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n326), .A2(new_n333), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n356), .B(KEYINPUT70), .C1(new_n357), .C2(new_n332), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT70), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT29), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n360), .B1(new_n340), .B2(new_n341), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n332), .B1(new_n326), .B2(new_n333), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n319), .A2(new_n225), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(new_n336), .B2(new_n338), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n341), .A2(new_n360), .ZN(new_n366));
  AOI21_X1  g180(.A(G902), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n358), .A2(new_n363), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G472), .ZN(new_n369));
  NOR2_X1   g183(.A1(G472), .A2(G902), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n345), .A2(new_n370), .ZN(new_n371));
  XOR2_X1   g185(.A(KEYINPUT69), .B(KEYINPUT32), .Z(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n352), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT20), .ZN(new_n375));
  XNOR2_X1  g189(.A(G113), .B(G122), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(new_n213), .ZN(new_n377));
  INV_X1    g191(.A(G237), .ZN(new_n378));
  INV_X1    g192(.A(G953), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n378), .A2(new_n379), .A3(G214), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(new_n191), .ZN(new_n381));
  NAND2_X1  g195(.A1(KEYINPUT18), .A2(G131), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n381), .B(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G140), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G125), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n199), .A2(G140), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT74), .ZN(new_n387));
  OR3_X1    g201(.A1(new_n199), .A2(KEYINPUT74), .A3(G140), .ZN(new_n388));
  AND2_X1   g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G146), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n385), .A2(new_n386), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n189), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n383), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n381), .A2(G131), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n380), .B(G143), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n309), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT17), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n395), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n395), .A2(new_n398), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT16), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT16), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n385), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G146), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n401), .A2(new_n189), .A3(new_n403), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(KEYINPUT75), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT75), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n404), .A2(new_n408), .A3(G146), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n400), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT90), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n399), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI211_X1 g226(.A(KEYINPUT90), .B(new_n400), .C1(new_n407), .C2(new_n409), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n377), .B(new_n394), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n395), .A2(new_n397), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT89), .ZN(new_n416));
  OR2_X1    g230(.A1(new_n391), .A2(KEYINPUT19), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT19), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n417), .B1(new_n389), .B2(new_n418), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n415), .A2(new_n416), .B1(new_n419), .B2(new_n189), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT77), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n405), .A2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n404), .A2(KEYINPUT77), .A3(G146), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n420), .B(new_n424), .C1(new_n416), .C2(new_n415), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n394), .ZN(new_n426));
  INV_X1    g240(.A(new_n377), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n414), .A2(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(G475), .A2(G902), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n375), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n430), .ZN(new_n432));
  AOI211_X1 g246(.A(KEYINPUT20), .B(new_n432), .C1(new_n414), .C2(new_n428), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n394), .B1(new_n412), .B2(new_n413), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n427), .ZN(new_n435));
  AOI21_X1  g249(.A(G902), .B1(new_n435), .B2(new_n414), .ZN(new_n436));
  INV_X1    g250(.A(G475), .ZN(new_n437));
  OAI22_X1  g251(.A1(new_n431), .A2(new_n433), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(G234), .A2(G237), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(G952), .A3(new_n379), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(G898), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n439), .A2(G902), .A3(G953), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n440), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n196), .A2(G143), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT13), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n196), .A2(G143), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(KEYINPUT92), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n446), .A2(KEYINPUT13), .ZN(new_n450));
  OAI221_X1 g264(.A(G134), .B1(KEYINPUT92), .B2(new_n447), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n446), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n452), .A2(new_n448), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n300), .ZN(new_n454));
  INV_X1    g268(.A(G122), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G116), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT91), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n246), .A2(G122), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n216), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n216), .B1(new_n458), .B2(new_n459), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n451), .B(new_n454), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n453), .B(new_n300), .ZN(new_n464));
  INV_X1    g278(.A(new_n458), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n459), .B(KEYINPUT14), .ZN(new_n466));
  OAI21_X1  g280(.A(G107), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n464), .A2(new_n460), .A3(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT9), .B(G234), .ZN(new_n469));
  INV_X1    g283(.A(G217), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n469), .A2(new_n470), .A3(G953), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n463), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT93), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n463), .A2(new_n468), .ZN(new_n475));
  INV_X1    g289(.A(new_n471), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n463), .A2(new_n468), .A3(KEYINPUT93), .A4(new_n471), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n474), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G902), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT15), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n481), .A2(new_n482), .A3(G478), .ZN(new_n483));
  INV_X1    g297(.A(G478), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n479), .B(new_n480), .C1(KEYINPUT15), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n438), .A2(new_n445), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n470), .B1(G234), .B2(new_n480), .ZN(new_n488));
  XNOR2_X1  g302(.A(KEYINPUT22), .B(G137), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n379), .A2(G221), .A3(G234), .ZN(new_n490));
  XOR2_X1   g304(.A(new_n489), .B(new_n490), .Z(new_n491));
  OR2_X1    g305(.A1(new_n196), .A2(G119), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n196), .A2(G119), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT24), .B(G110), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT73), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT23), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT23), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(KEYINPUT73), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n498), .A2(new_n493), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT72), .ZN(new_n502));
  NAND2_X1  g316(.A1(KEYINPUT23), .A2(G119), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n502), .B1(new_n503), .B2(G128), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n196), .A2(KEYINPUT72), .A3(KEYINPUT23), .A4(G119), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n501), .A2(new_n492), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n496), .B1(new_n506), .B2(G110), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n407), .A2(new_n409), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT76), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT76), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n407), .A2(new_n510), .A3(new_n409), .A4(new_n507), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n494), .A2(new_n495), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n506), .B2(G110), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n392), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n515), .B1(new_n422), .B2(new_n423), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n491), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n491), .ZN(new_n519));
  AOI211_X1 g333(.A(new_n516), .B(new_n519), .C1(new_n509), .C2(new_n511), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT25), .B1(new_n521), .B2(new_n480), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT25), .ZN(new_n523));
  NOR4_X1   g337(.A1(new_n518), .A2(new_n520), .A3(new_n523), .A4(G902), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n488), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(G221), .B1(new_n469), .B2(G902), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(G469), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n528), .A2(new_n480), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n379), .A2(G227), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(KEYINPUT78), .ZN(new_n531));
  XNOR2_X1  g345(.A(G110), .B(G140), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n240), .A2(new_n198), .ZN(new_n534));
  AOI22_X1  g348(.A1(new_n239), .A2(new_n229), .B1(new_n195), .B2(new_n197), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n311), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT12), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g352(.A(KEYINPUT12), .B(new_n311), .C1(new_n534), .C2(new_n535), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n221), .B(new_n208), .C1(new_n230), .C2(new_n232), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT10), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n240), .B2(new_n198), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n198), .A2(new_n542), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n242), .A2(new_n544), .A3(new_n243), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n311), .A2(KEYINPUT82), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT82), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n305), .A2(new_n310), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n541), .A2(new_n543), .A3(new_n545), .A4(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n533), .B1(new_n540), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n545), .A2(new_n543), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n221), .A2(new_n202), .A3(new_n206), .A4(new_n207), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n553), .B1(new_n269), .B2(new_n270), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT83), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT83), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n541), .A2(new_n556), .A3(new_n543), .A4(new_n545), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n557), .A3(new_n311), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n550), .A2(new_n533), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n551), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n529), .B1(new_n560), .B2(G469), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n533), .B1(new_n558), .B2(new_n550), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n540), .A2(new_n550), .A3(new_n533), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n528), .B(new_n480), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n527), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n488), .A2(G902), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n521), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n525), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n295), .A2(new_n374), .A3(new_n487), .A4(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(G101), .ZN(G3));
  NAND2_X1  g385(.A1(new_n345), .A2(new_n480), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT94), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n573), .A3(G472), .ZN(new_n574));
  INV_X1    g388(.A(G472), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(new_n345), .B2(new_n480), .ZN(new_n576));
  AOI21_X1  g390(.A(KEYINPUT94), .B1(new_n345), .B2(new_n370), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n574), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n578), .A2(new_n568), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n274), .A2(new_n282), .A3(new_n284), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n284), .B1(new_n274), .B2(new_n282), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n187), .B(new_n444), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n481), .A2(new_n484), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT33), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n479), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n477), .A2(KEYINPUT33), .A3(new_n472), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n484), .A2(G902), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n583), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n438), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n582), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n579), .A2(new_n592), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT34), .B(G104), .Z(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G6));
  INV_X1    g409(.A(KEYINPUT95), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n414), .A2(new_n428), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT20), .B1(new_n597), .B2(new_n432), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n429), .A2(new_n375), .A3(new_n430), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n435), .A2(new_n414), .ZN(new_n601));
  OAI21_X1  g415(.A(G475), .B1(new_n601), .B2(G902), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n600), .A2(new_n486), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n596), .B1(new_n582), .B2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n486), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n438), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n283), .A2(new_n285), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n188), .B1(new_n608), .B2(new_n290), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n607), .A2(new_n609), .A3(KEYINPUT95), .A4(new_n444), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n579), .B1(new_n605), .B2(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT35), .B(G107), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G9));
  INV_X1    g428(.A(new_n565), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n616));
  INV_X1    g430(.A(new_n488), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n512), .A2(new_n517), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n519), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n512), .A2(new_n517), .A3(new_n491), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(new_n480), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(new_n523), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n521), .A2(KEYINPUT25), .A3(new_n480), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n617), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n519), .A2(KEYINPUT36), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n618), .B(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n626), .A2(G902), .A3(new_n488), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n616), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n626), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n566), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n525), .A2(KEYINPUT96), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n615), .B1(new_n628), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n578), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n632), .A2(new_n633), .A3(new_n295), .A4(new_n487), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT97), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT37), .B(G110), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G12));
  AND2_X1   g451(.A1(new_n632), .A2(new_n374), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT98), .B(G900), .Z(new_n639));
  OR2_X1    g453(.A1(new_n639), .A2(new_n443), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n440), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n600), .A2(new_n602), .A3(new_n486), .A4(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n187), .B1(new_n580), .B2(new_n581), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n638), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G128), .ZN(G30));
  NAND2_X1  g460(.A1(new_n608), .A2(new_n287), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n581), .A2(KEYINPUT87), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n294), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT38), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n641), .B(KEYINPUT39), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n565), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT40), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n628), .A2(new_n631), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  AOI22_X1  g470(.A1(new_n349), .A2(new_n351), .B1(new_n372), .B2(new_n371), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n357), .A2(new_n341), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n333), .A2(new_n341), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n480), .B1(new_n364), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(G472), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n606), .B1(new_n600), .B2(new_n602), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n656), .A2(new_n662), .A3(new_n187), .A4(new_n663), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n654), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G143), .ZN(G45));
  NAND3_X1  g480(.A1(new_n438), .A2(new_n590), .A3(new_n641), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n643), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n638), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G146), .ZN(G48));
  INV_X1    g484(.A(new_n567), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n624), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n480), .B1(new_n562), .B2(new_n563), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(G469), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n564), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n527), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n374), .A2(new_n672), .A3(new_n592), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(KEYINPUT41), .B(G113), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT99), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n677), .B(new_n679), .ZN(G15));
  NAND2_X1  g494(.A1(new_n525), .A2(new_n567), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n681), .B1(new_n657), .B2(new_n369), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n682), .B(new_n676), .C1(new_n605), .C2(new_n611), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G116), .ZN(G18));
  NOR3_X1   g498(.A1(new_n643), .A2(new_n527), .A3(new_n675), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n374), .A2(new_n685), .A3(new_n655), .A4(new_n487), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G119), .ZN(G21));
  OAI211_X1 g501(.A(new_n335), .B(new_n344), .C1(new_n332), .C2(new_n365), .ZN(new_n688));
  AOI22_X1  g502(.A1(new_n572), .A2(G472), .B1(new_n370), .B2(new_n688), .ZN(new_n689));
  AND4_X1   g503(.A1(new_n444), .A2(new_n674), .A3(new_n526), .A4(new_n564), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n672), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n438), .A2(new_n486), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT100), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n692), .A2(new_n643), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(KEYINPUT100), .B1(new_n663), .B2(new_n609), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n691), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G122), .ZN(G24));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n667), .A2(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n438), .A2(KEYINPUT101), .A3(new_n590), .A4(new_n641), .ZN(new_n700));
  AND4_X1   g514(.A1(new_n655), .A2(new_n689), .A3(new_n699), .A4(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n685), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G125), .ZN(G27));
  NAND2_X1  g517(.A1(new_n371), .A2(new_n346), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n369), .A2(new_n348), .A3(new_n704), .ZN(new_n705));
  AND4_X1   g519(.A1(new_n672), .A2(new_n699), .A3(new_n705), .A4(new_n700), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n289), .A2(new_n187), .A3(new_n294), .A4(new_n565), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n707), .A2(KEYINPUT102), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(KEYINPUT102), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n706), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n374), .A2(new_n672), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n294), .A2(new_n647), .A3(new_n648), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT102), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n712), .A2(new_n713), .A3(new_n187), .A4(new_n565), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n707), .A2(KEYINPUT102), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n711), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n699), .A2(new_n700), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(KEYINPUT42), .ZN(new_n718));
  AOI22_X1  g532(.A1(new_n710), .A2(KEYINPUT42), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G131), .ZN(G33));
  XOR2_X1   g534(.A(new_n642), .B(KEYINPUT103), .Z(new_n721));
  OAI211_X1 g535(.A(new_n721), .B(new_n682), .C1(new_n708), .C2(new_n709), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(KEYINPUT104), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n716), .A2(new_n724), .A3(new_n721), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G134), .ZN(G36));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n728));
  INV_X1    g542(.A(new_n590), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n728), .B1(new_n438), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(KEYINPUT105), .ZN(new_n731));
  OR2_X1    g545(.A1(new_n438), .A2(KEYINPUT106), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n438), .A2(KEYINPUT106), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n732), .A2(KEYINPUT43), .A3(new_n590), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n656), .A2(new_n633), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n735), .A2(KEYINPUT44), .A3(new_n736), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n289), .A2(new_n187), .A3(new_n294), .ZN(new_n741));
  INV_X1    g555(.A(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n564), .ZN(new_n743));
  INV_X1    g557(.A(new_n529), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n560), .A2(KEYINPUT45), .ZN(new_n745));
  OAI21_X1  g559(.A(G469), .B1(new_n560), .B2(KEYINPUT45), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n743), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI211_X1 g563(.A(KEYINPUT46), .B(new_n744), .C1(new_n745), .C2(new_n746), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n527), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n742), .A2(new_n751), .A3(new_n651), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n739), .A2(new_n740), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G137), .ZN(G39));
  NOR2_X1   g568(.A1(new_n374), .A2(new_n672), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n741), .A2(new_n667), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n749), .A2(new_n750), .ZN(new_n757));
  AND3_X1   g571(.A1(new_n757), .A2(KEYINPUT47), .A3(new_n526), .ZN(new_n758));
  AOI21_X1  g572(.A(KEYINPUT47), .B1(new_n757), .B2(new_n526), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n755), .B(new_n756), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G140), .ZN(G42));
  NOR2_X1   g575(.A1(new_n675), .A2(KEYINPUT49), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT107), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n763), .A2(new_n733), .A3(new_n732), .ZN(new_n764));
  INV_X1    g578(.A(new_n650), .ZN(new_n765));
  INV_X1    g579(.A(new_n662), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n590), .A2(new_n187), .A3(new_n526), .ZN(new_n767));
  AOI211_X1 g581(.A(new_n767), .B(new_n681), .C1(KEYINPUT49), .C2(new_n675), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n764), .A2(new_n765), .A3(new_n766), .A4(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n701), .B1(new_n708), .B2(new_n709), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT109), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n600), .A2(new_n606), .A3(new_n602), .ZN(new_n773));
  INV_X1    g587(.A(new_n641), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n773), .A2(new_n772), .A3(new_n774), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n741), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n638), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n771), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n779), .B1(new_n723), .B2(new_n725), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n683), .A2(new_n677), .A3(new_n686), .A4(new_n696), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT108), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n782), .B1(new_n438), .B2(new_n606), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n600), .A2(new_n602), .A3(KEYINPUT108), .A4(new_n486), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n784), .A3(new_n591), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n579), .A2(new_n295), .A3(new_n444), .A4(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(new_n570), .A3(new_n634), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n781), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n780), .A2(new_n719), .A3(new_n788), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n694), .A2(new_n695), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n615), .A2(new_n624), .A3(new_n627), .A4(new_n774), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n790), .A2(new_n662), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n638), .B1(new_n644), .B2(new_n668), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(new_n793), .A3(new_n702), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT52), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n770), .B1(new_n789), .B2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n794), .B(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n781), .B(KEYINPUT112), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n710), .A2(KEYINPUT42), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n716), .A2(new_n718), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n786), .A2(new_n570), .A3(new_n634), .ZN(new_n802));
  AND4_X1   g616(.A1(KEYINPUT53), .A2(new_n800), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n798), .A2(new_n799), .A3(new_n780), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n796), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(KEYINPUT54), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT51), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n742), .A2(new_n676), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n440), .B1(new_n808), .B2(KEYINPUT114), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n742), .A2(new_n810), .A3(new_n676), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n662), .A2(new_n681), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n809), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n809), .A2(KEYINPUT116), .A3(new_n811), .A4(new_n812), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n438), .A2(new_n590), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n672), .A2(new_n689), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n440), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n735), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(KEYINPUT113), .A2(KEYINPUT50), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n675), .A2(new_n187), .A3(new_n527), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n821), .A2(new_n765), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n759), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n751), .A2(KEYINPUT47), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n825), .B(new_n826), .C1(new_n526), .C2(new_n675), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n821), .A2(new_n827), .A3(new_n742), .ZN(new_n828));
  XOR2_X1   g642(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n829));
  NAND2_X1  g643(.A1(new_n765), .A2(new_n823), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n735), .A2(new_n820), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n824), .A2(new_n828), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n818), .A2(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n655), .A2(new_n689), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n809), .A2(new_n835), .A3(new_n735), .A4(new_n811), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n836), .B(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n807), .B1(new_n834), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n833), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n807), .A2(new_n840), .A3(new_n838), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n379), .A2(G952), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(new_n821), .B2(new_n685), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n705), .A2(new_n672), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n809), .A2(new_n846), .A3(new_n735), .A4(new_n811), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n847), .A2(KEYINPUT48), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(KEYINPUT48), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n845), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n591), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n815), .A2(new_n852), .A3(new_n816), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT117), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n847), .A2(KEYINPUT48), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n844), .B1(new_n856), .B2(new_n848), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT117), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n857), .A2(new_n853), .A3(new_n858), .ZN(new_n859));
  OAI22_X1  g673(.A1(new_n839), .A2(new_n842), .B1(new_n855), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT110), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n771), .A2(new_n778), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n714), .A2(new_n715), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n724), .A2(new_n863), .A3(new_n682), .A4(new_n721), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n724), .B1(new_n716), .B2(new_n721), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n604), .A2(new_n610), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n374), .A2(new_n672), .A3(new_n676), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n696), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n677), .A2(new_n686), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n871), .A2(new_n800), .A3(new_n801), .A4(new_n802), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n861), .B1(new_n866), .B2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n780), .A2(new_n719), .A3(KEYINPUT110), .A4(new_n788), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(new_n874), .A3(new_n798), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n770), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT111), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT111), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n875), .A2(new_n878), .A3(new_n770), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n789), .A2(new_n795), .A3(new_n770), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n877), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  AOI211_X1 g696(.A(new_n806), .B(new_n860), .C1(new_n882), .C2(KEYINPUT54), .ZN(new_n883));
  NOR2_X1   g697(.A1(G952), .A2(G953), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT118), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n769), .B1(new_n883), .B2(new_n885), .ZN(G75));
  AND2_X1   g700(.A1(new_n796), .A2(new_n804), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n887), .A2(new_n328), .A3(new_n480), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(KEYINPUT56), .ZN(new_n889));
  INV_X1    g703(.A(new_n259), .ZN(new_n890));
  INV_X1    g704(.A(new_n273), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(new_n212), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT55), .Z(new_n894));
  NOR2_X1   g708(.A1(new_n889), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n379), .A2(G952), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  XOR2_X1   g711(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n898));
  NAND2_X1  g712(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n897), .B1(new_n888), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n895), .A2(new_n900), .ZN(G51));
  XNOR2_X1  g715(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(new_n529), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT54), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n796), .B2(new_n804), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n903), .B1(new_n806), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n906), .B1(new_n562), .B2(new_n563), .ZN(new_n907));
  OR4_X1    g721(.A1(new_n480), .A2(new_n887), .A3(new_n745), .A4(new_n746), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n896), .B1(new_n907), .B2(new_n908), .ZN(G54));
  NAND4_X1  g723(.A1(new_n805), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n910), .A2(new_n597), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n597), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n911), .A2(new_n912), .A3(new_n896), .ZN(G60));
  XNOR2_X1  g727(.A(new_n587), .B(KEYINPUT121), .ZN(new_n914));
  NAND2_X1  g728(.A1(G478), .A2(G902), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT59), .Z(new_n916));
  NOR2_X1   g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n917), .B1(new_n806), .B2(new_n905), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n897), .ZN(new_n919));
  INV_X1    g733(.A(new_n916), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n880), .B1(new_n876), .B2(KEYINPUT111), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n904), .B1(new_n921), .B2(new_n879), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n920), .B1(new_n922), .B2(new_n806), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n919), .B1(new_n923), .B2(new_n914), .ZN(G63));
  NAND2_X1  g738(.A1(G217), .A2(G902), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT60), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n796), .B2(new_n804), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n629), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n928), .B(new_n897), .C1(new_n521), .C2(new_n927), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT61), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n929), .B(new_n931), .ZN(G66));
  OAI21_X1  g746(.A(G953), .B1(new_n441), .B2(new_n210), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT123), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(new_n788), .B2(G953), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n890), .B(new_n891), .C1(G898), .C2(new_n379), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n935), .B(new_n936), .ZN(G69));
  AND2_X1   g751(.A1(new_n793), .A2(new_n702), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n790), .A2(new_n651), .A3(new_n846), .A4(new_n751), .ZN(new_n939));
  AND4_X1   g753(.A1(new_n719), .A2(new_n938), .A3(new_n760), .A4(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n940), .A2(KEYINPUT124), .A3(new_n726), .A4(new_n753), .ZN(new_n941));
  AND4_X1   g755(.A1(new_n702), .A2(new_n760), .A3(new_n939), .A4(new_n793), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n942), .A2(new_n753), .A3(new_n726), .A4(new_n719), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT124), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n379), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n379), .A2(G900), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n947), .A2(KEYINPUT125), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n951));
  AOI21_X1  g765(.A(G953), .B1(new_n941), .B2(new_n945), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n951), .B1(new_n952), .B2(new_n948), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n320), .B1(new_n325), .B2(KEYINPUT30), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(new_n419), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n938), .A2(new_n665), .A3(new_n959), .ZN(new_n960));
  OAI211_X1 g774(.A(new_n793), .B(new_n702), .C1(new_n654), .C2(new_n664), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(KEYINPUT62), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n682), .A2(new_n742), .A3(new_n652), .A4(new_n785), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n760), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n960), .A2(new_n962), .A3(new_n753), .A4(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n965), .A2(new_n379), .A3(new_n956), .ZN(new_n966));
  INV_X1    g780(.A(G227), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n948), .B1(new_n967), .B2(G953), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT126), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n958), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n969), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n956), .B1(new_n950), .B2(new_n953), .ZN(new_n972));
  INV_X1    g786(.A(new_n966), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n970), .A2(new_n974), .ZN(G72));
  NAND2_X1  g789(.A1(G472), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT63), .Z(new_n977));
  INV_X1    g791(.A(new_n788), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n977), .B1(new_n946), .B2(new_n978), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n326), .A2(new_n341), .A3(new_n333), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n977), .B1(new_n965), .B2(new_n978), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n658), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n981), .A2(new_n897), .A3(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n977), .ZN(new_n985));
  OR3_X1    g799(.A1(new_n658), .A2(new_n985), .A3(new_n980), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n986), .B1(new_n921), .B2(new_n879), .ZN(new_n987));
  OAI21_X1  g801(.A(KEYINPUT127), .B1(new_n984), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT127), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n983), .A2(new_n897), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n990), .B1(new_n980), .B2(new_n979), .ZN(new_n991));
  INV_X1    g805(.A(new_n882), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n989), .B(new_n991), .C1(new_n992), .C2(new_n986), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n988), .A2(new_n993), .ZN(G57));
endmodule


