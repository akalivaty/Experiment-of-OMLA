

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765;

  OR2_X1 U369 ( .A1(n670), .A2(n671), .ZN(n667) );
  AND2_X1 U370 ( .A1(G221), .A2(n513), .ZN(n448) );
  XNOR2_X1 U371 ( .A(n472), .B(n447), .ZN(n482) );
  XNOR2_X1 U372 ( .A(G119), .B(G110), .ZN(n493) );
  XNOR2_X1 U373 ( .A(G113), .B(G104), .ZN(n520) );
  XNOR2_X1 U374 ( .A(G122), .B(G116), .ZN(n507) );
  XNOR2_X1 U375 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n522) );
  BUF_X1 U376 ( .A(n450), .Z(n405) );
  INV_X1 U377 ( .A(KEYINPUT80), .ZN(n453) );
  XNOR2_X2 U378 ( .A(n497), .B(n496), .ZN(n735) );
  NAND2_X2 U379 ( .A1(n364), .A2(n363), .ZN(n362) );
  AND2_X2 U380 ( .A1(n598), .A2(n597), .ZN(n449) );
  XNOR2_X2 U381 ( .A(n385), .B(n384), .ZN(n513) );
  XNOR2_X2 U382 ( .A(n502), .B(n501), .ZN(n670) );
  INV_X2 U383 ( .A(n699), .ZN(n373) );
  BUF_X2 U384 ( .A(n405), .Z(n347) );
  NOR2_X2 U385 ( .A1(n347), .A2(G952), .ZN(n737) );
  XNOR2_X2 U386 ( .A(n585), .B(n464), .ZN(n573) );
  XNOR2_X2 U387 ( .A(n436), .B(n435), .ZN(n585) );
  XNOR2_X1 U388 ( .A(G146), .B(G137), .ZN(n473) );
  XNOR2_X1 U389 ( .A(G146), .B(G101), .ZN(n484) );
  AND2_X1 U390 ( .A1(n552), .A2(n360), .ZN(n640) );
  XNOR2_X2 U391 ( .A(n478), .B(n459), .ZN(n739) );
  XNOR2_X2 U392 ( .A(n430), .B(n452), .ZN(n440) );
  NOR2_X2 U393 ( .A1(n573), .A2(n469), .ZN(n471) );
  NOR2_X2 U394 ( .A1(G902), .A2(n721), .ZN(n529) );
  NAND2_X1 U395 ( .A1(n358), .A2(n357), .ZN(n356) );
  OR2_X1 U396 ( .A1(n702), .A2(n703), .ZN(n358) );
  XNOR2_X1 U397 ( .A(n482), .B(n490), .ZN(n751) );
  XNOR2_X1 U398 ( .A(n349), .B(n397), .ZN(n752) );
  XNOR2_X1 U399 ( .A(n354), .B(KEYINPUT94), .ZN(n451) );
  INV_X1 U400 ( .A(KEYINPUT79), .ZN(n352) );
  XNOR2_X1 U401 ( .A(G128), .B(KEYINPUT97), .ZN(n491) );
  XNOR2_X1 U402 ( .A(n356), .B(n355), .ZN(G75) );
  NOR2_X1 U403 ( .A1(n704), .A2(n705), .ZN(n357) );
  NOR2_X1 U404 ( .A1(n426), .A2(n602), .ZN(n382) );
  XNOR2_X1 U405 ( .A(n415), .B(n414), .ZN(n657) );
  OR2_X1 U406 ( .A1(G953), .A2(n666), .ZN(n705) );
  INV_X1 U407 ( .A(n539), .ZN(n348) );
  OR2_X1 U408 ( .A1(n389), .A2(n388), .ZN(n607) );
  XNOR2_X1 U409 ( .A(n538), .B(n537), .ZN(n692) );
  NAND2_X1 U410 ( .A1(n536), .A2(n548), .ZN(n538) );
  XNOR2_X1 U411 ( .A(n505), .B(n408), .ZN(n668) );
  XNOR2_X1 U412 ( .A(n516), .B(G478), .ZN(n533) );
  XOR2_X1 U413 ( .A(n716), .B(n715), .Z(n718) );
  XNOR2_X1 U414 ( .A(n488), .B(n489), .ZN(n505) );
  NOR2_X1 U415 ( .A1(G902), .A2(n712), .ZN(n488) );
  INV_X1 U416 ( .A(n451), .ZN(n452) );
  XNOR2_X1 U417 ( .A(n484), .B(n352), .ZN(n351) );
  XNOR2_X1 U418 ( .A(n491), .B(n403), .ZN(n402) );
  XOR2_X1 U419 ( .A(KEYINPUT9), .B(G134), .Z(n511) );
  XOR2_X2 U420 ( .A(G119), .B(KEYINPUT96), .Z(n458) );
  INV_X2 U421 ( .A(KEYINPUT18), .ZN(n354) );
  INV_X1 U422 ( .A(KEYINPUT24), .ZN(n403) );
  XOR2_X2 U423 ( .A(KEYINPUT77), .B(KEYINPUT5), .Z(n474) );
  XOR2_X2 U424 ( .A(KEYINPUT7), .B(G107), .Z(n508) );
  XOR2_X2 U425 ( .A(KEYINPUT104), .B(KEYINPUT103), .Z(n523) );
  NOR2_X1 U426 ( .A1(G953), .A2(G237), .ZN(n517) );
  XNOR2_X1 U427 ( .A(n349), .B(KEYINPUT17), .ZN(n439) );
  XNOR2_X2 U428 ( .A(n353), .B(G146), .ZN(n349) );
  NAND2_X1 U429 ( .A1(n450), .A2(G224), .ZN(n430) );
  XNOR2_X2 U430 ( .A(n383), .B(G953), .ZN(n450) );
  XNOR2_X2 U431 ( .A(G110), .B(G104), .ZN(n456) );
  XNOR2_X2 U432 ( .A(n456), .B(G107), .ZN(n483) );
  AND2_X1 U433 ( .A1(n350), .A2(n574), .ZN(n404) );
  NAND2_X1 U434 ( .A1(n657), .A2(n434), .ZN(n350) );
  INV_X2 U435 ( .A(G125), .ZN(n353) );
  INV_X2 U436 ( .A(KEYINPUT64), .ZN(n383) );
  XNOR2_X1 U437 ( .A(n483), .B(n351), .ZN(n486) );
  AND2_X2 U438 ( .A1(n367), .A2(n366), .ZN(n365) );
  NAND2_X2 U439 ( .A1(n365), .A2(n362), .ZN(n631) );
  INV_X1 U440 ( .A(KEYINPUT53), .ZN(n355) );
  NAND2_X1 U441 ( .A1(n603), .A2(n359), .ZN(n426) );
  XOR2_X1 U442 ( .A(G131), .B(G134), .Z(n447) );
  INV_X1 U443 ( .A(KEYINPUT19), .ZN(n464) );
  INV_X1 U444 ( .A(KEYINPUT83), .ZN(n416) );
  AND2_X1 U445 ( .A1(n382), .A2(n424), .ZN(n378) );
  NOR2_X2 U446 ( .A1(n668), .A2(n667), .ZN(n536) );
  AND2_X1 U447 ( .A1(n604), .A2(n444), .ZN(n443) );
  INV_X1 U448 ( .A(n671), .ZN(n444) );
  XNOR2_X1 U449 ( .A(n480), .B(n479), .ZN(n589) );
  INV_X1 U450 ( .A(G472), .ZN(n479) );
  XNOR2_X1 U451 ( .A(G137), .B(G140), .ZN(n481) );
  XNOR2_X1 U452 ( .A(n492), .B(n402), .ZN(n494) );
  INV_X1 U453 ( .A(KEYINPUT10), .ZN(n397) );
  AND2_X1 U454 ( .A1(n369), .A2(n368), .ZN(n367) );
  OR2_X1 U455 ( .A1(n627), .A2(n371), .ZN(n368) );
  NOR2_X1 U456 ( .A1(n372), .A2(n371), .ZN(n363) );
  INV_X1 U457 ( .A(KEYINPUT8), .ZN(n384) );
  XNOR2_X1 U458 ( .A(n572), .B(KEYINPUT110), .ZN(n388) );
  INV_X1 U459 ( .A(KEYINPUT28), .ZN(n390) );
  INV_X1 U460 ( .A(KEYINPUT92), .ZN(n435) );
  INV_X1 U461 ( .A(n684), .ZN(n437) );
  XNOR2_X1 U462 ( .A(n653), .B(KEYINPUT84), .ZN(n427) );
  INV_X1 U463 ( .A(KEYINPUT90), .ZN(n556) );
  AND2_X1 U464 ( .A1(n627), .A2(n371), .ZN(n370) );
  INV_X1 U465 ( .A(KEYINPUT65), .ZN(n371) );
  XOR2_X1 U466 ( .A(G140), .B(G131), .Z(n519) );
  NAND2_X1 U467 ( .A1(G237), .A2(G234), .ZN(n465) );
  INV_X1 U468 ( .A(KEYINPUT106), .ZN(n417) );
  NOR2_X1 U469 ( .A1(G902), .A2(G237), .ZN(n460) );
  XNOR2_X1 U470 ( .A(KEYINPUT31), .B(KEYINPUT101), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n590), .B(KEYINPUT30), .ZN(n591) );
  NAND2_X1 U472 ( .A1(n589), .A2(n684), .ZN(n590) );
  NOR2_X1 U473 ( .A1(n506), .A2(KEYINPUT100), .ZN(n413) );
  XNOR2_X1 U474 ( .A(n482), .B(n429), .ZN(n632) );
  NOR2_X2 U475 ( .A1(n376), .A2(n374), .ZN(n753) );
  NAND2_X1 U476 ( .A1(n375), .A2(n624), .ZN(n374) );
  XNOR2_X1 U477 ( .A(n534), .B(KEYINPUT66), .ZN(n441) );
  NAND2_X1 U478 ( .A1(n387), .A2(n386), .ZN(n578) );
  INV_X1 U479 ( .A(n607), .ZN(n387) );
  XNOR2_X1 U480 ( .A(n723), .B(n722), .ZN(n724) );
  NAND2_X1 U481 ( .A1(n449), .A2(n428), .ZN(n653) );
  AND2_X1 U482 ( .A1(n599), .A2(n605), .ZN(n428) );
  INV_X1 U483 ( .A(n643), .ZN(n660) );
  AND2_X1 U484 ( .A1(n588), .A2(n663), .ZN(n359) );
  XNOR2_X1 U485 ( .A(n688), .B(n416), .ZN(n577) );
  NOR2_X1 U486 ( .A1(n670), .A2(n548), .ZN(n360) );
  AND2_X1 U487 ( .A1(n411), .A2(n570), .ZN(n361) );
  XNOR2_X1 U488 ( .A(G902), .B(KEYINPUT15), .ZN(n625) );
  INV_X1 U489 ( .A(n746), .ZN(n364) );
  NAND2_X1 U490 ( .A1(n746), .A2(n370), .ZN(n366) );
  NAND2_X1 U491 ( .A1(n372), .A2(n370), .ZN(n369) );
  NAND2_X1 U492 ( .A1(n373), .A2(n626), .ZN(n372) );
  XNOR2_X2 U493 ( .A(n564), .B(n563), .ZN(n746) );
  INV_X1 U494 ( .A(n657), .ZN(n394) );
  OR2_X1 U495 ( .A1(n382), .A2(n424), .ZN(n375) );
  NAND2_X1 U496 ( .A1(n379), .A2(n377), .ZN(n376) );
  NAND2_X1 U497 ( .A1(n378), .A2(n381), .ZN(n377) );
  NAND2_X1 U498 ( .A1(n380), .A2(n614), .ZN(n379) );
  INV_X1 U499 ( .A(n381), .ZN(n380) );
  XNOR2_X2 U500 ( .A(n425), .B(KEYINPUT46), .ZN(n381) );
  NAND2_X1 U501 ( .A1(n405), .A2(G234), .ZN(n385) );
  INV_X1 U502 ( .A(n578), .ZN(n654) );
  INV_X1 U503 ( .A(n573), .ZN(n386) );
  XNOR2_X1 U504 ( .A(n571), .B(n390), .ZN(n389) );
  BUF_X1 U505 ( .A(n746), .Z(n391) );
  NAND2_X1 U506 ( .A1(n348), .A2(n443), .ZN(n442) );
  XNOR2_X1 U507 ( .A(n442), .B(n441), .ZN(n547) );
  BUF_X1 U508 ( .A(n585), .Z(n392) );
  BUF_X1 U509 ( .A(n621), .Z(n393) );
  NOR2_X2 U510 ( .A1(n533), .A2(n541), .ZN(n531) );
  XNOR2_X2 U511 ( .A(n530), .B(n529), .ZN(n541) );
  XNOR2_X1 U512 ( .A(n478), .B(n477), .ZN(n429) );
  NOR2_X2 U513 ( .A1(n410), .A2(n409), .ZN(n644) );
  INV_X1 U514 ( .A(n394), .ZN(n395) );
  BUF_X1 U515 ( .A(n739), .Z(n396) );
  BUF_X1 U516 ( .A(n706), .Z(n398) );
  XNOR2_X1 U517 ( .A(n400), .B(n739), .ZN(n706) );
  XNOR2_X1 U518 ( .A(n438), .B(n472), .ZN(n400) );
  XNOR2_X1 U519 ( .A(n440), .B(n439), .ZN(n438) );
  NOR2_X1 U520 ( .A1(n726), .A2(n737), .ZN(n728) );
  NOR2_X1 U521 ( .A1(n637), .A2(n737), .ZN(n639) );
  NOR2_X1 U522 ( .A1(n736), .A2(n737), .ZN(n738) );
  INV_X2 U523 ( .A(KEYINPUT3), .ZN(n401) );
  BUF_X1 U524 ( .A(n644), .Z(n399) );
  XNOR2_X2 U525 ( .A(n419), .B(n458), .ZN(n478) );
  NAND2_X1 U526 ( .A1(n733), .A2(G217), .ZN(n734) );
  NOR2_X4 U527 ( .A1(n702), .A2(n631), .ZN(n733) );
  XNOR2_X2 U528 ( .A(n401), .B(G101), .ZN(n421) );
  NAND2_X1 U529 ( .A1(n418), .A2(n404), .ZN(n431) );
  XNOR2_X1 U530 ( .A(n630), .B(KEYINPUT78), .ZN(n702) );
  NOR2_X1 U531 ( .A1(n615), .A2(n611), .ZN(n612) );
  XNOR2_X1 U532 ( .A(n448), .B(n495), .ZN(n496) );
  NAND2_X1 U533 ( .A1(n762), .A2(KEYINPUT44), .ZN(n544) );
  XNOR2_X2 U534 ( .A(n406), .B(KEYINPUT35), .ZN(n762) );
  NAND2_X1 U535 ( .A1(n407), .A2(n599), .ZN(n406) );
  XNOR2_X1 U536 ( .A(n540), .B(KEYINPUT34), .ZN(n407) );
  INV_X1 U537 ( .A(KEYINPUT1), .ZN(n408) );
  XNOR2_X2 U538 ( .A(n510), .B(KEYINPUT4), .ZN(n472) );
  XNOR2_X2 U539 ( .A(n454), .B(n453), .ZN(n510) );
  AND2_X1 U540 ( .A1(n539), .A2(KEYINPUT100), .ZN(n409) );
  NAND2_X1 U541 ( .A1(n412), .A2(n361), .ZN(n410) );
  NAND2_X1 U542 ( .A1(n506), .A2(KEYINPUT100), .ZN(n411) );
  NAND2_X1 U543 ( .A1(n348), .A2(n413), .ZN(n412) );
  XNOR2_X2 U544 ( .A(n471), .B(n470), .ZN(n539) );
  NOR2_X2 U545 ( .A1(n539), .A2(n677), .ZN(n415) );
  NAND2_X1 U546 ( .A1(n536), .A2(n674), .ZN(n677) );
  XNOR2_X2 U547 ( .A(n532), .B(n417), .ZN(n688) );
  NAND2_X1 U548 ( .A1(n644), .A2(n434), .ZN(n418) );
  XNOR2_X2 U549 ( .A(n421), .B(n420), .ZN(n419) );
  XNOR2_X2 U550 ( .A(G113), .B(G116), .ZN(n420) );
  NAND2_X1 U551 ( .A1(n593), .A2(n422), .ZN(n598) );
  NAND2_X1 U552 ( .A1(n423), .A2(n592), .ZN(n422) );
  INV_X1 U553 ( .A(n591), .ZN(n423) );
  INV_X1 U554 ( .A(n614), .ZN(n424) );
  NOR2_X2 U555 ( .A1(n764), .A2(n765), .ZN(n425) );
  NAND2_X1 U556 ( .A1(n600), .A2(n427), .ZN(n601) );
  NOR2_X1 U557 ( .A1(n432), .A2(n431), .ZN(n535) );
  AND2_X2 U558 ( .A1(n394), .A2(n433), .ZN(n432) );
  NOR2_X1 U559 ( .A1(n644), .A2(n434), .ZN(n433) );
  INV_X1 U560 ( .A(KEYINPUT102), .ZN(n434) );
  NOR2_X2 U561 ( .A1(n621), .A2(n437), .ZN(n436) );
  XNOR2_X2 U562 ( .A(n462), .B(n461), .ZN(n621) );
  XNOR2_X1 U563 ( .A(n398), .B(n446), .ZN(n707) );
  NAND2_X1 U564 ( .A1(n706), .A2(n625), .ZN(n462) );
  NOR2_X1 U565 ( .A1(n746), .A2(n629), .ZN(n630) );
  XOR2_X1 U566 ( .A(KEYINPUT98), .B(KEYINPUT25), .Z(n445) );
  XNOR2_X1 U567 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n446) );
  NAND2_X1 U568 ( .A1(n643), .A2(n611), .ZN(n532) );
  XNOR2_X1 U569 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U570 ( .A(n486), .B(n485), .ZN(n487) );
  INV_X1 U571 ( .A(n594), .ZN(n595) );
  XNOR2_X1 U572 ( .A(n455), .B(G122), .ZN(n457) );
  XNOR2_X1 U573 ( .A(n751), .B(n487), .ZN(n712) );
  XNOR2_X1 U574 ( .A(KEYINPUT93), .B(KEYINPUT33), .ZN(n537) );
  AND2_X1 U575 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U576 ( .A(n457), .B(n483), .ZN(n459) );
  INV_X1 U577 ( .A(n533), .ZN(n542) );
  XNOR2_X1 U578 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(n729) );
  XNOR2_X1 U580 ( .A(n610), .B(n609), .ZN(n615) );
  XNOR2_X1 U581 ( .A(n500), .B(n445), .ZN(n501) );
  XNOR2_X1 U582 ( .A(n708), .B(n707), .ZN(n709) );
  XNOR2_X2 U583 ( .A(G128), .B(G143), .ZN(n454) );
  XOR2_X1 U584 ( .A(KEYINPUT74), .B(KEYINPUT16), .Z(n455) );
  XOR2_X1 U585 ( .A(KEYINPUT76), .B(n460), .Z(n463) );
  NAND2_X1 U586 ( .A1(G210), .A2(n463), .ZN(n461) );
  NAND2_X1 U587 ( .A1(G214), .A2(n463), .ZN(n684) );
  XOR2_X1 U588 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n466) );
  XNOR2_X1 U589 ( .A(n466), .B(n465), .ZN(n467) );
  NAND2_X1 U590 ( .A1(G952), .A2(n467), .ZN(n698) );
  NOR2_X1 U591 ( .A1(G953), .A2(n698), .ZN(n568) );
  INV_X1 U592 ( .A(G898), .ZN(n745) );
  NAND2_X1 U593 ( .A1(G953), .A2(n745), .ZN(n740) );
  NAND2_X1 U594 ( .A1(G902), .A2(n467), .ZN(n565) );
  NOR2_X1 U595 ( .A1(n740), .A2(n565), .ZN(n468) );
  NOR2_X1 U596 ( .A1(n568), .A2(n468), .ZN(n469) );
  INV_X1 U597 ( .A(KEYINPUT0), .ZN(n470) );
  XNOR2_X1 U598 ( .A(n474), .B(n473), .ZN(n476) );
  NAND2_X1 U599 ( .A1(G210), .A2(n517), .ZN(n475) );
  NOR2_X1 U600 ( .A1(G902), .A2(n632), .ZN(n480) );
  INV_X1 U601 ( .A(n589), .ZN(n570) );
  INV_X1 U602 ( .A(n570), .ZN(n674) );
  INV_X1 U603 ( .A(G469), .ZN(n489) );
  XNOR2_X1 U604 ( .A(n481), .B(KEYINPUT70), .ZN(n490) );
  AND2_X1 U605 ( .A1(G227), .A2(n347), .ZN(n485) );
  XOR2_X1 U606 ( .A(n752), .B(n490), .Z(n497) );
  XOR2_X1 U607 ( .A(KEYINPUT23), .B(KEYINPUT85), .Z(n492) );
  XNOR2_X1 U608 ( .A(n494), .B(n493), .ZN(n495) );
  NOR2_X1 U609 ( .A1(n735), .A2(G902), .ZN(n502) );
  XOR2_X1 U610 ( .A(KEYINPUT99), .B(KEYINPUT20), .Z(n499) );
  NAND2_X1 U611 ( .A1(G234), .A2(n625), .ZN(n498) );
  XNOR2_X1 U612 ( .A(n499), .B(n498), .ZN(n503) );
  NAND2_X1 U613 ( .A1(n503), .A2(G217), .ZN(n500) );
  NAND2_X1 U614 ( .A1(n503), .A2(G221), .ZN(n504) );
  XNOR2_X1 U615 ( .A(KEYINPUT21), .B(n504), .ZN(n671) );
  INV_X1 U616 ( .A(n505), .ZN(n572) );
  NOR2_X2 U617 ( .A1(n667), .A2(n572), .ZN(n596) );
  INV_X1 U618 ( .A(n596), .ZN(n506) );
  XNOR2_X1 U619 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U620 ( .A(n510), .B(n509), .Z(n512) );
  XNOR2_X1 U621 ( .A(n512), .B(n511), .ZN(n515) );
  NAND2_X1 U622 ( .A1(G217), .A2(n513), .ZN(n514) );
  NOR2_X1 U623 ( .A1(n729), .A2(G902), .ZN(n516) );
  XNOR2_X1 U624 ( .A(KEYINPUT13), .B(G475), .ZN(n530) );
  NAND2_X1 U625 ( .A1(n517), .A2(G214), .ZN(n518) );
  XNOR2_X1 U626 ( .A(n519), .B(n518), .ZN(n527) );
  XOR2_X1 U627 ( .A(G143), .B(G122), .Z(n521) );
  XNOR2_X1 U628 ( .A(n521), .B(n520), .ZN(n525) );
  XNOR2_X1 U629 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U630 ( .A(n525), .B(n524), .Z(n526) );
  XNOR2_X1 U631 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U632 ( .A(n752), .B(n528), .ZN(n721) );
  XNOR2_X2 U633 ( .A(n531), .B(KEYINPUT105), .ZN(n643) );
  NAND2_X1 U634 ( .A1(n541), .A2(n533), .ZN(n611) );
  INV_X1 U635 ( .A(n668), .ZN(n618) );
  NOR2_X1 U636 ( .A1(n541), .A2(n542), .ZN(n604) );
  XOR2_X1 U637 ( .A(KEYINPUT22), .B(KEYINPUT73), .Z(n534) );
  NOR2_X1 U638 ( .A1(n618), .A2(n547), .ZN(n552) );
  XOR2_X1 U639 ( .A(n570), .B(KEYINPUT6), .Z(n582) );
  INV_X1 U640 ( .A(n582), .ZN(n548) );
  NOR2_X1 U641 ( .A1(n535), .A2(n640), .ZN(n545) );
  NOR2_X1 U642 ( .A1(n539), .A2(n692), .ZN(n540) );
  NAND2_X1 U643 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U644 ( .A(n543), .B(KEYINPUT107), .ZN(n599) );
  NAND2_X1 U645 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U646 ( .A(n546), .B(KEYINPUT91), .ZN(n555) );
  NOR2_X1 U647 ( .A1(n548), .A2(n547), .ZN(n550) );
  AND2_X1 U648 ( .A1(n670), .A2(n618), .ZN(n549) );
  NAND2_X1 U649 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U650 ( .A(KEYINPUT32), .B(n551), .ZN(n763) );
  AND2_X1 U651 ( .A1(n552), .A2(n570), .ZN(n553) );
  NAND2_X1 U652 ( .A1(n553), .A2(n670), .ZN(n648) );
  NAND2_X1 U653 ( .A1(n763), .A2(n648), .ZN(n558) );
  NAND2_X1 U654 ( .A1(KEYINPUT44), .A2(n558), .ZN(n554) );
  NAND2_X1 U655 ( .A1(n555), .A2(n554), .ZN(n557) );
  XNOR2_X1 U656 ( .A(n557), .B(n556), .ZN(n562) );
  INV_X1 U657 ( .A(n558), .ZN(n560) );
  NOR2_X1 U658 ( .A1(n762), .A2(KEYINPUT44), .ZN(n559) );
  NAND2_X1 U659 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U660 ( .A1(n562), .A2(n561), .ZN(n564) );
  XOR2_X1 U661 ( .A(KEYINPUT86), .B(KEYINPUT45), .Z(n563) );
  OR2_X1 U662 ( .A1(n347), .A2(n565), .ZN(n566) );
  NOR2_X1 U663 ( .A1(G900), .A2(n566), .ZN(n567) );
  NOR2_X1 U664 ( .A1(n568), .A2(n567), .ZN(n594) );
  NOR2_X1 U665 ( .A1(n671), .A2(n594), .ZN(n569) );
  NAND2_X1 U666 ( .A1(n569), .A2(n670), .ZN(n581) );
  NOR2_X1 U667 ( .A1(n570), .A2(n581), .ZN(n571) );
  INV_X1 U668 ( .A(n577), .ZN(n574) );
  NAND2_X1 U669 ( .A1(n574), .A2(KEYINPUT69), .ZN(n575) );
  NAND2_X1 U670 ( .A1(n654), .A2(n575), .ZN(n576) );
  NAND2_X1 U671 ( .A1(n576), .A2(KEYINPUT47), .ZN(n603) );
  NOR2_X1 U672 ( .A1(KEYINPUT47), .A2(n577), .ZN(n580) );
  NOR2_X1 U673 ( .A1(KEYINPUT69), .A2(n578), .ZN(n579) );
  NAND2_X1 U674 ( .A1(n580), .A2(n579), .ZN(n588) );
  NOR2_X1 U675 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U676 ( .A(KEYINPUT108), .B(n583), .ZN(n584) );
  INV_X1 U677 ( .A(n611), .ZN(n658) );
  NAND2_X1 U678 ( .A1(n584), .A2(n658), .ZN(n617) );
  NOR2_X1 U679 ( .A1(n617), .A2(n392), .ZN(n586) );
  XNOR2_X1 U680 ( .A(n586), .B(KEYINPUT36), .ZN(n587) );
  NAND2_X1 U681 ( .A1(n587), .A2(n618), .ZN(n663) );
  INV_X1 U682 ( .A(n621), .ZN(n605) );
  NAND2_X1 U683 ( .A1(n591), .A2(KEYINPUT109), .ZN(n593) );
  INV_X1 U684 ( .A(KEYINPUT109), .ZN(n592) );
  NAND2_X1 U685 ( .A1(KEYINPUT47), .A2(n688), .ZN(n600) );
  XOR2_X1 U686 ( .A(KEYINPUT81), .B(n601), .Z(n602) );
  INV_X1 U687 ( .A(n604), .ZN(n687) );
  XOR2_X1 U688 ( .A(KEYINPUT38), .B(n605), .Z(n685) );
  NAND2_X1 U689 ( .A1(n685), .A2(n684), .ZN(n689) );
  NOR2_X1 U690 ( .A1(n687), .A2(n689), .ZN(n606) );
  XNOR2_X1 U691 ( .A(KEYINPUT41), .B(n606), .ZN(n682) );
  NOR2_X1 U692 ( .A1(n607), .A2(n682), .ZN(n608) );
  XNOR2_X1 U693 ( .A(KEYINPUT42), .B(n608), .ZN(n765) );
  NAND2_X1 U694 ( .A1(n449), .A2(n685), .ZN(n610) );
  XOR2_X1 U695 ( .A(KEYINPUT72), .B(KEYINPUT39), .Z(n609) );
  XNOR2_X1 U696 ( .A(n612), .B(KEYINPUT40), .ZN(n764) );
  XNOR2_X1 U697 ( .A(KEYINPUT89), .B(KEYINPUT48), .ZN(n613) );
  XNOR2_X1 U698 ( .A(n613), .B(KEYINPUT71), .ZN(n614) );
  NOR2_X1 U699 ( .A1(n643), .A2(n615), .ZN(n616) );
  XOR2_X1 U700 ( .A(KEYINPUT111), .B(n616), .Z(n761) );
  NOR2_X1 U701 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U702 ( .A1(n619), .A2(n684), .ZN(n620) );
  XNOR2_X1 U703 ( .A(n620), .B(KEYINPUT43), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n622), .A2(n393), .ZN(n665) );
  INV_X1 U705 ( .A(n665), .ZN(n623) );
  NOR2_X1 U706 ( .A1(n761), .A2(n623), .ZN(n624) );
  INV_X1 U707 ( .A(n753), .ZN(n699) );
  INV_X1 U708 ( .A(n625), .ZN(n626) );
  NAND2_X1 U709 ( .A1(n626), .A2(KEYINPUT2), .ZN(n627) );
  NAND2_X1 U710 ( .A1(n753), .A2(KEYINPUT2), .ZN(n628) );
  XOR2_X1 U711 ( .A(KEYINPUT87), .B(n628), .Z(n629) );
  NAND2_X1 U712 ( .A1(n733), .A2(G472), .ZN(n636) );
  INV_X1 U713 ( .A(n632), .ZN(n634) );
  XOR2_X1 U714 ( .A(KEYINPUT62), .B(KEYINPUT112), .Z(n633) );
  XNOR2_X1 U715 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U716 ( .A(KEYINPUT95), .B(KEYINPUT63), .ZN(n638) );
  XNOR2_X1 U717 ( .A(n639), .B(n638), .ZN(G57) );
  XNOR2_X1 U718 ( .A(G101), .B(n640), .ZN(n641) );
  XNOR2_X1 U719 ( .A(n641), .B(KEYINPUT113), .ZN(G3) );
  NAND2_X1 U720 ( .A1(n658), .A2(n399), .ZN(n642) );
  XNOR2_X1 U721 ( .A(n642), .B(G104), .ZN(G6) );
  XOR2_X1 U722 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n646) );
  NAND2_X1 U723 ( .A1(n660), .A2(n399), .ZN(n645) );
  XNOR2_X1 U724 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U725 ( .A(G107), .B(n647), .ZN(G9) );
  XNOR2_X1 U726 ( .A(G110), .B(KEYINPUT114), .ZN(n649) );
  XNOR2_X1 U727 ( .A(n649), .B(n648), .ZN(G12) );
  XOR2_X1 U728 ( .A(KEYINPUT29), .B(KEYINPUT115), .Z(n651) );
  NAND2_X1 U729 ( .A1(n654), .A2(n660), .ZN(n650) );
  XNOR2_X1 U730 ( .A(n651), .B(n650), .ZN(n652) );
  XOR2_X1 U731 ( .A(G128), .B(n652), .Z(G30) );
  XNOR2_X1 U732 ( .A(G143), .B(n653), .ZN(G45) );
  NAND2_X1 U733 ( .A1(n654), .A2(n658), .ZN(n655) );
  XNOR2_X1 U734 ( .A(n655), .B(KEYINPUT116), .ZN(n656) );
  XNOR2_X1 U735 ( .A(G146), .B(n656), .ZN(G48) );
  NAND2_X1 U736 ( .A1(n395), .A2(n658), .ZN(n659) );
  XNOR2_X1 U737 ( .A(n659), .B(G113), .ZN(G15) );
  NAND2_X1 U738 ( .A1(n395), .A2(n660), .ZN(n661) );
  XNOR2_X1 U739 ( .A(n661), .B(G116), .ZN(G18) );
  XOR2_X1 U740 ( .A(G125), .B(KEYINPUT37), .Z(n662) );
  XNOR2_X1 U741 ( .A(n663), .B(n662), .ZN(G27) );
  XOR2_X1 U742 ( .A(G140), .B(KEYINPUT117), .Z(n664) );
  XNOR2_X1 U743 ( .A(n665), .B(n664), .ZN(G42) );
  NOR2_X1 U744 ( .A1(n692), .A2(n682), .ZN(n666) );
  XOR2_X1 U745 ( .A(KEYINPUT118), .B(KEYINPUT51), .Z(n680) );
  NAND2_X1 U746 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U747 ( .A(n669), .B(KEYINPUT50), .ZN(n676) );
  AND2_X1 U748 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U749 ( .A(KEYINPUT49), .B(n672), .Z(n673) );
  NOR2_X1 U750 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U751 ( .A1(n676), .A2(n675), .ZN(n678) );
  NAND2_X1 U752 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U753 ( .A(n680), .B(n679), .Z(n681) );
  NOR2_X1 U754 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U755 ( .A(KEYINPUT119), .B(n683), .Z(n695) );
  NOR2_X1 U756 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U757 ( .A1(n687), .A2(n686), .ZN(n691) );
  NOR2_X1 U758 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U759 ( .A1(n691), .A2(n690), .ZN(n693) );
  NOR2_X1 U760 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U761 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U762 ( .A(n696), .B(KEYINPUT52), .ZN(n697) );
  NOR2_X1 U763 ( .A1(n698), .A2(n697), .ZN(n704) );
  NOR2_X1 U764 ( .A1(n391), .A2(n699), .ZN(n701) );
  XNOR2_X1 U765 ( .A(KEYINPUT82), .B(KEYINPUT2), .ZN(n700) );
  NOR2_X1 U766 ( .A1(n701), .A2(n700), .ZN(n703) );
  NAND2_X1 U767 ( .A1(n733), .A2(G210), .ZN(n708) );
  NOR2_X1 U768 ( .A1(n709), .A2(n737), .ZN(n711) );
  XNOR2_X1 U769 ( .A(KEYINPUT88), .B(KEYINPUT56), .ZN(n710) );
  XNOR2_X1 U770 ( .A(n711), .B(n710), .ZN(G51) );
  BUF_X1 U771 ( .A(n712), .Z(n716) );
  XOR2_X1 U772 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n714) );
  XNOR2_X1 U773 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n713) );
  XNOR2_X1 U774 ( .A(n714), .B(n713), .ZN(n715) );
  NAND2_X1 U775 ( .A1(n733), .A2(G469), .ZN(n717) );
  XNOR2_X1 U776 ( .A(n717), .B(n718), .ZN(n719) );
  NOR2_X1 U777 ( .A1(n719), .A2(n737), .ZN(n720) );
  XNOR2_X1 U778 ( .A(n720), .B(KEYINPUT122), .ZN(G54) );
  NAND2_X1 U779 ( .A1(n733), .A2(G475), .ZN(n725) );
  INV_X1 U780 ( .A(n721), .ZN(n723) );
  XOR2_X1 U781 ( .A(KEYINPUT59), .B(KEYINPUT67), .Z(n722) );
  XNOR2_X1 U782 ( .A(n725), .B(n724), .ZN(n726) );
  XNOR2_X1 U783 ( .A(KEYINPUT68), .B(KEYINPUT60), .ZN(n727) );
  XNOR2_X1 U784 ( .A(n728), .B(n727), .ZN(G60) );
  XOR2_X1 U785 ( .A(n729), .B(KEYINPUT123), .Z(n731) );
  NAND2_X1 U786 ( .A1(n733), .A2(G478), .ZN(n730) );
  XNOR2_X1 U787 ( .A(n731), .B(n730), .ZN(n732) );
  NOR2_X1 U788 ( .A1(n737), .A2(n732), .ZN(G63) );
  XNOR2_X1 U789 ( .A(n734), .B(n735), .ZN(n736) );
  XNOR2_X1 U790 ( .A(KEYINPUT124), .B(n738), .ZN(G66) );
  XNOR2_X1 U791 ( .A(n396), .B(KEYINPUT126), .ZN(n741) );
  NAND2_X1 U792 ( .A1(n741), .A2(n740), .ZN(n750) );
  NAND2_X1 U793 ( .A1(G224), .A2(G953), .ZN(n742) );
  XNOR2_X1 U794 ( .A(n742), .B(KEYINPUT125), .ZN(n743) );
  XNOR2_X1 U795 ( .A(n743), .B(KEYINPUT61), .ZN(n744) );
  NOR2_X1 U796 ( .A1(n745), .A2(n744), .ZN(n748) );
  NOR2_X1 U797 ( .A1(G953), .A2(n391), .ZN(n747) );
  NOR2_X1 U798 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U799 ( .A(n750), .B(n749), .ZN(G69) );
  XOR2_X1 U800 ( .A(n752), .B(n751), .Z(n755) );
  XOR2_X1 U801 ( .A(n755), .B(n373), .Z(n754) );
  NAND2_X1 U802 ( .A1(n754), .A2(n347), .ZN(n759) );
  XNOR2_X1 U803 ( .A(G227), .B(n755), .ZN(n756) );
  NAND2_X1 U804 ( .A1(n756), .A2(G900), .ZN(n757) );
  NAND2_X1 U805 ( .A1(n757), .A2(G953), .ZN(n758) );
  NAND2_X1 U806 ( .A1(n759), .A2(n758), .ZN(n760) );
  XOR2_X1 U807 ( .A(KEYINPUT127), .B(n760), .Z(G72) );
  XOR2_X1 U808 ( .A(G134), .B(n761), .Z(G36) );
  XOR2_X1 U809 ( .A(G122), .B(n762), .Z(G24) );
  XNOR2_X1 U810 ( .A(G119), .B(n763), .ZN(G21) );
  XOR2_X1 U811 ( .A(n764), .B(G131), .Z(G33) );
  XOR2_X1 U812 ( .A(G137), .B(n765), .Z(G39) );
endmodule

