//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n547, new_n548, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n595,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n462), .A2(G137), .A3(new_n461), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n461), .A2(KEYINPUT66), .A3(G101), .A4(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(KEYINPUT67), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n466), .A2(new_n471), .A3(KEYINPUT67), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n465), .B1(new_n473), .B2(new_n474), .ZN(G160));
  NOR2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n461), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n477), .B2(new_n478), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  AND2_X1   g061(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n487));
  OAI211_X1 g062(.A(G138), .B(new_n461), .C1(new_n487), .C2(new_n476), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n462), .A2(KEYINPUT68), .A3(G138), .A4(new_n461), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n462), .A2(G126), .A3(G2105), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(G2104), .C1(G114), .C2(new_n461), .ZN(new_n495));
  AND2_X1   g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n488), .A2(new_n489), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n492), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT69), .B1(new_n501), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n506), .A2(G88), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(G50), .A3(G543), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n507), .B1(new_n502), .B2(new_n505), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OAI211_X1 g089(.A(new_n510), .B(new_n511), .C1(new_n513), .C2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  AND2_X1   g091(.A1(new_n512), .A2(new_n509), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G89), .ZN(new_n518));
  AND2_X1   g093(.A1(new_n509), .A2(G543), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n520), .A2(KEYINPUT7), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n519), .A2(G51), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n518), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g099(.A1(G63), .A2(G651), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n512), .A2(KEYINPUT70), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(KEYINPUT70), .B1(new_n512), .B2(new_n525), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n524), .A2(new_n528), .ZN(G168));
  AOI22_X1  g104(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n514), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n512), .A2(new_n509), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n509), .A2(G543), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n532), .A2(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n531), .A2(new_n536), .ZN(G171));
  AOI22_X1  g112(.A1(new_n512), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n538));
  OR3_X1    g113(.A1(new_n538), .A2(KEYINPUT71), .A3(new_n514), .ZN(new_n539));
  OAI21_X1  g114(.A(KEYINPUT71), .B1(new_n538), .B2(new_n514), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n517), .A2(G81), .B1(G43), .B2(new_n519), .ZN(new_n541));
  AND3_X1   g116(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT73), .ZN(new_n546));
  XOR2_X1   g121(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n547));
  XNOR2_X1  g122(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  XNOR2_X1  g124(.A(KEYINPUT74), .B(KEYINPUT9), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n519), .A2(G53), .A3(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT9), .ZN(new_n552));
  INV_X1    g127(.A(G53), .ZN(new_n553));
  OAI211_X1 g128(.A(KEYINPUT74), .B(new_n552), .C1(new_n535), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n512), .A2(G65), .ZN(new_n556));
  INV_X1    g131(.A(G78), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n557), .B2(new_n504), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n555), .B1(G651), .B2(new_n558), .ZN(new_n559));
  AND3_X1   g134(.A1(new_n512), .A2(G91), .A3(new_n509), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  INV_X1    g139(.A(G168), .ZN(G286));
  NAND4_X1  g140(.A1(new_n506), .A2(G87), .A3(new_n508), .A4(new_n509), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n509), .A2(G49), .A3(G543), .ZN(new_n567));
  AOI21_X1  g142(.A(G74), .B1(new_n506), .B2(new_n508), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n566), .B(new_n567), .C1(new_n568), .C2(new_n514), .ZN(G288));
  AND2_X1   g144(.A1(G73), .A2(G543), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(new_n512), .B2(G61), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n571), .A2(new_n514), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n506), .A2(G86), .A3(new_n508), .A4(new_n509), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n509), .A2(G48), .A3(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G305));
  AOI22_X1  g152(.A1(new_n517), .A2(G85), .B1(G47), .B2(new_n519), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n514), .B2(new_n579), .ZN(G290));
  NAND2_X1  g155(.A1(G301), .A2(G868), .ZN(new_n581));
  XOR2_X1   g156(.A(KEYINPUT76), .B(KEYINPUT10), .Z(new_n582));
  NAND3_X1  g157(.A1(new_n517), .A2(G92), .A3(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n582), .ZN(new_n584));
  INV_X1    g159(.A(G92), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n532), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n519), .A2(G54), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n512), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n589), .B2(new_n514), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n581), .B1(G868), .B2(new_n591), .ZN(G284));
  OAI21_X1  g167(.A(new_n581), .B1(G868), .B2(new_n591), .ZN(G321));
  INV_X1    g168(.A(G868), .ZN(new_n594));
  NAND2_X1  g169(.A1(G299), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n595), .B1(new_n594), .B2(G168), .ZN(G297));
  OAI21_X1  g171(.A(new_n595), .B1(new_n594), .B2(G168), .ZN(G280));
  INV_X1    g172(.A(G559), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n591), .B1(new_n598), .B2(G860), .ZN(G148));
  AND2_X1   g174(.A1(new_n583), .A2(new_n586), .ZN(new_n600));
  INV_X1    g175(.A(new_n590), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(G559), .ZN(new_n603));
  OR3_X1    g178(.A1(new_n603), .A2(KEYINPUT77), .A3(new_n594), .ZN(new_n604));
  OAI21_X1  g179(.A(KEYINPUT77), .B1(new_n603), .B2(new_n594), .ZN(new_n605));
  OAI211_X1 g180(.A(new_n604), .B(new_n605), .C1(G868), .C2(new_n542), .ZN(G323));
  XNOR2_X1  g181(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g182(.A1(new_n481), .A2(G135), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n479), .A2(G123), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n461), .A2(G111), .ZN(new_n610));
  OAI21_X1  g185(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n608), .B(new_n609), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(G2096), .Z(new_n613));
  NAND3_X1  g188(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT78), .B(KEYINPUT13), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(G2100), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n613), .A2(new_n619), .A3(new_n620), .ZN(G156));
  XNOR2_X1  g196(.A(G1341), .B(G1348), .ZN(new_n622));
  XOR2_X1   g197(.A(G2443), .B(G2446), .Z(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(KEYINPUT15), .B(G2435), .ZN(new_n625));
  INV_X1    g200(.A(G2438), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2427), .B(G2430), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT14), .ZN(new_n631));
  OAI21_X1  g206(.A(KEYINPUT79), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n625), .B(G2438), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(new_n628), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT79), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(new_n635), .A3(KEYINPUT14), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n633), .A2(new_n628), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n624), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  AOI211_X1 g215(.A(new_n638), .B(new_n623), .C1(new_n632), .C2(new_n636), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n622), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NOR3_X1   g217(.A1(new_n630), .A2(KEYINPUT79), .A3(new_n631), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n635), .B1(new_n634), .B2(KEYINPUT14), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n639), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(new_n623), .ZN(new_n646));
  INV_X1    g221(.A(new_n622), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n637), .A2(new_n639), .A3(new_n624), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n642), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(G14), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n651), .B1(new_n642), .B2(new_n649), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(G401));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT18), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2096), .B(G2100), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT80), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n661), .B(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT18), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n658), .A2(KEYINPUT17), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n656), .A2(new_n657), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n664), .B(new_n668), .Z(G227));
  XOR2_X1   g244(.A(G1991), .B(G1996), .Z(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT19), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT81), .B(KEYINPUT20), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n676), .A2(new_n677), .ZN(new_n682));
  OR3_X1    g257(.A1(new_n675), .A2(new_n678), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n675), .A2(new_n682), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n672), .B1(new_n681), .B2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  NOR3_X1   g262(.A1(new_n681), .A2(new_n685), .A3(new_n672), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n670), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1981), .B(G1986), .ZN(new_n690));
  INV_X1    g265(.A(new_n681), .ZN(new_n691));
  INV_X1    g266(.A(new_n685), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n691), .A2(new_n692), .A3(new_n671), .ZN(new_n693));
  INV_X1    g268(.A(new_n670), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n693), .A2(new_n694), .A3(new_n686), .ZN(new_n695));
  AND3_X1   g270(.A1(new_n689), .A2(new_n690), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n690), .B1(new_n689), .B2(new_n695), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(G229));
  INV_X1    g273(.A(G29), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G32), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT93), .B(KEYINPUT26), .Z(new_n701));
  NAND3_X1  g276(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n481), .A2(G141), .ZN(new_n706));
  INV_X1    g281(.A(G129), .ZN(new_n707));
  INV_X1    g282(.A(new_n479), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n700), .B1(new_n710), .B2(new_n699), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT27), .ZN(new_n712));
  INV_X1    g287(.A(G1996), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n699), .A2(G33), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n481), .A2(G139), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT25), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n462), .A2(G127), .ZN(new_n721));
  NAND2_X1  g296(.A1(G115), .A2(G2104), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n461), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT92), .ZN(new_n724));
  OR3_X1    g299(.A1(new_n720), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n720), .B2(new_n723), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n715), .B1(new_n728), .B2(new_n699), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G2072), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n699), .A2(G27), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G164), .B2(new_n699), .ZN(new_n732));
  INV_X1    g307(.A(G2078), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT31), .B(G11), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT94), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT30), .ZN(new_n737));
  AND2_X1   g312(.A1(new_n737), .A2(G28), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n699), .B1(new_n737), .B2(G28), .ZN(new_n739));
  OAI221_X1 g314(.A(new_n736), .B1(new_n738), .B2(new_n739), .C1(new_n612), .C2(new_n699), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT95), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n730), .A2(new_n734), .A3(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G16), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G5), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G171), .B2(new_n743), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT96), .B(G1961), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  NOR3_X1   g322(.A1(new_n714), .A2(new_n742), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n699), .A2(G35), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT97), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G162), .B2(new_n699), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G2090), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT99), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n743), .A2(G4), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n591), .B2(new_n743), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT88), .B(G1348), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n758), .B(new_n760), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n743), .A2(KEYINPUT83), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n743), .A2(KEYINPUT83), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n765), .A2(G20), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT100), .B(KEYINPUT23), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(G299), .B2(G16), .ZN(new_n769));
  INV_X1    g344(.A(G1956), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR3_X1   g346(.A1(new_n756), .A2(new_n761), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n765), .A2(G19), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT89), .Z(new_n774));
  NAND3_X1  g349(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(new_n764), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT90), .B(G1341), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n481), .A2(G140), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n479), .A2(G128), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n461), .A2(G116), .ZN(new_n781));
  OAI21_X1  g356(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n779), .B(new_n780), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G29), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n699), .A2(G26), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT28), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT91), .ZN(new_n788));
  INV_X1    g363(.A(G2067), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(G2084), .ZN(new_n791));
  NAND2_X1  g366(.A1(G160), .A2(G29), .ZN(new_n792));
  INV_X1    g367(.A(G34), .ZN(new_n793));
  AOI21_X1  g368(.A(G29), .B1(new_n793), .B2(KEYINPUT24), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(KEYINPUT24), .B2(new_n793), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  OAI22_X1  g371(.A1(new_n729), .A2(G2072), .B1(new_n791), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n743), .A2(G21), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G168), .B2(new_n743), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1966), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n796), .A2(new_n791), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n753), .B2(new_n754), .ZN(new_n802));
  NOR4_X1   g377(.A1(new_n790), .A2(new_n797), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n748), .A2(new_n772), .A3(new_n778), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n743), .A2(G6), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT32), .B(G1981), .ZN(new_n806));
  OAI211_X1 g381(.A(new_n805), .B(new_n806), .C1(new_n576), .C2(new_n743), .ZN(new_n807));
  INV_X1    g382(.A(new_n806), .ZN(new_n808));
  INV_X1    g383(.A(G61), .ZN(new_n809));
  AOI211_X1 g384(.A(new_n809), .B(new_n507), .C1(new_n502), .C2(new_n505), .ZN(new_n810));
  OAI21_X1  g385(.A(G651), .B1(new_n810), .B2(new_n570), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n573), .A2(new_n574), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n743), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n805), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n808), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT84), .B(G1971), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n506), .A2(G62), .A3(new_n508), .ZN(new_n818));
  NAND2_X1  g393(.A1(G75), .A2(G543), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n514), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n510), .A2(new_n511), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n820), .A2(new_n821), .A3(new_n765), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n764), .A2(G22), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n817), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n823), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n825), .B(new_n816), .C1(G303), .C2(new_n765), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n807), .A2(new_n815), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(G1976), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n566), .A2(new_n567), .ZN(new_n829));
  OAI21_X1  g404(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n743), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n743), .A2(G23), .ZN(new_n832));
  OAI21_X1  g407(.A(KEYINPUT33), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n832), .B1(G288), .B2(G16), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT33), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n828), .B1(new_n833), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n834), .A2(new_n835), .ZN(new_n838));
  AOI211_X1 g413(.A(KEYINPUT33), .B(new_n832), .C1(G288), .C2(G16), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n838), .A2(new_n839), .A3(G1976), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n827), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT85), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(G1976), .B1(new_n838), .B2(new_n839), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n833), .A2(new_n828), .A3(new_n836), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n846), .A2(KEYINPUT85), .A3(new_n827), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n843), .A2(KEYINPUT34), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(KEYINPUT34), .B1(new_n843), .B2(new_n847), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT86), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n699), .A2(G25), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n479), .A2(G119), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT82), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n854));
  INV_X1    g429(.A(G107), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n854), .B1(new_n855), .B2(G2105), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(G131), .B2(new_n481), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n853), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n851), .B1(new_n858), .B2(G29), .ZN(new_n859));
  XOR2_X1   g434(.A(KEYINPUT35), .B(G1991), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n764), .A2(G24), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(G290), .B2(new_n765), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(G1986), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(G1986), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n849), .A2(new_n850), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT34), .ZN(new_n870));
  AND3_X1   g445(.A1(new_n846), .A2(KEYINPUT85), .A3(new_n827), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT85), .B1(new_n846), .B2(new_n827), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n868), .ZN(new_n874));
  AOI21_X1  g449(.A(KEYINPUT86), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n848), .B1(new_n869), .B2(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(KEYINPUT87), .B(KEYINPUT36), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n848), .B(new_n877), .C1(new_n869), .C2(new_n875), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n804), .B1(new_n879), .B2(new_n880), .ZN(G311));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n879), .A2(new_n880), .ZN(new_n883));
  INV_X1    g458(.A(new_n804), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI211_X1 g460(.A(KEYINPUT101), .B(new_n804), .C1(new_n879), .C2(new_n880), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(G150));
  AOI22_X1  g462(.A1(new_n517), .A2(G93), .B1(G55), .B2(new_n519), .ZN(new_n888));
  AOI22_X1  g463(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n889), .A2(KEYINPUT102), .ZN(new_n890));
  OAI21_X1  g465(.A(G651), .B1(new_n889), .B2(KEYINPUT102), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(KEYINPUT103), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n894));
  OAI211_X1 g469(.A(new_n894), .B(new_n888), .C1(new_n890), .C2(new_n891), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n893), .A2(new_n542), .A3(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n775), .A2(KEYINPUT103), .A3(new_n892), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT38), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n591), .A2(G559), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n899), .B(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT39), .ZN(new_n902));
  AOI21_X1  g477(.A(G860), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(new_n902), .B2(new_n901), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n892), .A2(G860), .ZN(new_n905));
  XOR2_X1   g480(.A(new_n905), .B(KEYINPUT37), .Z(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(G145));
  NAND2_X1  g482(.A1(new_n481), .A2(G142), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n479), .A2(G130), .ZN(new_n909));
  OR2_X1    g484(.A1(G106), .A2(G2105), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n910), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n908), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT104), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n908), .A2(new_n909), .A3(new_n914), .A4(new_n911), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n615), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(new_n615), .A3(new_n915), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n917), .A2(new_n853), .A3(new_n857), .A4(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n918), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n858), .B1(new_n920), .B2(new_n916), .ZN(new_n921));
  AOI21_X1  g496(.A(KEYINPUT105), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n919), .A2(new_n921), .A3(KEYINPUT105), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n499), .A2(new_n783), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n499), .A2(new_n783), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n728), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n727), .A2(new_n925), .A3(new_n926), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(new_n710), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n710), .B1(new_n928), .B2(new_n929), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n923), .B(new_n924), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n932), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n919), .A2(new_n921), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n934), .A2(new_n930), .A3(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(G160), .B(new_n485), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(new_n612), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n933), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n924), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n934), .B(new_n930), .C1(new_n940), .C2(new_n922), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n938), .B1(new_n933), .B2(new_n941), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n939), .A2(new_n942), .A3(G37), .ZN(new_n943));
  XOR2_X1   g518(.A(new_n943), .B(KEYINPUT40), .Z(G395));
  AOI21_X1  g519(.A(KEYINPUT108), .B1(new_n892), .B2(new_n594), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n591), .A2(new_n562), .A3(new_n559), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n591), .B1(new_n562), .B2(new_n559), .ZN(new_n948));
  OAI21_X1  g523(.A(KEYINPUT41), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(G299), .A2(new_n602), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT41), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n946), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n896), .A2(new_n603), .A3(new_n897), .ZN(new_n954));
  INV_X1    g529(.A(new_n603), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n898), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n953), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n947), .A2(new_n948), .ZN(new_n958));
  INV_X1    g533(.A(new_n954), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n603), .B1(new_n896), .B2(new_n897), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n957), .A2(new_n961), .A3(KEYINPUT106), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n964), .B(new_n958), .C1(new_n959), .C2(new_n960), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(G290), .B(new_n576), .ZN(new_n967));
  INV_X1    g542(.A(G288), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(G303), .ZN(new_n969));
  OR2_X1    g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n967), .A2(new_n969), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n972), .B(KEYINPUT42), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n966), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n963), .B1(new_n962), .B2(new_n965), .ZN(new_n975));
  OAI21_X1  g550(.A(G868), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n962), .A2(new_n965), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT107), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n966), .B2(new_n973), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n945), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n974), .A2(new_n975), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n978), .A2(new_n966), .A3(new_n973), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n981), .A2(new_n982), .A3(KEYINPUT108), .A4(G868), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n980), .A2(new_n983), .ZN(G295));
  AND2_X1   g559(.A1(new_n980), .A2(new_n983), .ZN(G331));
  INV_X1    g560(.A(KEYINPUT43), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n987));
  NAND2_X1  g562(.A1(G171), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT109), .B1(new_n531), .B2(new_n536), .ZN(new_n989));
  NAND3_X1  g564(.A1(G286), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(G168), .A2(new_n987), .A3(G171), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n898), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n896), .A2(new_n897), .A3(new_n990), .A4(new_n991), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n953), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n993), .A2(new_n994), .A3(new_n958), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(new_n972), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G37), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n972), .B1(new_n996), .B2(new_n997), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n986), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n951), .B1(new_n950), .B2(new_n946), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1003), .B1(new_n1004), .B2(new_n952), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n958), .A2(KEYINPUT110), .A3(new_n951), .ZN(new_n1006));
  AOI22_X1  g581(.A1(new_n1005), .A2(new_n1006), .B1(new_n994), .B2(new_n993), .ZN(new_n1007));
  INV_X1    g582(.A(new_n997), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n970), .B(new_n971), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1009), .A2(KEYINPUT43), .A3(new_n999), .A4(new_n998), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1002), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT44), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT43), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1009), .A2(new_n986), .A3(new_n999), .A4(new_n998), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT44), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1012), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1016), .B1(new_n1002), .B2(new_n1010), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT44), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT111), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1019), .A2(new_n1022), .ZN(G397));
  XNOR2_X1  g598(.A(new_n783), .B(new_n789), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(new_n713), .B2(new_n710), .ZN(new_n1025));
  INV_X1    g600(.A(G1384), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n499), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n465), .ZN(new_n1030));
  INV_X1    g605(.A(new_n474), .ZN(new_n1031));
  OAI211_X1 g606(.A(G40), .B(new_n1030), .C1(new_n1031), .C2(new_n472), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1025), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n713), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n1035), .B(KEYINPUT113), .ZN(new_n1036));
  INV_X1    g611(.A(new_n710), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1034), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n860), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n858), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n853), .A2(new_n860), .A3(new_n857), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1038), .B1(new_n1033), .B2(new_n1042), .ZN(new_n1043));
  AND2_X1   g618(.A1(G290), .A2(G1986), .ZN(new_n1044));
  NOR2_X1   g619(.A1(G290), .A2(G1986), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1033), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g621(.A(new_n1046), .B(KEYINPUT112), .Z(new_n1047));
  AND2_X1   g622(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n498), .A2(new_n493), .A3(new_n495), .ZN(new_n1050));
  AOI21_X1  g625(.A(G1384), .B1(new_n1050), .B2(new_n492), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT45), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1032), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1029), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1049), .B1(new_n1054), .B2(G2078), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1032), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1056), .A2(KEYINPUT53), .A3(new_n733), .A4(new_n1052), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1032), .B1(new_n1027), .B2(KEYINPUT50), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT50), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n490), .A2(new_n491), .A3(KEYINPUT4), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n498), .A2(new_n493), .A3(new_n495), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1059), .B(new_n1026), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1058), .A2(new_n1062), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT125), .B(G1961), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1055), .A2(new_n1057), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(G171), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1055), .A2(new_n1065), .A3(G301), .A4(new_n1057), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT54), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G1966), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1054), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(G2084), .B2(new_n1063), .ZN(new_n1072));
  OAI21_X1  g647(.A(G8), .B1(new_n1072), .B2(G286), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1058), .A2(new_n1062), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1074), .A2(new_n791), .B1(new_n1070), .B2(new_n1054), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(G168), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT51), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G8), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1078), .B1(new_n1075), .B2(G168), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1069), .B1(new_n1077), .B2(new_n1081), .ZN(new_n1082));
  OR3_X1    g657(.A1(new_n572), .A2(G1981), .A3(new_n575), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT118), .B(G86), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n574), .B1(new_n532), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(G1981), .B1(new_n572), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT49), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1027), .A2(new_n1032), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1090), .A2(new_n1078), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1083), .A2(new_n1086), .A3(KEYINPUT49), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1089), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1091), .B1(new_n828), .B2(G288), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT52), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n968), .B2(G1976), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1093), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(KEYINPUT52), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT117), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT117), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1094), .A2(new_n1100), .A3(KEYINPUT52), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1097), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G1971), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1054), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT114), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT115), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n1063), .B2(G2090), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1058), .A2(KEYINPUT115), .A3(new_n754), .A4(new_n1062), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT114), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1054), .A2(new_n1109), .A3(new_n1103), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1105), .A2(new_n1107), .A3(new_n1108), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(G303), .A2(G8), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1112), .B(KEYINPUT55), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT116), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1113), .B(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1111), .A2(G8), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1062), .A2(KEYINPUT119), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n499), .A2(new_n1118), .A3(new_n1059), .A4(new_n1026), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1058), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1104), .B1(G2090), .B2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(G8), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(new_n1113), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1102), .A2(new_n1116), .A3(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1067), .A2(KEYINPUT54), .A3(new_n1068), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1082), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n558), .A2(G651), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1129), .A2(new_n551), .A3(new_n554), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n560), .B(KEYINPUT75), .ZN(new_n1131));
  OAI21_X1  g706(.A(KEYINPUT57), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT57), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n559), .A2(new_n562), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1121), .A2(new_n770), .ZN(new_n1137));
  XNOR2_X1  g712(.A(KEYINPUT56), .B(G2072), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1056), .A2(new_n1052), .A3(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1136), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(G1956), .B1(new_n1120), .B2(new_n1058), .ZN(new_n1141));
  AND4_X1   g716(.A1(new_n1052), .A2(new_n1029), .A3(new_n1053), .A4(new_n1138), .ZN(new_n1142));
  NOR3_X1   g717(.A1(new_n1141), .A2(new_n1142), .A3(new_n1135), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1128), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1063), .A2(new_n759), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1090), .A2(new_n789), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n600), .A2(KEYINPUT123), .A3(new_n601), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT123), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1148), .B1(new_n587), .B2(new_n590), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1145), .A2(KEYINPUT60), .A3(new_n1146), .A4(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT60), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n760), .B1(new_n1058), .B2(new_n1062), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1146), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1152), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1153), .A2(new_n1154), .A3(new_n1152), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1151), .B(new_n1155), .C1(new_n1156), .C2(new_n1149), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1137), .A2(new_n1136), .A3(new_n1139), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1135), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1158), .A2(KEYINPUT61), .A3(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1144), .A2(new_n1157), .A3(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1029), .A2(new_n1052), .A3(new_n713), .A4(new_n1053), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT121), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT121), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1056), .A2(new_n1164), .A3(new_n713), .A4(new_n1052), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1053), .A2(new_n1051), .ZN(new_n1166));
  XNOR2_X1  g741(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n1167));
  XNOR2_X1  g742(.A(new_n1167), .B(G1341), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1163), .A2(new_n1165), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT59), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1170), .A2(new_n1171), .A3(new_n542), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1171), .B1(new_n1170), .B2(new_n542), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1161), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n591), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1159), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n1158), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT120), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1178), .A2(KEYINPUT120), .A3(new_n1158), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g758(.A(KEYINPUT124), .B1(new_n1176), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1170), .A2(new_n542), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(KEYINPUT59), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(new_n1172), .ZN(new_n1187));
  NAND4_X1  g762(.A1(new_n1187), .A2(new_n1160), .A3(new_n1157), .A4(new_n1144), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT124), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1188), .A2(new_n1189), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1127), .B1(new_n1184), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1072), .A2(G286), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1080), .B1(new_n1079), .B2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1073), .A2(KEYINPUT51), .ZN(new_n1194));
  OAI21_X1  g769(.A(KEYINPUT62), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1077), .A2(new_n1196), .A3(new_n1081), .ZN(new_n1197));
  INV_X1    g772(.A(new_n1067), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1195), .A2(new_n1125), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  NOR3_X1   g774(.A1(new_n1075), .A2(new_n1078), .A3(G286), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1102), .A2(new_n1116), .A3(new_n1124), .A4(new_n1200), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT63), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AND2_X1   g778(.A1(new_n1200), .A2(KEYINPUT63), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1111), .A2(G8), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1205), .A2(new_n1113), .ZN(new_n1206));
  NAND4_X1  g781(.A1(new_n1204), .A2(new_n1206), .A3(new_n1116), .A4(new_n1102), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1203), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(new_n1116), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1093), .A2(new_n828), .A3(new_n968), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1210), .A2(new_n1083), .ZN(new_n1211));
  AOI22_X1  g786(.A1(new_n1209), .A2(new_n1102), .B1(new_n1091), .B2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1199), .A2(new_n1208), .A3(new_n1212), .ZN(new_n1213));
  OAI21_X1  g788(.A(new_n1048), .B1(new_n1191), .B2(new_n1213), .ZN(new_n1214));
  NOR2_X1   g789(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n783), .A2(G2067), .ZN(new_n1216));
  OAI21_X1  g791(.A(new_n1033), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n1033), .A2(new_n1045), .ZN(new_n1218));
  XNOR2_X1  g793(.A(new_n1218), .B(KEYINPUT48), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1043), .A2(new_n1219), .ZN(new_n1220));
  XNOR2_X1  g795(.A(new_n1036), .B(KEYINPUT46), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1024), .A2(new_n710), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1033), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  AND2_X1   g799(.A1(new_n1224), .A2(KEYINPUT47), .ZN(new_n1225));
  NOR2_X1   g800(.A1(new_n1224), .A2(KEYINPUT47), .ZN(new_n1226));
  OAI211_X1 g801(.A(new_n1217), .B(new_n1220), .C1(new_n1225), .C2(new_n1226), .ZN(new_n1227));
  INV_X1    g802(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1214), .A2(new_n1228), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g804(.A1(G227), .A2(new_n459), .ZN(new_n1231));
  OAI21_X1  g805(.A(new_n1231), .B1(new_n653), .B2(new_n654), .ZN(new_n1232));
  INV_X1    g806(.A(KEYINPUT126), .ZN(new_n1233));
  AOI21_X1  g807(.A(G229), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g808(.A(new_n1234), .B1(new_n1233), .B2(new_n1232), .ZN(new_n1235));
  NOR2_X1   g809(.A1(new_n1235), .A2(new_n943), .ZN(new_n1236));
  AND3_X1   g810(.A1(new_n1236), .A2(KEYINPUT127), .A3(new_n1015), .ZN(new_n1237));
  AOI21_X1  g811(.A(KEYINPUT127), .B1(new_n1236), .B2(new_n1015), .ZN(new_n1238));
  NOR2_X1   g812(.A1(new_n1237), .A2(new_n1238), .ZN(G308));
  NAND2_X1  g813(.A1(new_n1236), .A2(new_n1015), .ZN(G225));
endmodule


