

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593;

  XOR2_X2 U326 ( .A(n457), .B(KEYINPUT28), .Z(n529) );
  XNOR2_X2 U327 ( .A(KEYINPUT104), .B(n297), .ZN(n504) );
  XOR2_X1 U328 ( .A(KEYINPUT92), .B(n465), .Z(n575) );
  XOR2_X1 U329 ( .A(KEYINPUT40), .B(n505), .Z(n294) );
  XOR2_X1 U330 ( .A(n426), .B(n425), .Z(n295) );
  NOR2_X1 U331 ( .A1(n460), .A2(n451), .ZN(n296) );
  XOR2_X1 U332 ( .A(n478), .B(KEYINPUT38), .Z(n297) );
  XOR2_X1 U333 ( .A(G50GAT), .B(G162GAT), .Z(n424) );
  INV_X1 U334 ( .A(n357), .ZN(n358) );
  XNOR2_X1 U335 ( .A(n359), .B(n358), .ZN(n360) );
  INV_X1 U336 ( .A(KEYINPUT74), .ZN(n364) );
  XNOR2_X1 U337 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U338 ( .A(n448), .B(n432), .Z(n460) );
  XNOR2_X1 U339 ( .A(n559), .B(n364), .ZN(n482) );
  INV_X1 U340 ( .A(n482), .ZN(n454) );
  XNOR2_X1 U341 ( .A(n482), .B(KEYINPUT36), .ZN(n591) );
  XOR2_X1 U342 ( .A(n582), .B(KEYINPUT41), .Z(n565) );
  INV_X1 U343 ( .A(KEYINPUT106), .ZN(n479) );
  XNOR2_X1 U344 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n455) );
  XNOR2_X1 U345 ( .A(n479), .B(G50GAT), .ZN(n480) );
  XNOR2_X1 U346 ( .A(n456), .B(n455), .ZN(G1351GAT) );
  XNOR2_X1 U347 ( .A(n481), .B(n480), .ZN(G1331GAT) );
  XOR2_X1 U348 ( .A(G134GAT), .B(G43GAT), .Z(n299) );
  NAND2_X1 U349 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U350 ( .A(n299), .B(n298), .ZN(n302) );
  XOR2_X1 U351 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n301) );
  XNOR2_X1 U352 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n301), .B(n300), .ZN(n323) );
  XOR2_X1 U354 ( .A(n302), .B(n323), .Z(n310) );
  XOR2_X1 U355 ( .A(KEYINPUT83), .B(KEYINPUT84), .Z(n304) );
  XNOR2_X1 U356 ( .A(G99GAT), .B(G190GAT), .ZN(n303) );
  XNOR2_X1 U357 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U358 ( .A(KEYINPUT20), .B(G176GAT), .Z(n306) );
  XNOR2_X1 U359 ( .A(G15GAT), .B(G183GAT), .ZN(n305) );
  XNOR2_X1 U360 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U362 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U363 ( .A(n311), .B(G71GAT), .Z(n315) );
  XOR2_X1 U364 ( .A(G127GAT), .B(KEYINPUT82), .Z(n313) );
  XNOR2_X1 U365 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n313), .B(n312), .ZN(n440) );
  XNOR2_X1 U367 ( .A(n440), .B(G120GAT), .ZN(n314) );
  XNOR2_X2 U368 ( .A(n315), .B(n314), .ZN(n531) );
  XOR2_X1 U369 ( .A(G176GAT), .B(G64GAT), .Z(n332) );
  XNOR2_X1 U370 ( .A(G8GAT), .B(G183GAT), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n316), .B(KEYINPUT75), .ZN(n376) );
  XOR2_X1 U372 ( .A(n332), .B(n376), .Z(n318) );
  XNOR2_X1 U373 ( .A(G204GAT), .B(KEYINPUT94), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n318), .B(n317), .ZN(n327) );
  XOR2_X1 U375 ( .A(KEYINPUT96), .B(KEYINPUT93), .Z(n320) );
  NAND2_X1 U376 ( .A1(G226GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U377 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U378 ( .A(n321), .B(KEYINPUT95), .Z(n325) );
  XNOR2_X1 U379 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n322) );
  XNOR2_X1 U380 ( .A(n322), .B(G211GAT), .ZN(n419) );
  XNOR2_X1 U381 ( .A(n323), .B(n419), .ZN(n324) );
  XNOR2_X1 U382 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U383 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U384 ( .A(G92GAT), .B(KEYINPUT72), .Z(n329) );
  XNOR2_X1 U385 ( .A(G190GAT), .B(G218GAT), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U387 ( .A(G36GAT), .B(n330), .Z(n347) );
  XOR2_X1 U388 ( .A(n331), .B(n347), .Z(n520) );
  XOR2_X1 U389 ( .A(G99GAT), .B(G106GAT), .Z(n357) );
  XOR2_X1 U390 ( .A(n357), .B(n332), .Z(n334) );
  NAND2_X1 U391 ( .A1(G230GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U392 ( .A(n334), .B(n333), .ZN(n345) );
  XOR2_X1 U393 ( .A(KEYINPUT31), .B(KEYINPUT70), .Z(n340) );
  XNOR2_X1 U394 ( .A(G120GAT), .B(G148GAT), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n335), .B(G57GAT), .ZN(n443) );
  XOR2_X1 U396 ( .A(KEYINPUT32), .B(KEYINPUT68), .Z(n337) );
  XNOR2_X1 U397 ( .A(KEYINPUT69), .B(KEYINPUT33), .ZN(n336) );
  XNOR2_X1 U398 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U399 ( .A(n443), .B(n338), .ZN(n339) );
  XNOR2_X1 U400 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U401 ( .A(G71GAT), .B(KEYINPUT13), .Z(n367) );
  XOR2_X1 U402 ( .A(n341), .B(n367), .Z(n343) );
  XNOR2_X1 U403 ( .A(G85GAT), .B(G92GAT), .ZN(n342) );
  XNOR2_X1 U404 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U405 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U406 ( .A(G204GAT), .B(G78GAT), .ZN(n423) );
  XOR2_X1 U407 ( .A(n346), .B(n423), .Z(n477) );
  INV_X1 U408 ( .A(n477), .ZN(n582) );
  INV_X1 U409 ( .A(n347), .ZN(n351) );
  XOR2_X1 U410 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n349) );
  XNOR2_X1 U411 ( .A(KEYINPUT9), .B(KEYINPUT11), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U413 ( .A(n351), .B(n350), .Z(n363) );
  XNOR2_X1 U414 ( .A(G29GAT), .B(G134GAT), .ZN(n352) );
  XNOR2_X1 U415 ( .A(n352), .B(G85GAT), .ZN(n439) );
  INV_X1 U416 ( .A(KEYINPUT73), .ZN(n353) );
  XNOR2_X1 U417 ( .A(n439), .B(n353), .ZN(n355) );
  NAND2_X1 U418 ( .A1(G232GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n355), .B(n354), .ZN(n361) );
  XNOR2_X1 U420 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n356) );
  XNOR2_X1 U421 ( .A(n356), .B(KEYINPUT7), .ZN(n396) );
  XNOR2_X1 U422 ( .A(n396), .B(n424), .ZN(n359) );
  XOR2_X1 U423 ( .A(n363), .B(n362), .Z(n559) );
  XOR2_X1 U424 ( .A(G64GAT), .B(G57GAT), .Z(n366) );
  XNOR2_X1 U425 ( .A(G155GAT), .B(G78GAT), .ZN(n365) );
  XNOR2_X1 U426 ( .A(n366), .B(n365), .ZN(n368) );
  XOR2_X1 U427 ( .A(n368), .B(n367), .Z(n370) );
  XNOR2_X1 U428 ( .A(G127GAT), .B(G211GAT), .ZN(n369) );
  XNOR2_X1 U429 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U430 ( .A(KEYINPUT79), .B(KEYINPUT78), .Z(n372) );
  XNOR2_X1 U431 ( .A(KEYINPUT77), .B(KEYINPUT15), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U433 ( .A(n374), .B(n373), .Z(n378) );
  XNOR2_X1 U434 ( .A(G22GAT), .B(G15GAT), .ZN(n375) );
  XNOR2_X1 U435 ( .A(n375), .B(G1GAT), .ZN(n393) );
  XNOR2_X1 U436 ( .A(n393), .B(n376), .ZN(n377) );
  XNOR2_X1 U437 ( .A(n378), .B(n377), .ZN(n383) );
  XOR2_X1 U438 ( .A(KEYINPUT76), .B(KEYINPUT12), .Z(n380) );
  NAND2_X1 U439 ( .A1(G231GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U440 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U441 ( .A(KEYINPUT14), .B(n381), .Z(n382) );
  XOR2_X1 U442 ( .A(n383), .B(n382), .Z(n585) );
  INV_X1 U443 ( .A(n585), .ZN(n556) );
  NOR2_X1 U444 ( .A1(n591), .A2(n556), .ZN(n384) );
  XOR2_X1 U445 ( .A(KEYINPUT45), .B(n384), .Z(n385) );
  NOR2_X1 U446 ( .A1(n582), .A2(n385), .ZN(n386) );
  XNOR2_X1 U447 ( .A(KEYINPUT112), .B(n386), .ZN(n404) );
  XOR2_X1 U448 ( .A(G8GAT), .B(G113GAT), .Z(n388) );
  XNOR2_X1 U449 ( .A(G169GAT), .B(G197GAT), .ZN(n387) );
  XNOR2_X1 U450 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U451 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n390) );
  XNOR2_X1 U452 ( .A(KEYINPUT66), .B(KEYINPUT65), .ZN(n389) );
  XNOR2_X1 U453 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U454 ( .A(n392), .B(n391), .ZN(n403) );
  XOR2_X1 U455 ( .A(G50GAT), .B(G29GAT), .Z(n395) );
  XNOR2_X1 U456 ( .A(G141GAT), .B(n393), .ZN(n394) );
  XNOR2_X1 U457 ( .A(n395), .B(n394), .ZN(n401) );
  XOR2_X1 U458 ( .A(n396), .B(KEYINPUT67), .Z(n398) );
  NAND2_X1 U459 ( .A1(G229GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U460 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U461 ( .A(n399), .B(G36GAT), .Z(n400) );
  XNOR2_X1 U462 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U463 ( .A(n403), .B(n402), .Z(n547) );
  AND2_X1 U464 ( .A1(n404), .A2(n547), .ZN(n411) );
  XOR2_X1 U465 ( .A(KEYINPUT46), .B(KEYINPUT111), .Z(n406) );
  INV_X1 U466 ( .A(n547), .ZN(n579) );
  NAND2_X1 U467 ( .A1(n565), .A2(n579), .ZN(n405) );
  XNOR2_X1 U468 ( .A(n406), .B(n405), .ZN(n407) );
  NAND2_X1 U469 ( .A1(n407), .A2(n556), .ZN(n408) );
  NOR2_X1 U470 ( .A1(n559), .A2(n408), .ZN(n409) );
  XOR2_X1 U471 ( .A(KEYINPUT47), .B(n409), .Z(n410) );
  NOR2_X1 U472 ( .A1(n411), .A2(n410), .ZN(n412) );
  XNOR2_X1 U473 ( .A(n412), .B(KEYINPUT48), .ZN(n528) );
  NOR2_X1 U474 ( .A1(n520), .A2(n528), .ZN(n413) );
  XNOR2_X1 U475 ( .A(KEYINPUT54), .B(n413), .ZN(n576) );
  XOR2_X1 U476 ( .A(KEYINPUT2), .B(KEYINPUT86), .Z(n415) );
  XNOR2_X1 U477 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n414) );
  XNOR2_X1 U478 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U479 ( .A(G141GAT), .B(n416), .Z(n448) );
  XOR2_X1 U480 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n418) );
  XNOR2_X1 U481 ( .A(G22GAT), .B(KEYINPUT24), .ZN(n417) );
  XNOR2_X1 U482 ( .A(n418), .B(n417), .ZN(n430) );
  XNOR2_X1 U483 ( .A(n419), .B(G148GAT), .ZN(n421) );
  AND2_X1 U484 ( .A1(G228GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U485 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U486 ( .A(n422), .B(G218GAT), .ZN(n428) );
  XOR2_X1 U487 ( .A(KEYINPUT23), .B(KEYINPUT85), .Z(n426) );
  XOR2_X1 U488 ( .A(n424), .B(n423), .Z(n425) );
  XNOR2_X1 U489 ( .A(n295), .B(G106GAT), .ZN(n427) );
  XNOR2_X1 U490 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U491 ( .A(n430), .B(n429), .ZN(n431) );
  INV_X1 U492 ( .A(n431), .ZN(n432) );
  XOR2_X1 U493 ( .A(KEYINPUT4), .B(KEYINPUT89), .Z(n434) );
  XNOR2_X1 U494 ( .A(KEYINPUT90), .B(KEYINPUT6), .ZN(n433) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U496 ( .A(KEYINPUT91), .B(KEYINPUT1), .Z(n436) );
  XNOR2_X1 U497 ( .A(KEYINPUT5), .B(KEYINPUT88), .ZN(n435) );
  XNOR2_X1 U498 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U499 ( .A(n438), .B(n437), .Z(n442) );
  XNOR2_X1 U500 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U501 ( .A(n442), .B(n441), .ZN(n447) );
  XOR2_X1 U502 ( .A(n443), .B(G162GAT), .Z(n445) );
  NAND2_X1 U503 ( .A1(G225GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U504 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U505 ( .A(n447), .B(n446), .Z(n450) );
  XNOR2_X1 U506 ( .A(G1GAT), .B(n448), .ZN(n449) );
  XNOR2_X1 U507 ( .A(n450), .B(n449), .ZN(n465) );
  INV_X1 U508 ( .A(n575), .ZN(n451) );
  AND2_X1 U509 ( .A1(n576), .A2(n296), .ZN(n452) );
  XNOR2_X1 U510 ( .A(n452), .B(KEYINPUT55), .ZN(n453) );
  NOR2_X2 U511 ( .A1(n531), .A2(n453), .ZN(n570) );
  NAND2_X1 U512 ( .A1(n570), .A2(n454), .ZN(n456) );
  XNOR2_X1 U513 ( .A(n460), .B(KEYINPUT64), .ZN(n457) );
  NAND2_X1 U514 ( .A1(n460), .A2(n531), .ZN(n458) );
  XNOR2_X1 U515 ( .A(n458), .B(KEYINPUT26), .ZN(n578) );
  XNOR2_X1 U516 ( .A(KEYINPUT27), .B(n520), .ZN(n467) );
  NOR2_X1 U517 ( .A1(n578), .A2(n467), .ZN(n463) );
  NOR2_X1 U518 ( .A1(n531), .A2(n520), .ZN(n459) );
  NOR2_X1 U519 ( .A1(n460), .A2(n459), .ZN(n461) );
  XOR2_X1 U520 ( .A(KEYINPUT25), .B(n461), .Z(n462) );
  NOR2_X1 U521 ( .A1(n463), .A2(n462), .ZN(n464) );
  NOR2_X1 U522 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U523 ( .A(n466), .B(KEYINPUT98), .ZN(n473) );
  INV_X1 U524 ( .A(n529), .ZN(n471) );
  NOR2_X1 U525 ( .A1(n575), .A2(n467), .ZN(n468) );
  XNOR2_X1 U526 ( .A(KEYINPUT97), .B(n468), .ZN(n527) );
  INV_X1 U527 ( .A(n527), .ZN(n469) );
  NAND2_X1 U528 ( .A1(n469), .A2(n531), .ZN(n470) );
  NOR2_X1 U529 ( .A1(n471), .A2(n470), .ZN(n472) );
  NOR2_X1 U530 ( .A1(n473), .A2(n472), .ZN(n474) );
  XNOR2_X1 U531 ( .A(n474), .B(KEYINPUT99), .ZN(n486) );
  NAND2_X1 U532 ( .A1(n486), .A2(n556), .ZN(n475) );
  NOR2_X1 U533 ( .A1(n475), .A2(n591), .ZN(n476) );
  XNOR2_X1 U534 ( .A(n476), .B(KEYINPUT37), .ZN(n516) );
  NAND2_X1 U535 ( .A1(n477), .A2(n579), .ZN(n489) );
  NOR2_X1 U536 ( .A1(n516), .A2(n489), .ZN(n478) );
  NOR2_X1 U537 ( .A1(n529), .A2(n504), .ZN(n481) );
  NAND2_X1 U538 ( .A1(n482), .A2(n585), .ZN(n485) );
  XNOR2_X1 U539 ( .A(KEYINPUT80), .B(KEYINPUT16), .ZN(n483) );
  XNOR2_X1 U540 ( .A(n483), .B(KEYINPUT81), .ZN(n484) );
  XNOR2_X1 U541 ( .A(n485), .B(n484), .ZN(n487) );
  NAND2_X1 U542 ( .A1(n487), .A2(n486), .ZN(n488) );
  XNOR2_X1 U543 ( .A(KEYINPUT100), .B(n488), .ZN(n508) );
  OR2_X1 U544 ( .A1(n508), .A2(n489), .ZN(n498) );
  NOR2_X1 U545 ( .A1(n575), .A2(n498), .ZN(n494) );
  XOR2_X1 U546 ( .A(KEYINPUT34), .B(KEYINPUT103), .Z(n491) );
  XNOR2_X1 U547 ( .A(G1GAT), .B(KEYINPUT102), .ZN(n490) );
  XNOR2_X1 U548 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U549 ( .A(KEYINPUT101), .B(n492), .ZN(n493) );
  XNOR2_X1 U550 ( .A(n494), .B(n493), .ZN(G1324GAT) );
  NOR2_X1 U551 ( .A1(n520), .A2(n498), .ZN(n495) );
  XOR2_X1 U552 ( .A(G8GAT), .B(n495), .Z(G1325GAT) );
  NOR2_X1 U553 ( .A1(n531), .A2(n498), .ZN(n497) );
  XNOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n496) );
  XNOR2_X1 U555 ( .A(n497), .B(n496), .ZN(G1326GAT) );
  NOR2_X1 U556 ( .A1(n529), .A2(n498), .ZN(n499) );
  XOR2_X1 U557 ( .A(G22GAT), .B(n499), .Z(G1327GAT) );
  NOR2_X1 U558 ( .A1(n575), .A2(n504), .ZN(n500) );
  XNOR2_X1 U559 ( .A(n500), .B(KEYINPUT39), .ZN(n501) );
  XNOR2_X1 U560 ( .A(G29GAT), .B(n501), .ZN(G1328GAT) );
  NOR2_X1 U561 ( .A1(n520), .A2(n504), .ZN(n503) );
  XNOR2_X1 U562 ( .A(G36GAT), .B(KEYINPUT105), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n503), .B(n502), .ZN(G1329GAT) );
  NOR2_X1 U564 ( .A1(n531), .A2(n504), .ZN(n505) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n294), .ZN(G1330GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n507) );
  XNOR2_X1 U567 ( .A(G57GAT), .B(KEYINPUT107), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n507), .B(n506), .ZN(n510) );
  NAND2_X1 U569 ( .A1(n547), .A2(n565), .ZN(n517) );
  OR2_X1 U570 ( .A1(n508), .A2(n517), .ZN(n513) );
  NOR2_X1 U571 ( .A1(n575), .A2(n513), .ZN(n509) );
  XOR2_X1 U572 ( .A(n510), .B(n509), .Z(G1332GAT) );
  NOR2_X1 U573 ( .A1(n520), .A2(n513), .ZN(n511) );
  XOR2_X1 U574 ( .A(G64GAT), .B(n511), .Z(G1333GAT) );
  NOR2_X1 U575 ( .A1(n531), .A2(n513), .ZN(n512) );
  XOR2_X1 U576 ( .A(G71GAT), .B(n512), .Z(G1334GAT) );
  NOR2_X1 U577 ( .A1(n529), .A2(n513), .ZN(n515) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(G1335GAT) );
  NOR2_X1 U580 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n518), .B(KEYINPUT109), .ZN(n524) );
  NOR2_X1 U582 ( .A1(n575), .A2(n524), .ZN(n519) );
  XOR2_X1 U583 ( .A(G85GAT), .B(n519), .Z(G1336GAT) );
  NOR2_X1 U584 ( .A1(n520), .A2(n524), .ZN(n521) );
  XOR2_X1 U585 ( .A(G92GAT), .B(n521), .Z(G1337GAT) );
  NOR2_X1 U586 ( .A1(n531), .A2(n524), .ZN(n522) );
  XOR2_X1 U587 ( .A(KEYINPUT110), .B(n522), .Z(n523) );
  XNOR2_X1 U588 ( .A(G99GAT), .B(n523), .ZN(G1338GAT) );
  NOR2_X1 U589 ( .A1(n529), .A2(n524), .ZN(n525) );
  XOR2_X1 U590 ( .A(KEYINPUT44), .B(n525), .Z(n526) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  XOR2_X1 U592 ( .A(G113GAT), .B(KEYINPUT113), .Z(n533) );
  NOR2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n546) );
  NAND2_X1 U594 ( .A1(n546), .A2(n529), .ZN(n530) );
  NOR2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n540) );
  NAND2_X1 U596 ( .A1(n540), .A2(n579), .ZN(n532) );
  XNOR2_X1 U597 ( .A(n533), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U599 ( .A1(n540), .A2(n565), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(KEYINPUT114), .ZN(n539) );
  XOR2_X1 U602 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n537) );
  NAND2_X1 U603 ( .A1(n540), .A2(n585), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n542) );
  NAND2_X1 U607 ( .A1(n540), .A2(n454), .ZN(n541) );
  XNOR2_X1 U608 ( .A(n542), .B(n541), .ZN(n544) );
  XOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT116), .Z(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  INV_X1 U611 ( .A(n578), .ZN(n545) );
  NAND2_X1 U612 ( .A1(n546), .A2(n545), .ZN(n560) );
  NOR2_X1 U613 ( .A1(n547), .A2(n560), .ZN(n548) );
  XOR2_X1 U614 ( .A(G141GAT), .B(n548), .Z(n549) );
  XNOR2_X1 U615 ( .A(KEYINPUT118), .B(n549), .ZN(G1344GAT) );
  INV_X1 U616 ( .A(n565), .ZN(n550) );
  NOR2_X1 U617 ( .A1(n550), .A2(n560), .ZN(n555) );
  XOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n552) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(KEYINPUT119), .B(n553), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  NOR2_X1 U623 ( .A1(n556), .A2(n560), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1346GAT) );
  INV_X1 U626 ( .A(n559), .ZN(n561) );
  NOR2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U628 ( .A(G162GAT), .B(n562), .Z(G1347GAT) );
  NAND2_X1 U629 ( .A1(n579), .A2(n570), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(KEYINPUT122), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U632 ( .A1(n570), .A2(n565), .ZN(n567) );
  XOR2_X1 U633 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n569) );
  XOR2_X1 U635 ( .A(G176GAT), .B(KEYINPUT56), .Z(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  NAND2_X1 U637 ( .A1(n570), .A2(n585), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n573) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n572) );
  XNOR2_X1 U641 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U642 ( .A(KEYINPUT59), .B(n574), .Z(n581) );
  NAND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n589) );
  NAND2_X1 U645 ( .A1(n589), .A2(n579), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  NAND2_X1 U648 ( .A1(n589), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NAND2_X1 U650 ( .A1(n589), .A2(n585), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT126), .B(KEYINPUT62), .Z(n588) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n587) );
  XNOR2_X1 U654 ( .A(n588), .B(n587), .ZN(n593) );
  INV_X1 U655 ( .A(n589), .ZN(n590) );
  NOR2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U657 ( .A(n593), .B(n592), .Z(G1355GAT) );
endmodule

