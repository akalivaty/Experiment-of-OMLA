

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U319 ( .A(n344), .B(n343), .ZN(n346) );
  OR2_X1 U320 ( .A1(n462), .A2(n461), .ZN(n463) );
  XNOR2_X1 U321 ( .A(n311), .B(n310), .ZN(n336) );
  NOR2_X1 U322 ( .A1(n394), .A2(n393), .ZN(n395) );
  XNOR2_X1 U323 ( .A(n409), .B(n290), .ZN(n410) );
  INV_X1 U324 ( .A(KEYINPUT55), .ZN(n471) );
  NOR2_X1 U325 ( .A1(n470), .A2(n565), .ZN(n472) );
  XOR2_X1 U326 ( .A(n429), .B(n428), .Z(n287) );
  XOR2_X1 U327 ( .A(G43GAT), .B(G50GAT), .Z(n288) );
  XOR2_X1 U328 ( .A(n372), .B(n402), .Z(n289) );
  XOR2_X1 U329 ( .A(n408), .B(n407), .Z(n290) );
  XOR2_X1 U330 ( .A(n463), .B(KEYINPUT47), .Z(n291) );
  OR2_X1 U331 ( .A1(n456), .A2(n459), .ZN(n292) );
  NOR2_X1 U332 ( .A1(n529), .A2(n526), .ZN(n380) );
  XNOR2_X1 U333 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U334 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U335 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U336 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U337 ( .A(n430), .B(n287), .ZN(n431) );
  NAND2_X1 U338 ( .A1(n292), .A2(n291), .ZN(n464) );
  INV_X1 U339 ( .A(KEYINPUT97), .ZN(n374) );
  XNOR2_X1 U340 ( .A(n432), .B(n431), .ZN(n456) );
  XNOR2_X1 U341 ( .A(n464), .B(KEYINPUT48), .ZN(n533) );
  XNOR2_X1 U342 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U343 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U344 ( .A(n377), .B(n376), .ZN(n378) );
  INV_X1 U345 ( .A(KEYINPUT44), .ZN(n453) );
  XNOR2_X1 U346 ( .A(n480), .B(n479), .ZN(n508) );
  XNOR2_X1 U347 ( .A(n483), .B(G190GAT), .ZN(n484) );
  XNOR2_X1 U348 ( .A(n453), .B(G106GAT), .ZN(n454) );
  XNOR2_X1 U349 ( .A(n450), .B(G85GAT), .ZN(n451) );
  XNOR2_X1 U350 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n481) );
  XNOR2_X1 U351 ( .A(n485), .B(n484), .ZN(G1351GAT) );
  XNOR2_X1 U352 ( .A(n452), .B(n451), .ZN(G1336GAT) );
  XOR2_X1 U353 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n294) );
  XNOR2_X1 U354 ( .A(G85GAT), .B(KEYINPUT95), .ZN(n293) );
  XNOR2_X1 U355 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U356 ( .A(G120GAT), .B(G57GAT), .Z(n422) );
  XOR2_X1 U357 ( .A(n295), .B(n422), .Z(n300) );
  XOR2_X1 U358 ( .A(KEYINPUT0), .B(KEYINPUT84), .Z(n297) );
  XNOR2_X1 U359 ( .A(G127GAT), .B(G113GAT), .ZN(n296) );
  XNOR2_X1 U360 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U361 ( .A(KEYINPUT83), .B(n298), .Z(n365) );
  XOR2_X1 U362 ( .A(G29GAT), .B(G134GAT), .Z(n408) );
  XNOR2_X1 U363 ( .A(n365), .B(n408), .ZN(n299) );
  XNOR2_X1 U364 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U365 ( .A(KEYINPUT6), .B(G1GAT), .Z(n302) );
  NAND2_X1 U366 ( .A1(G225GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U367 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U368 ( .A(n304), .B(n303), .Z(n313) );
  XOR2_X1 U369 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n306) );
  XNOR2_X1 U370 ( .A(KEYINPUT90), .B(KEYINPUT2), .ZN(n305) );
  XNOR2_X1 U371 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U372 ( .A(n307), .B(G148GAT), .Z(n311) );
  XNOR2_X1 U373 ( .A(G155GAT), .B(G141GAT), .ZN(n309) );
  XNOR2_X1 U374 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n308) );
  XNOR2_X1 U375 ( .A(n336), .B(KEYINPUT4), .ZN(n312) );
  XNOR2_X1 U376 ( .A(n313), .B(n312), .ZN(n387) );
  XNOR2_X1 U377 ( .A(KEYINPUT96), .B(n387), .ZN(n514) );
  XOR2_X1 U378 ( .A(KEYINPUT13), .B(G71GAT), .Z(n421) );
  XOR2_X1 U379 ( .A(G8GAT), .B(G57GAT), .Z(n315) );
  XNOR2_X1 U380 ( .A(G155GAT), .B(G127GAT), .ZN(n314) );
  XNOR2_X1 U381 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U382 ( .A(n421), .B(n316), .Z(n318) );
  NAND2_X1 U383 ( .A1(G231GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U384 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U385 ( .A(n319), .B(KEYINPUT82), .Z(n322) );
  XNOR2_X1 U386 ( .A(G1GAT), .B(G22GAT), .ZN(n320) );
  XNOR2_X1 U387 ( .A(n320), .B(G15GAT), .ZN(n440) );
  XNOR2_X1 U388 ( .A(n440), .B(KEYINPUT81), .ZN(n321) );
  XNOR2_X1 U389 ( .A(n322), .B(n321), .ZN(n330) );
  XOR2_X1 U390 ( .A(KEYINPUT80), .B(G183GAT), .Z(n324) );
  XNOR2_X1 U391 ( .A(G64GAT), .B(G211GAT), .ZN(n323) );
  XNOR2_X1 U392 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U393 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n326) );
  XNOR2_X1 U394 ( .A(G78GAT), .B(KEYINPUT15), .ZN(n325) );
  XNOR2_X1 U395 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U396 ( .A(n328), .B(n327), .Z(n329) );
  XOR2_X1 U397 ( .A(n330), .B(n329), .Z(n575) );
  INV_X1 U398 ( .A(n575), .ZN(n563) );
  XOR2_X1 U399 ( .A(KEYINPUT89), .B(G197GAT), .Z(n332) );
  XNOR2_X1 U400 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n331) );
  XNOR2_X1 U401 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U402 ( .A(G211GAT), .B(n333), .Z(n371) );
  XOR2_X1 U403 ( .A(KEYINPUT70), .B(KEYINPUT71), .Z(n335) );
  XNOR2_X1 U404 ( .A(G106GAT), .B(G78GAT), .ZN(n334) );
  XNOR2_X1 U405 ( .A(n335), .B(n334), .ZN(n419) );
  XNOR2_X1 U406 ( .A(n336), .B(n419), .ZN(n344) );
  XOR2_X1 U407 ( .A(KEYINPUT94), .B(KEYINPUT22), .Z(n338) );
  XNOR2_X1 U408 ( .A(G22GAT), .B(KEYINPUT23), .ZN(n337) );
  XNOR2_X1 U409 ( .A(n338), .B(n337), .ZN(n340) );
  XOR2_X1 U410 ( .A(G50GAT), .B(G204GAT), .Z(n339) );
  XNOR2_X1 U411 ( .A(n340), .B(n339), .ZN(n342) );
  XOR2_X1 U412 ( .A(KEYINPUT24), .B(KEYINPUT93), .Z(n341) );
  NAND2_X1 U413 ( .A1(G228GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U414 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U415 ( .A(n371), .B(n347), .ZN(n470) );
  XOR2_X1 U416 ( .A(G176GAT), .B(G169GAT), .Z(n349) );
  XNOR2_X1 U417 ( .A(G120GAT), .B(G15GAT), .ZN(n348) );
  XNOR2_X1 U418 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U419 ( .A(KEYINPUT85), .B(KEYINPUT86), .Z(n351) );
  XNOR2_X1 U420 ( .A(G71GAT), .B(KEYINPUT66), .ZN(n350) );
  XNOR2_X1 U421 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U422 ( .A(n353), .B(n352), .Z(n358) );
  XOR2_X1 U423 ( .A(KEYINPUT87), .B(KEYINPUT20), .Z(n355) );
  NAND2_X1 U424 ( .A1(G227GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U425 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U426 ( .A(KEYINPUT88), .B(n356), .ZN(n357) );
  XNOR2_X1 U427 ( .A(n358), .B(n357), .ZN(n364) );
  XOR2_X1 U428 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n360) );
  XNOR2_X1 U429 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n359) );
  XNOR2_X1 U430 ( .A(n360), .B(n359), .ZN(n372) );
  XOR2_X1 U431 ( .A(n372), .B(G99GAT), .Z(n362) );
  XNOR2_X1 U432 ( .A(G134GAT), .B(G190GAT), .ZN(n361) );
  XNOR2_X1 U433 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U434 ( .A(n364), .B(n363), .Z(n367) );
  XNOR2_X1 U435 ( .A(n365), .B(G43GAT), .ZN(n366) );
  XOR2_X1 U436 ( .A(n367), .B(n366), .Z(n535) );
  INV_X1 U437 ( .A(n535), .ZN(n529) );
  XOR2_X1 U438 ( .A(G204GAT), .B(KEYINPUT72), .Z(n369) );
  XNOR2_X1 U439 ( .A(G92GAT), .B(G176GAT), .ZN(n368) );
  XNOR2_X1 U440 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U441 ( .A(G64GAT), .B(n370), .ZN(n430) );
  XOR2_X1 U442 ( .A(n430), .B(n371), .Z(n379) );
  XOR2_X1 U443 ( .A(G190GAT), .B(G36GAT), .Z(n402) );
  NAND2_X1 U444 ( .A1(G226GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U445 ( .A(n289), .B(n373), .ZN(n377) );
  XOR2_X1 U446 ( .A(G8GAT), .B(G169GAT), .Z(n444) );
  XNOR2_X1 U447 ( .A(KEYINPUT80), .B(n444), .ZN(n375) );
  XOR2_X1 U448 ( .A(n379), .B(n378), .Z(n504) );
  INV_X1 U449 ( .A(n504), .ZN(n526) );
  XOR2_X1 U450 ( .A(KEYINPUT99), .B(n380), .Z(n381) );
  NOR2_X1 U451 ( .A1(n470), .A2(n381), .ZN(n382) );
  XNOR2_X1 U452 ( .A(n382), .B(KEYINPUT25), .ZN(n386) );
  NAND2_X1 U453 ( .A1(n470), .A2(n529), .ZN(n383) );
  XNOR2_X1 U454 ( .A(KEYINPUT26), .B(n383), .ZN(n566) );
  INV_X1 U455 ( .A(n566), .ZN(n384) );
  XOR2_X1 U456 ( .A(KEYINPUT27), .B(n526), .Z(n390) );
  NAND2_X1 U457 ( .A1(n384), .A2(n390), .ZN(n385) );
  NAND2_X1 U458 ( .A1(n386), .A2(n385), .ZN(n388) );
  NAND2_X1 U459 ( .A1(n388), .A2(n387), .ZN(n389) );
  XOR2_X1 U460 ( .A(KEYINPUT100), .B(n389), .Z(n394) );
  XOR2_X1 U461 ( .A(KEYINPUT28), .B(n470), .Z(n534) );
  INV_X1 U462 ( .A(n534), .ZN(n507) );
  INV_X1 U463 ( .A(n514), .ZN(n501) );
  AND2_X1 U464 ( .A1(n390), .A2(n501), .ZN(n391) );
  XNOR2_X1 U465 ( .A(n391), .B(KEYINPUT98), .ZN(n532) );
  NAND2_X1 U466 ( .A1(n529), .A2(n532), .ZN(n392) );
  NOR2_X1 U467 ( .A1(n507), .A2(n392), .ZN(n393) );
  XNOR2_X1 U468 ( .A(KEYINPUT101), .B(n395), .ZN(n489) );
  NAND2_X1 U469 ( .A1(n563), .A2(n489), .ZN(n396) );
  XNOR2_X1 U470 ( .A(n396), .B(KEYINPUT105), .ZN(n414) );
  XOR2_X1 U471 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n398) );
  XNOR2_X1 U472 ( .A(KEYINPUT77), .B(KEYINPUT76), .ZN(n397) );
  XNOR2_X1 U473 ( .A(n398), .B(n397), .ZN(n413) );
  XNOR2_X1 U474 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n399) );
  XNOR2_X1 U475 ( .A(n288), .B(n399), .ZN(n441) );
  XOR2_X1 U476 ( .A(G106GAT), .B(n441), .Z(n401) );
  NAND2_X1 U477 ( .A1(G232GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U478 ( .A(n401), .B(n400), .ZN(n411) );
  XOR2_X1 U479 ( .A(KEYINPUT9), .B(G218GAT), .Z(n404) );
  XOR2_X1 U480 ( .A(G85GAT), .B(G99GAT), .Z(n417) );
  XNOR2_X1 U481 ( .A(n402), .B(n417), .ZN(n403) );
  XNOR2_X1 U482 ( .A(n404), .B(n403), .ZN(n409) );
  XOR2_X1 U483 ( .A(G92GAT), .B(KEYINPUT78), .Z(n406) );
  XNOR2_X1 U484 ( .A(G162GAT), .B(KEYINPUT79), .ZN(n405) );
  XNOR2_X1 U485 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U486 ( .A(n413), .B(n412), .ZN(n486) );
  XOR2_X1 U487 ( .A(KEYINPUT36), .B(n486), .Z(n579) );
  NAND2_X1 U488 ( .A1(n414), .A2(n579), .ZN(n415) );
  XNOR2_X1 U489 ( .A(KEYINPUT37), .B(n415), .ZN(n478) );
  AND2_X1 U490 ( .A1(G230GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U491 ( .A(n420), .B(G148GAT), .ZN(n427) );
  XOR2_X1 U492 ( .A(KEYINPUT74), .B(KEYINPUT32), .Z(n424) );
  XNOR2_X1 U493 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U494 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U495 ( .A(n425), .B(KEYINPUT73), .Z(n426) );
  XNOR2_X1 U496 ( .A(n427), .B(n426), .ZN(n432) );
  XOR2_X1 U497 ( .A(KEYINPUT31), .B(KEYINPUT69), .Z(n429) );
  XNOR2_X1 U498 ( .A(KEYINPUT75), .B(KEYINPUT33), .ZN(n428) );
  XNOR2_X1 U499 ( .A(n456), .B(KEYINPUT41), .ZN(n434) );
  INV_X1 U500 ( .A(KEYINPUT64), .ZN(n433) );
  XNOR2_X1 U501 ( .A(n434), .B(n433), .ZN(n549) );
  INV_X1 U502 ( .A(n549), .ZN(n474) );
  XOR2_X1 U503 ( .A(KEYINPUT67), .B(G197GAT), .Z(n436) );
  XNOR2_X1 U504 ( .A(G141GAT), .B(G113GAT), .ZN(n435) );
  XNOR2_X1 U505 ( .A(n436), .B(n435), .ZN(n449) );
  XOR2_X1 U506 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n438) );
  NAND2_X1 U507 ( .A1(G229GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U508 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U509 ( .A(n439), .B(KEYINPUT29), .Z(n443) );
  XNOR2_X1 U510 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U511 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U512 ( .A(n445), .B(n444), .Z(n447) );
  XNOR2_X1 U513 ( .A(G29GAT), .B(G36GAT), .ZN(n446) );
  XNOR2_X1 U514 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U515 ( .A(n449), .B(n448), .ZN(n567) );
  NOR2_X1 U516 ( .A1(n474), .A2(n567), .ZN(n513) );
  NAND2_X1 U517 ( .A1(n478), .A2(n513), .ZN(n528) );
  NOR2_X1 U518 ( .A1(n514), .A2(n528), .ZN(n452) );
  INV_X1 U519 ( .A(KEYINPUT114), .ZN(n450) );
  NOR2_X1 U520 ( .A1(n534), .A2(n528), .ZN(n455) );
  XNOR2_X1 U521 ( .A(n455), .B(n454), .ZN(G1339GAT) );
  XOR2_X1 U522 ( .A(n504), .B(KEYINPUT121), .Z(n465) );
  NAND2_X1 U523 ( .A1(n575), .A2(n579), .ZN(n457) );
  XOR2_X1 U524 ( .A(KEYINPUT45), .B(n457), .Z(n458) );
  INV_X1 U525 ( .A(n567), .ZN(n560) );
  NAND2_X1 U526 ( .A1(n458), .A2(n560), .ZN(n459) );
  AND2_X1 U527 ( .A1(n549), .A2(n567), .ZN(n460) );
  XNOR2_X1 U528 ( .A(n460), .B(KEYINPUT46), .ZN(n462) );
  INV_X1 U529 ( .A(n486), .ZN(n557) );
  OR2_X1 U530 ( .A1(n557), .A2(n575), .ZN(n461) );
  NAND2_X1 U531 ( .A1(n465), .A2(n533), .ZN(n466) );
  XNOR2_X1 U532 ( .A(n466), .B(KEYINPUT122), .ZN(n467) );
  XNOR2_X1 U533 ( .A(n467), .B(KEYINPUT54), .ZN(n468) );
  NOR2_X1 U534 ( .A1(n468), .A2(n501), .ZN(n469) );
  XNOR2_X1 U535 ( .A(n469), .B(KEYINPUT65), .ZN(n565) );
  XNOR2_X1 U536 ( .A(n472), .B(n471), .ZN(n473) );
  NAND2_X1 U537 ( .A1(n473), .A2(n535), .ZN(n562) );
  NOR2_X1 U538 ( .A1(n562), .A2(n474), .ZN(n477) );
  XNOR2_X1 U539 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n475) );
  XNOR2_X1 U540 ( .A(n475), .B(G176GAT), .ZN(n476) );
  XNOR2_X1 U541 ( .A(n477), .B(n476), .ZN(G1349GAT) );
  XOR2_X1 U542 ( .A(KEYINPUT38), .B(KEYINPUT106), .Z(n480) );
  NOR2_X1 U543 ( .A1(n560), .A2(n456), .ZN(n490) );
  NAND2_X1 U544 ( .A1(n490), .A2(n478), .ZN(n479) );
  NAND2_X1 U545 ( .A1(n535), .A2(n508), .ZN(n482) );
  XNOR2_X1 U546 ( .A(n482), .B(n481), .ZN(G1330GAT) );
  NOR2_X1 U547 ( .A1(n486), .A2(n562), .ZN(n485) );
  XNOR2_X1 U548 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n483) );
  NAND2_X1 U549 ( .A1(n575), .A2(n486), .ZN(n487) );
  XOR2_X1 U550 ( .A(KEYINPUT16), .B(n487), .Z(n488) );
  AND2_X1 U551 ( .A1(n489), .A2(n488), .ZN(n512) );
  NAND2_X1 U552 ( .A1(n490), .A2(n512), .ZN(n499) );
  NOR2_X1 U553 ( .A1(n514), .A2(n499), .ZN(n492) );
  XNOR2_X1 U554 ( .A(KEYINPUT102), .B(KEYINPUT34), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U556 ( .A(G1GAT), .B(n493), .Z(G1324GAT) );
  NOR2_X1 U557 ( .A1(n526), .A2(n499), .ZN(n495) );
  XNOR2_X1 U558 ( .A(G8GAT), .B(KEYINPUT103), .ZN(n494) );
  XNOR2_X1 U559 ( .A(n495), .B(n494), .ZN(G1325GAT) );
  NOR2_X1 U560 ( .A1(n529), .A2(n499), .ZN(n497) );
  XNOR2_X1 U561 ( .A(KEYINPUT35), .B(KEYINPUT104), .ZN(n496) );
  XNOR2_X1 U562 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U563 ( .A(G15GAT), .B(n498), .ZN(G1326GAT) );
  NOR2_X1 U564 ( .A1(n534), .A2(n499), .ZN(n500) );
  XOR2_X1 U565 ( .A(G22GAT), .B(n500), .Z(G1327GAT) );
  XOR2_X1 U566 ( .A(G29GAT), .B(KEYINPUT39), .Z(n503) );
  NAND2_X1 U567 ( .A1(n508), .A2(n501), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  XOR2_X1 U569 ( .A(G36GAT), .B(KEYINPUT107), .Z(n506) );
  NAND2_X1 U570 ( .A1(n508), .A2(n504), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(G1329GAT) );
  NAND2_X1 U572 ( .A1(n508), .A2(n507), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n509), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n511) );
  XNOR2_X1 U575 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(n516) );
  NAND2_X1 U577 ( .A1(n513), .A2(n512), .ZN(n522) );
  NOR2_X1 U578 ( .A1(n514), .A2(n522), .ZN(n515) );
  XOR2_X1 U579 ( .A(n516), .B(n515), .Z(n517) );
  XNOR2_X1 U580 ( .A(KEYINPUT108), .B(n517), .ZN(G1332GAT) );
  NOR2_X1 U581 ( .A1(n526), .A2(n522), .ZN(n519) );
  XNOR2_X1 U582 ( .A(G64GAT), .B(KEYINPUT111), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(G1333GAT) );
  NOR2_X1 U584 ( .A1(n529), .A2(n522), .ZN(n520) );
  XOR2_X1 U585 ( .A(KEYINPUT112), .B(n520), .Z(n521) );
  XNOR2_X1 U586 ( .A(G71GAT), .B(n521), .ZN(G1334GAT) );
  NOR2_X1 U587 ( .A1(n534), .A2(n522), .ZN(n524) );
  XNOR2_X1 U588 ( .A(KEYINPUT113), .B(KEYINPUT43), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U590 ( .A(G78GAT), .B(n525), .Z(G1335GAT) );
  NOR2_X1 U591 ( .A1(n526), .A2(n528), .ZN(n527) );
  XOR2_X1 U592 ( .A(G92GAT), .B(n527), .Z(G1337GAT) );
  NOR2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n531) );
  XNOR2_X1 U594 ( .A(G99GAT), .B(KEYINPUT115), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(G1338GAT) );
  NAND2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n547) );
  NAND2_X1 U597 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U598 ( .A1(n547), .A2(n536), .ZN(n544) );
  NAND2_X1 U599 ( .A1(n544), .A2(n567), .ZN(n537) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U602 ( .A1(n544), .A2(n549), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U604 ( .A(G120GAT), .B(n540), .ZN(G1341GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n542) );
  NAND2_X1 U606 ( .A1(n544), .A2(n575), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U609 ( .A(G134GAT), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U610 ( .A1(n544), .A2(n557), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  NOR2_X1 U612 ( .A1(n566), .A2(n547), .ZN(n558) );
  NAND2_X1 U613 ( .A1(n558), .A2(n567), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(n548), .ZN(G1344GAT) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n553) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n551) );
  NAND2_X1 U617 ( .A1(n558), .A2(n549), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n555) );
  NAND2_X1 U621 ( .A1(n558), .A2(n575), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(G155GAT), .B(n556), .ZN(G1346GAT) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U626 ( .A1(n560), .A2(n562), .ZN(n561) );
  XOR2_X1 U627 ( .A(G169GAT), .B(n561), .Z(G1348GAT) );
  NOR2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U629 ( .A(G183GAT), .B(n564), .Z(G1350GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n569) );
  NOR2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n578) );
  NAND2_X1 U632 ( .A1(n578), .A2(n567), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n570), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n572) );
  NAND2_X1 U636 ( .A1(n578), .A2(n456), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n574) );
  XOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT124), .Z(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  NAND2_X1 U640 ( .A1(n578), .A2(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(KEYINPUT126), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G211GAT), .B(n577), .ZN(G1354GAT) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(n580), .B(KEYINPUT62), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

