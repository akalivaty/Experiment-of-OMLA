

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U550 ( .A1(G651), .A2(n683), .ZN(n697) );
  AND2_X1 U551 ( .A1(G2105), .A2(G2104), .ZN(n601) );
  XNOR2_X1 U552 ( .A(n585), .B(n584), .ZN(n661) );
  NOR2_X2 U553 ( .A1(n732), .A2(n731), .ZN(n734) );
  XNOR2_X2 U554 ( .A(G2104), .B(KEYINPUT64), .ZN(n594) );
  AND2_X2 U555 ( .A1(G101), .A2(n661), .ZN(n587) );
  INV_X1 U556 ( .A(KEYINPUT65), .ZN(n584) );
  INV_X1 U557 ( .A(G40), .ZN(n731) );
  NOR2_X2 U558 ( .A1(G2105), .A2(G2104), .ZN(n589) );
  AND2_X1 U559 ( .A1(n522), .A2(n520), .ZN(n519) );
  AND2_X1 U560 ( .A1(n592), .A2(n524), .ZN(n521) );
  AND2_X2 U561 ( .A1(n595), .A2(G2105), .ZN(n925) );
  XNOR2_X1 U562 ( .A(n591), .B(KEYINPUT66), .ZN(n592) );
  AND2_X1 U563 ( .A1(n594), .A2(n583), .ZN(n585) );
  NAND2_X1 U564 ( .A1(n601), .A2(G113), .ZN(n591) );
  NOR2_X1 U565 ( .A1(n532), .A2(n528), .ZN(n527) );
  NOR2_X1 U566 ( .A1(n784), .A2(n533), .ZN(n532) );
  OR2_X4 U567 ( .A1(n819), .A2(n818), .ZN(n740) );
  XNOR2_X2 U568 ( .A(n590), .B(n589), .ZN(n598) );
  AND2_X1 U569 ( .A1(n556), .A2(G8), .ZN(n555) );
  NAND2_X1 U570 ( .A1(n779), .A2(KEYINPUT97), .ZN(n533) );
  OR2_X1 U571 ( .A1(G286), .A2(n533), .ZN(n531) );
  NOR2_X1 U572 ( .A1(n544), .A2(n545), .ZN(n735) );
  NAND2_X1 U573 ( .A1(n550), .A2(n546), .ZN(n545) );
  NAND2_X1 U574 ( .A1(n547), .A2(n554), .ZN(n544) );
  INV_X1 U575 ( .A(KEYINPUT96), .ZN(n774) );
  INV_X1 U576 ( .A(G1384), .ZN(n729) );
  NOR2_X1 U577 ( .A1(n536), .A2(KEYINPUT101), .ZN(n535) );
  NOR2_X1 U578 ( .A1(n850), .A2(n852), .ZN(n541) );
  BUF_X1 U579 ( .A(n601), .Z(n926) );
  NAND2_X1 U580 ( .A1(n523), .A2(KEYINPUT68), .ZN(n522) );
  NAND2_X1 U581 ( .A1(n518), .A2(KEYINPUT68), .ZN(n517) );
  NOR2_X1 U582 ( .A1(n740), .A2(n1039), .ZN(n751) );
  INV_X1 U583 ( .A(G1966), .ZN(n546) );
  NAND2_X1 U584 ( .A1(n531), .A2(n529), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n530), .A2(n780), .ZN(n529) );
  AND2_X1 U586 ( .A1(G286), .A2(n780), .ZN(n526) );
  OR2_X1 U587 ( .A1(n548), .A2(n819), .ZN(n547) );
  AND2_X1 U588 ( .A1(n553), .A2(n551), .ZN(n550) );
  NAND2_X1 U589 ( .A1(n552), .A2(KEYINPUT92), .ZN(n551) );
  AND2_X1 U590 ( .A1(n542), .A2(n540), .ZN(n539) );
  NOR2_X1 U591 ( .A1(n541), .A2(n515), .ZN(n540) );
  NAND2_X1 U592 ( .A1(n538), .A2(KEYINPUT101), .ZN(n537) );
  OR2_X1 U593 ( .A1(n605), .A2(n604), .ZN(n730) );
  AND2_X1 U594 ( .A1(n596), .A2(n517), .ZN(n516) );
  XOR2_X1 U595 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U596 ( .A1(n550), .A2(n554), .ZN(n514) );
  INV_X1 U597 ( .A(KEYINPUT97), .ZN(n780) );
  NAND2_X1 U598 ( .A1(n730), .A2(n729), .ZN(n818) );
  INV_X1 U599 ( .A(n818), .ZN(n549) );
  INV_X1 U600 ( .A(G8), .ZN(n552) );
  NAND2_X1 U601 ( .A1(n519), .A2(n516), .ZN(n732) );
  AND2_X1 U602 ( .A1(n1014), .A2(n864), .ZN(n515) );
  INV_X1 U603 ( .A(KEYINPUT101), .ZN(n852) );
  INV_X1 U604 ( .A(n592), .ZN(n518) );
  NAND2_X1 U605 ( .A1(n593), .A2(n521), .ZN(n520) );
  INV_X1 U606 ( .A(n593), .ZN(n523) );
  INV_X1 U607 ( .A(KEYINPUT68), .ZN(n524) );
  NAND2_X1 U608 ( .A1(n527), .A2(n525), .ZN(n534) );
  NAND2_X1 U609 ( .A1(n784), .A2(n526), .ZN(n525) );
  INV_X1 U610 ( .A(n779), .ZN(n530) );
  NAND2_X1 U611 ( .A1(n534), .A2(G8), .ZN(n782) );
  NAND2_X1 U612 ( .A1(n851), .A2(n535), .ZN(n542) );
  INV_X1 U613 ( .A(n850), .ZN(n536) );
  NAND2_X1 U614 ( .A1(n539), .A2(n537), .ZN(n543) );
  INV_X1 U615 ( .A(n851), .ZN(n538) );
  NAND2_X1 U616 ( .A1(n543), .A2(n866), .ZN(n867) );
  NAND2_X1 U617 ( .A1(n547), .A2(n514), .ZN(n799) );
  NAND2_X1 U618 ( .A1(n549), .A2(KEYINPUT92), .ZN(n548) );
  NAND2_X1 U619 ( .A1(n818), .A2(n555), .ZN(n553) );
  NAND2_X1 U620 ( .A1(n819), .A2(n555), .ZN(n554) );
  INV_X1 U621 ( .A(KEYINPUT92), .ZN(n556) );
  INV_X2 U622 ( .A(n740), .ZN(n755) );
  NOR2_X1 U623 ( .A1(n785), .A2(n552), .ZN(n557) );
  OR2_X1 U624 ( .A1(n846), .A2(n845), .ZN(n558) );
  INV_X1 U625 ( .A(KEYINPUT26), .ZN(n750) );
  XOR2_X1 U626 ( .A(KEYINPUT30), .B(KEYINPUT95), .Z(n737) );
  BUF_X1 U627 ( .A(n598), .Z(n921) );
  INV_X1 U628 ( .A(G651), .ZN(n565) );
  NOR2_X1 U629 ( .A1(G543), .A2(n565), .ZN(n560) );
  XNOR2_X1 U630 ( .A(KEYINPUT1), .B(KEYINPUT69), .ZN(n559) );
  XNOR2_X2 U631 ( .A(n560), .B(n559), .ZN(n700) );
  NAND2_X1 U632 ( .A1(G63), .A2(n700), .ZN(n562) );
  XOR2_X1 U633 ( .A(KEYINPUT0), .B(G543), .Z(n683) );
  NAND2_X1 U634 ( .A1(G51), .A2(n697), .ZN(n561) );
  NAND2_X1 U635 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U636 ( .A(KEYINPUT6), .B(n563), .ZN(n571) );
  NOR2_X1 U637 ( .A1(G651), .A2(G543), .ZN(n701) );
  NAND2_X1 U638 ( .A1(n701), .A2(G89), .ZN(n564) );
  XNOR2_X1 U639 ( .A(n564), .B(KEYINPUT4), .ZN(n567) );
  NOR2_X1 U640 ( .A1(n683), .A2(n565), .ZN(n696) );
  NAND2_X1 U641 ( .A1(G76), .A2(n696), .ZN(n566) );
  NAND2_X1 U642 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U643 ( .A(KEYINPUT5), .B(n568), .ZN(n569) );
  XNOR2_X1 U644 ( .A(KEYINPUT75), .B(n569), .ZN(n570) );
  NOR2_X1 U645 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U646 ( .A(KEYINPUT7), .B(n572), .Z(G168) );
  XOR2_X1 U647 ( .A(G2438), .B(G2454), .Z(n574) );
  XNOR2_X1 U648 ( .A(G2435), .B(G2430), .ZN(n573) );
  XNOR2_X1 U649 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U650 ( .A(n575), .B(G2427), .Z(n577) );
  XNOR2_X1 U651 ( .A(G1341), .B(G1348), .ZN(n576) );
  XNOR2_X1 U652 ( .A(n577), .B(n576), .ZN(n581) );
  XOR2_X1 U653 ( .A(G2443), .B(G2446), .Z(n579) );
  XNOR2_X1 U654 ( .A(KEYINPUT104), .B(G2451), .ZN(n578) );
  XNOR2_X1 U655 ( .A(n579), .B(n578), .ZN(n580) );
  XOR2_X1 U656 ( .A(n581), .B(n580), .Z(n582) );
  AND2_X1 U657 ( .A1(G14), .A2(n582), .ZN(G401) );
  INV_X1 U658 ( .A(G2105), .ZN(n583) );
  INV_X1 U659 ( .A(KEYINPUT23), .ZN(n586) );
  XNOR2_X1 U660 ( .A(n587), .B(n586), .ZN(n588) );
  INV_X1 U661 ( .A(n588), .ZN(n733) );
  XNOR2_X2 U662 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n590) );
  NAND2_X1 U663 ( .A1(n598), .A2(G137), .ZN(n593) );
  INV_X1 U664 ( .A(n594), .ZN(n595) );
  NAND2_X1 U665 ( .A1(n925), .A2(G125), .ZN(n596) );
  INV_X1 U666 ( .A(n732), .ZN(n597) );
  AND2_X1 U667 ( .A1(n733), .A2(n597), .ZN(G160) );
  AND2_X1 U668 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U669 ( .A(G69), .ZN(G235) );
  INV_X1 U670 ( .A(G132), .ZN(G219) );
  INV_X1 U671 ( .A(G82), .ZN(G220) );
  NAND2_X1 U672 ( .A1(n598), .A2(G138), .ZN(n600) );
  NAND2_X1 U673 ( .A1(n661), .A2(G102), .ZN(n599) );
  NAND2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n605) );
  NAND2_X1 U675 ( .A1(G126), .A2(n925), .ZN(n603) );
  NAND2_X1 U676 ( .A1(G114), .A2(n926), .ZN(n602) );
  NAND2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n604) );
  INV_X1 U678 ( .A(n730), .ZN(G164) );
  NAND2_X1 U679 ( .A1(G64), .A2(n700), .ZN(n608) );
  NAND2_X1 U680 ( .A1(G52), .A2(n697), .ZN(n607) );
  NAND2_X1 U681 ( .A1(n608), .A2(n607), .ZN(n613) );
  NAND2_X1 U682 ( .A1(G90), .A2(n701), .ZN(n610) );
  NAND2_X1 U683 ( .A1(G77), .A2(n696), .ZN(n609) );
  NAND2_X1 U684 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U685 ( .A(KEYINPUT9), .B(n611), .Z(n612) );
  NOR2_X1 U686 ( .A1(n613), .A2(n612), .ZN(G171) );
  NAND2_X1 U687 ( .A1(G7), .A2(G661), .ZN(n614) );
  XNOR2_X1 U688 ( .A(n614), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U689 ( .A(G223), .ZN(n868) );
  NAND2_X1 U690 ( .A1(n868), .A2(G567), .ZN(n615) );
  XNOR2_X1 U691 ( .A(n615), .B(KEYINPUT71), .ZN(n616) );
  XNOR2_X1 U692 ( .A(KEYINPUT11), .B(n616), .ZN(G234) );
  XOR2_X1 U693 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n618) );
  NAND2_X1 U694 ( .A1(G56), .A2(n700), .ZN(n617) );
  XNOR2_X1 U695 ( .A(n618), .B(n617), .ZN(n625) );
  XNOR2_X1 U696 ( .A(KEYINPUT13), .B(KEYINPUT73), .ZN(n623) );
  NAND2_X1 U697 ( .A1(n701), .A2(G81), .ZN(n619) );
  XNOR2_X1 U698 ( .A(n619), .B(KEYINPUT12), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G68), .A2(n696), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U701 ( .A(n623), .B(n622), .ZN(n624) );
  NOR2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n697), .A2(G43), .ZN(n626) );
  NAND2_X1 U704 ( .A1(n627), .A2(n626), .ZN(n1022) );
  INV_X1 U705 ( .A(G860), .ZN(n649) );
  OR2_X1 U706 ( .A1(n1022), .A2(n649), .ZN(G153) );
  INV_X1 U707 ( .A(G171), .ZN(G301) );
  NAND2_X1 U708 ( .A1(G868), .A2(G301), .ZN(n637) );
  NAND2_X1 U709 ( .A1(G79), .A2(n696), .ZN(n629) );
  NAND2_X1 U710 ( .A1(G54), .A2(n697), .ZN(n628) );
  NAND2_X1 U711 ( .A1(n629), .A2(n628), .ZN(n634) );
  NAND2_X1 U712 ( .A1(G66), .A2(n700), .ZN(n631) );
  NAND2_X1 U713 ( .A1(G92), .A2(n701), .ZN(n630) );
  NAND2_X1 U714 ( .A1(n631), .A2(n630), .ZN(n632) );
  XNOR2_X1 U715 ( .A(KEYINPUT74), .B(n632), .ZN(n633) );
  NOR2_X1 U716 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X2 U717 ( .A(n635), .B(KEYINPUT15), .ZN(n1017) );
  INV_X1 U718 ( .A(G868), .ZN(n653) );
  NAND2_X1 U719 ( .A1(n1017), .A2(n653), .ZN(n636) );
  NAND2_X1 U720 ( .A1(n637), .A2(n636), .ZN(G284) );
  NAND2_X1 U721 ( .A1(G65), .A2(n700), .ZN(n639) );
  NAND2_X1 U722 ( .A1(G78), .A2(n696), .ZN(n638) );
  NAND2_X1 U723 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U724 ( .A1(n701), .A2(G91), .ZN(n640) );
  XOR2_X1 U725 ( .A(KEYINPUT70), .B(n640), .Z(n641) );
  NOR2_X1 U726 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U727 ( .A1(n697), .A2(G53), .ZN(n643) );
  NAND2_X1 U728 ( .A1(n644), .A2(n643), .ZN(G299) );
  NOR2_X1 U729 ( .A1(G286), .A2(n653), .ZN(n645) );
  XNOR2_X1 U730 ( .A(n645), .B(KEYINPUT76), .ZN(n647) );
  NOR2_X1 U731 ( .A1(G299), .A2(G868), .ZN(n646) );
  NOR2_X1 U732 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U733 ( .A(KEYINPUT77), .B(n648), .Z(G297) );
  NAND2_X1 U734 ( .A1(n649), .A2(G559), .ZN(n650) );
  INV_X1 U735 ( .A(n1017), .ZN(n711) );
  NAND2_X1 U736 ( .A1(n650), .A2(n711), .ZN(n651) );
  XNOR2_X1 U737 ( .A(n651), .B(KEYINPUT16), .ZN(n652) );
  XNOR2_X1 U738 ( .A(KEYINPUT78), .B(n652), .ZN(G148) );
  NOR2_X1 U739 ( .A1(n1017), .A2(n653), .ZN(n654) );
  XNOR2_X1 U740 ( .A(n654), .B(KEYINPUT79), .ZN(n655) );
  NOR2_X1 U741 ( .A1(G559), .A2(n655), .ZN(n657) );
  NOR2_X1 U742 ( .A1(G868), .A2(n1022), .ZN(n656) );
  NOR2_X1 U743 ( .A1(n657), .A2(n656), .ZN(G282) );
  NAND2_X1 U744 ( .A1(n925), .A2(G123), .ZN(n658) );
  XNOR2_X1 U745 ( .A(n658), .B(KEYINPUT18), .ZN(n660) );
  NAND2_X1 U746 ( .A1(G111), .A2(n926), .ZN(n659) );
  NAND2_X1 U747 ( .A1(n660), .A2(n659), .ZN(n665) );
  NAND2_X1 U748 ( .A1(G135), .A2(n921), .ZN(n663) );
  BUF_X1 U749 ( .A(n661), .Z(n922) );
  NAND2_X1 U750 ( .A1(G99), .A2(n922), .ZN(n662) );
  NAND2_X1 U751 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U752 ( .A1(n665), .A2(n664), .ZN(n968) );
  XOR2_X1 U753 ( .A(n968), .B(G2096), .Z(n666) );
  NOR2_X1 U754 ( .A1(G2100), .A2(n666), .ZN(n667) );
  XOR2_X1 U755 ( .A(KEYINPUT80), .B(n667), .Z(G156) );
  NAND2_X1 U756 ( .A1(G62), .A2(n700), .ZN(n669) );
  NAND2_X1 U757 ( .A1(G88), .A2(n701), .ZN(n668) );
  NAND2_X1 U758 ( .A1(n669), .A2(n668), .ZN(n672) );
  NAND2_X1 U759 ( .A1(n696), .A2(G75), .ZN(n670) );
  XOR2_X1 U760 ( .A(KEYINPUT84), .B(n670), .Z(n671) );
  NOR2_X1 U761 ( .A1(n672), .A2(n671), .ZN(n674) );
  NAND2_X1 U762 ( .A1(n697), .A2(G50), .ZN(n673) );
  NAND2_X1 U763 ( .A1(n674), .A2(n673), .ZN(G303) );
  INV_X1 U764 ( .A(G303), .ZN(G166) );
  NAND2_X1 U765 ( .A1(G61), .A2(n700), .ZN(n676) );
  NAND2_X1 U766 ( .A1(G86), .A2(n701), .ZN(n675) );
  NAND2_X1 U767 ( .A1(n676), .A2(n675), .ZN(n680) );
  NAND2_X1 U768 ( .A1(G73), .A2(n696), .ZN(n677) );
  XNOR2_X1 U769 ( .A(n677), .B(KEYINPUT83), .ZN(n678) );
  XNOR2_X1 U770 ( .A(n678), .B(KEYINPUT2), .ZN(n679) );
  NOR2_X1 U771 ( .A1(n680), .A2(n679), .ZN(n682) );
  NAND2_X1 U772 ( .A1(n697), .A2(G48), .ZN(n681) );
  NAND2_X1 U773 ( .A1(n682), .A2(n681), .ZN(G305) );
  NAND2_X1 U774 ( .A1(G87), .A2(n683), .ZN(n684) );
  XNOR2_X1 U775 ( .A(n684), .B(KEYINPUT82), .ZN(n689) );
  NAND2_X1 U776 ( .A1(G49), .A2(n697), .ZN(n686) );
  NAND2_X1 U777 ( .A1(G74), .A2(G651), .ZN(n685) );
  NAND2_X1 U778 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U779 ( .A1(n700), .A2(n687), .ZN(n688) );
  NAND2_X1 U780 ( .A1(n689), .A2(n688), .ZN(G288) );
  AND2_X1 U781 ( .A1(n700), .A2(G60), .ZN(n693) );
  NAND2_X1 U782 ( .A1(G85), .A2(n701), .ZN(n691) );
  NAND2_X1 U783 ( .A1(G72), .A2(n696), .ZN(n690) );
  NAND2_X1 U784 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U785 ( .A1(n693), .A2(n692), .ZN(n695) );
  NAND2_X1 U786 ( .A1(n697), .A2(G47), .ZN(n694) );
  NAND2_X1 U787 ( .A1(n695), .A2(n694), .ZN(G290) );
  NAND2_X1 U788 ( .A1(G80), .A2(n696), .ZN(n699) );
  NAND2_X1 U789 ( .A1(G55), .A2(n697), .ZN(n698) );
  NAND2_X1 U790 ( .A1(n699), .A2(n698), .ZN(n705) );
  NAND2_X1 U791 ( .A1(G67), .A2(n700), .ZN(n703) );
  NAND2_X1 U792 ( .A1(G93), .A2(n701), .ZN(n702) );
  NAND2_X1 U793 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U794 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U795 ( .A(n706), .B(KEYINPUT81), .ZN(n945) );
  XNOR2_X1 U796 ( .A(KEYINPUT19), .B(G305), .ZN(n707) );
  XNOR2_X1 U797 ( .A(n707), .B(G288), .ZN(n708) );
  XNOR2_X1 U798 ( .A(G166), .B(n708), .ZN(n710) );
  INV_X1 U799 ( .A(G299), .ZN(n1012) );
  XNOR2_X1 U800 ( .A(G290), .B(n1012), .ZN(n709) );
  XNOR2_X1 U801 ( .A(n710), .B(n709), .ZN(n944) );
  NAND2_X1 U802 ( .A1(G559), .A2(n711), .ZN(n712) );
  XNOR2_X1 U803 ( .A(n712), .B(n1022), .ZN(n874) );
  XNOR2_X1 U804 ( .A(n944), .B(n874), .ZN(n713) );
  NAND2_X1 U805 ( .A1(n713), .A2(G868), .ZN(n714) );
  XNOR2_X1 U806 ( .A(n945), .B(n714), .ZN(G295) );
  NAND2_X1 U807 ( .A1(G2078), .A2(G2084), .ZN(n715) );
  XNOR2_X1 U808 ( .A(n715), .B(KEYINPUT85), .ZN(n716) );
  XNOR2_X1 U809 ( .A(KEYINPUT20), .B(n716), .ZN(n717) );
  NAND2_X1 U810 ( .A1(n717), .A2(G2090), .ZN(n718) );
  XNOR2_X1 U811 ( .A(n718), .B(KEYINPUT86), .ZN(n719) );
  XNOR2_X1 U812 ( .A(KEYINPUT21), .B(n719), .ZN(n720) );
  NAND2_X1 U813 ( .A1(n720), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U814 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U815 ( .A1(G220), .A2(G219), .ZN(n721) );
  XOR2_X1 U816 ( .A(KEYINPUT22), .B(n721), .Z(n722) );
  NOR2_X1 U817 ( .A1(G218), .A2(n722), .ZN(n723) );
  NAND2_X1 U818 ( .A1(G96), .A2(n723), .ZN(n872) );
  NAND2_X1 U819 ( .A1(G2106), .A2(n872), .ZN(n727) );
  NAND2_X1 U820 ( .A1(G120), .A2(G108), .ZN(n724) );
  NOR2_X1 U821 ( .A1(G235), .A2(n724), .ZN(n725) );
  NAND2_X1 U822 ( .A1(G57), .A2(n725), .ZN(n873) );
  NAND2_X1 U823 ( .A1(G567), .A2(n873), .ZN(n726) );
  NAND2_X1 U824 ( .A1(n727), .A2(n726), .ZN(n876) );
  NAND2_X1 U825 ( .A1(G483), .A2(G661), .ZN(n728) );
  NOR2_X1 U826 ( .A1(n876), .A2(n728), .ZN(n871) );
  NAND2_X1 U827 ( .A1(n871), .A2(G36), .ZN(G176) );
  NAND2_X1 U828 ( .A1(n734), .A2(n733), .ZN(n819) );
  XNOR2_X1 U829 ( .A(n735), .B(KEYINPUT94), .ZN(n783) );
  INV_X1 U830 ( .A(n783), .ZN(n736) );
  NOR2_X1 U831 ( .A1(G2084), .A2(n740), .ZN(n785) );
  NAND2_X1 U832 ( .A1(n736), .A2(n557), .ZN(n738) );
  XNOR2_X1 U833 ( .A(n738), .B(n737), .ZN(n739) );
  NOR2_X1 U834 ( .A1(n739), .A2(G168), .ZN(n744) );
  XOR2_X1 U835 ( .A(G2078), .B(KEYINPUT25), .Z(n1044) );
  NOR2_X1 U836 ( .A1(n1044), .A2(n740), .ZN(n742) );
  NOR2_X1 U837 ( .A1(n755), .A2(G1961), .ZN(n741) );
  NOR2_X1 U838 ( .A1(n742), .A2(n741), .ZN(n769) );
  AND2_X1 U839 ( .A1(G301), .A2(n769), .ZN(n743) );
  NOR2_X1 U840 ( .A1(n744), .A2(n743), .ZN(n745) );
  XNOR2_X1 U841 ( .A(n745), .B(KEYINPUT31), .ZN(n773) );
  NAND2_X1 U842 ( .A1(n755), .A2(G2072), .ZN(n746) );
  XNOR2_X1 U843 ( .A(n746), .B(KEYINPUT27), .ZN(n748) );
  INV_X1 U844 ( .A(G1956), .ZN(n983) );
  NOR2_X1 U845 ( .A1(n983), .A2(n755), .ZN(n747) );
  NOR2_X1 U846 ( .A1(n748), .A2(n747), .ZN(n763) );
  NOR2_X1 U847 ( .A1(n1012), .A2(n763), .ZN(n749) );
  XOR2_X1 U848 ( .A(n749), .B(KEYINPUT28), .Z(n767) );
  INV_X1 U849 ( .A(G1996), .ZN(n1039) );
  XNOR2_X1 U850 ( .A(n751), .B(n750), .ZN(n753) );
  NAND2_X1 U851 ( .A1(n740), .A2(G1341), .ZN(n752) );
  NAND2_X1 U852 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U853 ( .A1(n1022), .A2(n754), .ZN(n759) );
  NAND2_X1 U854 ( .A1(G1348), .A2(n740), .ZN(n757) );
  NAND2_X1 U855 ( .A1(G2067), .A2(n755), .ZN(n756) );
  NAND2_X1 U856 ( .A1(n757), .A2(n756), .ZN(n760) );
  NOR2_X1 U857 ( .A1(n1017), .A2(n760), .ZN(n758) );
  OR2_X1 U858 ( .A1(n759), .A2(n758), .ZN(n762) );
  NAND2_X1 U859 ( .A1(n1017), .A2(n760), .ZN(n761) );
  NAND2_X1 U860 ( .A1(n762), .A2(n761), .ZN(n765) );
  NAND2_X1 U861 ( .A1(n1012), .A2(n763), .ZN(n764) );
  NAND2_X1 U862 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U863 ( .A1(n767), .A2(n766), .ZN(n768) );
  XNOR2_X1 U864 ( .A(n768), .B(KEYINPUT29), .ZN(n771) );
  NOR2_X1 U865 ( .A1(G301), .A2(n769), .ZN(n770) );
  NOR2_X1 U866 ( .A1(n771), .A2(n770), .ZN(n772) );
  NOR2_X2 U867 ( .A1(n773), .A2(n772), .ZN(n775) );
  XNOR2_X2 U868 ( .A(n775), .B(n774), .ZN(n784) );
  NOR2_X1 U869 ( .A1(n799), .A2(G1971), .ZN(n777) );
  NOR2_X1 U870 ( .A1(G2090), .A2(n740), .ZN(n776) );
  NOR2_X1 U871 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U872 ( .A1(n778), .A2(G303), .ZN(n779) );
  INV_X1 U873 ( .A(KEYINPUT32), .ZN(n781) );
  XNOR2_X1 U874 ( .A(n782), .B(n781), .ZN(n840) );
  NAND2_X1 U875 ( .A1(G8), .A2(n785), .ZN(n786) );
  NAND2_X1 U876 ( .A1(n784), .A2(n786), .ZN(n787) );
  NOR2_X1 U877 ( .A1(n783), .A2(n787), .ZN(n841) );
  NAND2_X1 U878 ( .A1(G1976), .A2(G288), .ZN(n1025) );
  INV_X1 U879 ( .A(n1025), .ZN(n790) );
  OR2_X1 U880 ( .A1(n841), .A2(n790), .ZN(n788) );
  NOR2_X1 U881 ( .A1(n840), .A2(n788), .ZN(n792) );
  NOR2_X1 U882 ( .A1(G1976), .A2(G288), .ZN(n798) );
  NOR2_X1 U883 ( .A1(G1971), .A2(G303), .ZN(n789) );
  NOR2_X1 U884 ( .A1(n798), .A2(n789), .ZN(n1028) );
  NOR2_X1 U885 ( .A1(n790), .A2(n1028), .ZN(n791) );
  NOR2_X2 U886 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U887 ( .A(n793), .B(KEYINPUT98), .ZN(n794) );
  NOR2_X1 U888 ( .A1(n799), .A2(n794), .ZN(n795) );
  NOR2_X1 U889 ( .A1(n795), .A2(KEYINPUT33), .ZN(n796) );
  XNOR2_X1 U890 ( .A(n796), .B(KEYINPUT99), .ZN(n836) );
  XNOR2_X1 U891 ( .A(G1981), .B(KEYINPUT100), .ZN(n797) );
  XNOR2_X1 U892 ( .A(n797), .B(G305), .ZN(n1010) );
  AND2_X1 U893 ( .A1(n798), .A2(KEYINPUT33), .ZN(n800) );
  INV_X1 U894 ( .A(n799), .ZN(n845) );
  NAND2_X1 U895 ( .A1(n800), .A2(n845), .ZN(n833) );
  NAND2_X1 U896 ( .A1(G131), .A2(n921), .ZN(n802) );
  NAND2_X1 U897 ( .A1(G119), .A2(n925), .ZN(n801) );
  NAND2_X1 U898 ( .A1(n802), .A2(n801), .ZN(n806) );
  NAND2_X1 U899 ( .A1(G95), .A2(n922), .ZN(n804) );
  NAND2_X1 U900 ( .A1(G107), .A2(n926), .ZN(n803) );
  NAND2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n938) );
  XNOR2_X1 U903 ( .A(KEYINPUT89), .B(G1991), .ZN(n1043) );
  NOR2_X1 U904 ( .A1(n938), .A2(n1043), .ZN(n817) );
  NAND2_X1 U905 ( .A1(n922), .A2(G105), .ZN(n808) );
  XNOR2_X1 U906 ( .A(KEYINPUT38), .B(KEYINPUT90), .ZN(n807) );
  XNOR2_X1 U907 ( .A(n808), .B(n807), .ZN(n815) );
  NAND2_X1 U908 ( .A1(G129), .A2(n925), .ZN(n810) );
  NAND2_X1 U909 ( .A1(G117), .A2(n926), .ZN(n809) );
  NAND2_X1 U910 ( .A1(n810), .A2(n809), .ZN(n813) );
  NAND2_X1 U911 ( .A1(G141), .A2(n921), .ZN(n811) );
  XNOR2_X1 U912 ( .A(KEYINPUT91), .B(n811), .ZN(n812) );
  NOR2_X1 U913 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U914 ( .A1(n815), .A2(n814), .ZN(n920) );
  AND2_X1 U915 ( .A1(n920), .A2(G1996), .ZN(n816) );
  NOR2_X1 U916 ( .A1(n817), .A2(n816), .ZN(n973) );
  NOR2_X1 U917 ( .A1(n549), .A2(n819), .ZN(n864) );
  INV_X1 U918 ( .A(n864), .ZN(n820) );
  NOR2_X1 U919 ( .A1(n973), .A2(n820), .ZN(n856) );
  INV_X1 U920 ( .A(n856), .ZN(n832) );
  NAND2_X1 U921 ( .A1(n925), .A2(G128), .ZN(n821) );
  XOR2_X1 U922 ( .A(KEYINPUT87), .B(n821), .Z(n823) );
  NAND2_X1 U923 ( .A1(n926), .A2(G116), .ZN(n822) );
  NAND2_X1 U924 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U925 ( .A(n824), .B(KEYINPUT35), .ZN(n829) );
  NAND2_X1 U926 ( .A1(G140), .A2(n921), .ZN(n826) );
  NAND2_X1 U927 ( .A1(G104), .A2(n922), .ZN(n825) );
  NAND2_X1 U928 ( .A1(n826), .A2(n825), .ZN(n827) );
  XOR2_X1 U929 ( .A(KEYINPUT34), .B(n827), .Z(n828) );
  NAND2_X1 U930 ( .A1(n829), .A2(n828), .ZN(n830) );
  XOR2_X1 U931 ( .A(n830), .B(KEYINPUT36), .Z(n941) );
  XNOR2_X1 U932 ( .A(KEYINPUT37), .B(G2067), .ZN(n862) );
  OR2_X1 U933 ( .A1(n941), .A2(n862), .ZN(n831) );
  XOR2_X1 U934 ( .A(KEYINPUT88), .B(n831), .Z(n967) );
  NAND2_X1 U935 ( .A1(n864), .A2(n967), .ZN(n860) );
  AND2_X1 U936 ( .A1(n832), .A2(n860), .ZN(n849) );
  NAND2_X1 U937 ( .A1(n833), .A2(n849), .ZN(n834) );
  NOR2_X1 U938 ( .A1(n1010), .A2(n834), .ZN(n835) );
  NAND2_X1 U939 ( .A1(n836), .A2(n835), .ZN(n851) );
  NOR2_X1 U940 ( .A1(G1981), .A2(G305), .ZN(n837) );
  XOR2_X1 U941 ( .A(n837), .B(KEYINPUT93), .Z(n838) );
  XNOR2_X1 U942 ( .A(KEYINPUT24), .B(n838), .ZN(n839) );
  NAND2_X1 U943 ( .A1(n839), .A2(n845), .ZN(n847) );
  NOR2_X1 U944 ( .A1(n840), .A2(n841), .ZN(n844) );
  NAND2_X1 U945 ( .A1(G166), .A2(G8), .ZN(n842) );
  NOR2_X1 U946 ( .A1(G2090), .A2(n842), .ZN(n843) );
  NOR2_X1 U947 ( .A1(n844), .A2(n843), .ZN(n846) );
  NAND2_X1 U948 ( .A1(n847), .A2(n558), .ZN(n848) );
  NAND2_X1 U949 ( .A1(n849), .A2(n848), .ZN(n850) );
  XNOR2_X1 U950 ( .A(G1986), .B(G290), .ZN(n1014) );
  NOR2_X1 U951 ( .A1(G1996), .A2(n920), .ZN(n962) );
  AND2_X1 U952 ( .A1(n1043), .A2(n938), .ZN(n969) );
  NOR2_X1 U953 ( .A1(G1986), .A2(G290), .ZN(n853) );
  NOR2_X1 U954 ( .A1(n969), .A2(n853), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n854), .B(KEYINPUT102), .ZN(n855) );
  NOR2_X1 U956 ( .A1(n856), .A2(n855), .ZN(n857) );
  NOR2_X1 U957 ( .A1(n962), .A2(n857), .ZN(n858) );
  XOR2_X1 U958 ( .A(KEYINPUT39), .B(n858), .Z(n859) );
  XNOR2_X1 U959 ( .A(n859), .B(KEYINPUT103), .ZN(n861) );
  NAND2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n863) );
  NAND2_X1 U961 ( .A1(n941), .A2(n862), .ZN(n972) );
  NAND2_X1 U962 ( .A1(n863), .A2(n972), .ZN(n865) );
  NAND2_X1 U963 ( .A1(n865), .A2(n864), .ZN(n866) );
  XNOR2_X1 U964 ( .A(n867), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U965 ( .A1(G2106), .A2(n868), .ZN(G217) );
  AND2_X1 U966 ( .A1(G15), .A2(G2), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G661), .A2(n869), .ZN(G259) );
  NAND2_X1 U968 ( .A1(G3), .A2(G1), .ZN(n870) );
  NAND2_X1 U969 ( .A1(n871), .A2(n870), .ZN(G188) );
  XNOR2_X1 U970 ( .A(G120), .B(KEYINPUT105), .ZN(G236) );
  XNOR2_X1 U971 ( .A(G108), .B(KEYINPUT119), .ZN(G238) );
  INV_X1 U973 ( .A(G96), .ZN(G221) );
  NOR2_X1 U974 ( .A1(n873), .A2(n872), .ZN(G325) );
  INV_X1 U975 ( .A(G325), .ZN(G261) );
  NOR2_X1 U976 ( .A1(G860), .A2(n874), .ZN(n875) );
  XOR2_X1 U977 ( .A(n945), .B(n875), .Z(G145) );
  XOR2_X1 U978 ( .A(KEYINPUT106), .B(n876), .Z(G319) );
  XNOR2_X1 U979 ( .A(G2067), .B(G2072), .ZN(n877) );
  XNOR2_X1 U980 ( .A(n877), .B(KEYINPUT42), .ZN(n887) );
  XOR2_X1 U981 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n879) );
  XNOR2_X1 U982 ( .A(G2678), .B(G2096), .ZN(n878) );
  XNOR2_X1 U983 ( .A(n879), .B(n878), .ZN(n883) );
  XOR2_X1 U984 ( .A(G2100), .B(G2090), .Z(n881) );
  XNOR2_X1 U985 ( .A(G2084), .B(G2078), .ZN(n880) );
  XNOR2_X1 U986 ( .A(n881), .B(n880), .ZN(n882) );
  XOR2_X1 U987 ( .A(n883), .B(n882), .Z(n885) );
  XNOR2_X1 U988 ( .A(KEYINPUT109), .B(KEYINPUT43), .ZN(n884) );
  XNOR2_X1 U989 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U990 ( .A(n887), .B(n886), .ZN(G227) );
  XOR2_X1 U991 ( .A(KEYINPUT111), .B(G1956), .Z(n889) );
  XNOR2_X1 U992 ( .A(G1981), .B(G1961), .ZN(n888) );
  XNOR2_X1 U993 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U994 ( .A(n890), .B(KEYINPUT41), .Z(n892) );
  XNOR2_X1 U995 ( .A(G1996), .B(G1991), .ZN(n891) );
  XNOR2_X1 U996 ( .A(n892), .B(n891), .ZN(n896) );
  XOR2_X1 U997 ( .A(G1976), .B(G1971), .Z(n894) );
  XNOR2_X1 U998 ( .A(G1986), .B(G1966), .ZN(n893) );
  XNOR2_X1 U999 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U1000 ( .A(n896), .B(n895), .Z(n898) );
  XNOR2_X1 U1001 ( .A(KEYINPUT110), .B(G2474), .ZN(n897) );
  XNOR2_X1 U1002 ( .A(n898), .B(n897), .ZN(G229) );
  NAND2_X1 U1003 ( .A1(G100), .A2(n922), .ZN(n900) );
  NAND2_X1 U1004 ( .A1(G112), .A2(n926), .ZN(n899) );
  NAND2_X1 U1005 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U1006 ( .A(KEYINPUT112), .B(n901), .ZN(n906) );
  NAND2_X1 U1007 ( .A1(G124), .A2(n925), .ZN(n902) );
  XNOR2_X1 U1008 ( .A(n902), .B(KEYINPUT44), .ZN(n904) );
  NAND2_X1 U1009 ( .A1(n921), .A2(G136), .ZN(n903) );
  NAND2_X1 U1010 ( .A1(n904), .A2(n903), .ZN(n905) );
  NOR2_X1 U1011 ( .A1(n906), .A2(n905), .ZN(G162) );
  XNOR2_X1 U1012 ( .A(KEYINPUT115), .B(KEYINPUT45), .ZN(n911) );
  NAND2_X1 U1013 ( .A1(n922), .A2(G106), .ZN(n907) );
  XNOR2_X1 U1014 ( .A(n907), .B(KEYINPUT114), .ZN(n909) );
  NAND2_X1 U1015 ( .A1(G142), .A2(n921), .ZN(n908) );
  NAND2_X1 U1016 ( .A1(n909), .A2(n908), .ZN(n910) );
  XNOR2_X1 U1017 ( .A(n911), .B(n910), .ZN(n916) );
  NAND2_X1 U1018 ( .A1(G130), .A2(n925), .ZN(n913) );
  NAND2_X1 U1019 ( .A1(G118), .A2(n926), .ZN(n912) );
  NAND2_X1 U1020 ( .A1(n913), .A2(n912), .ZN(n914) );
  XOR2_X1 U1021 ( .A(KEYINPUT113), .B(n914), .Z(n915) );
  NOR2_X1 U1022 ( .A1(n916), .A2(n915), .ZN(n917) );
  XOR2_X1 U1023 ( .A(n917), .B(n968), .Z(n919) );
  XNOR2_X1 U1024 ( .A(G164), .B(G162), .ZN(n918) );
  XNOR2_X1 U1025 ( .A(n919), .B(n918), .ZN(n934) );
  XOR2_X1 U1026 ( .A(G160), .B(n920), .Z(n932) );
  NAND2_X1 U1027 ( .A1(G139), .A2(n921), .ZN(n924) );
  NAND2_X1 U1028 ( .A1(G103), .A2(n922), .ZN(n923) );
  NAND2_X1 U1029 ( .A1(n924), .A2(n923), .ZN(n931) );
  NAND2_X1 U1030 ( .A1(G127), .A2(n925), .ZN(n928) );
  NAND2_X1 U1031 ( .A1(G115), .A2(n926), .ZN(n927) );
  NAND2_X1 U1032 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1033 ( .A(KEYINPUT47), .B(n929), .Z(n930) );
  NOR2_X1 U1034 ( .A1(n931), .A2(n930), .ZN(n957) );
  XNOR2_X1 U1035 ( .A(n932), .B(n957), .ZN(n933) );
  XOR2_X1 U1036 ( .A(n934), .B(n933), .Z(n940) );
  XOR2_X1 U1037 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n936) );
  XNOR2_X1 U1038 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n935) );
  XNOR2_X1 U1039 ( .A(n936), .B(n935), .ZN(n937) );
  XNOR2_X1 U1040 ( .A(n938), .B(n937), .ZN(n939) );
  XNOR2_X1 U1041 ( .A(n940), .B(n939), .ZN(n942) );
  XNOR2_X1 U1042 ( .A(n942), .B(n941), .ZN(n943) );
  NOR2_X1 U1043 ( .A1(G37), .A2(n943), .ZN(G395) );
  XNOR2_X1 U1044 ( .A(G286), .B(n944), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(G171), .B(n1022), .ZN(n946) );
  XNOR2_X1 U1046 ( .A(n946), .B(n945), .ZN(n947) );
  XNOR2_X1 U1047 ( .A(n948), .B(n947), .ZN(n949) );
  XOR2_X1 U1048 ( .A(n949), .B(n1017), .Z(n950) );
  NOR2_X1 U1049 ( .A1(G37), .A2(n950), .ZN(G397) );
  NOR2_X1 U1050 ( .A1(G227), .A2(G229), .ZN(n951) );
  XOR2_X1 U1051 ( .A(KEYINPUT49), .B(n951), .Z(n952) );
  NAND2_X1 U1052 ( .A1(G319), .A2(n952), .ZN(n953) );
  NOR2_X1 U1053 ( .A1(G401), .A2(n953), .ZN(n956) );
  NOR2_X1 U1054 ( .A1(G395), .A2(G397), .ZN(n954) );
  XNOR2_X1 U1055 ( .A(n954), .B(KEYINPUT118), .ZN(n955) );
  NAND2_X1 U1056 ( .A1(n956), .A2(n955), .ZN(G225) );
  INV_X1 U1057 ( .A(G225), .ZN(G308) );
  INV_X1 U1058 ( .A(G57), .ZN(G237) );
  INV_X1 U1059 ( .A(KEYINPUT55), .ZN(n1058) );
  XOR2_X1 U1060 ( .A(G2072), .B(n957), .Z(n959) );
  XOR2_X1 U1061 ( .A(G164), .B(G2078), .Z(n958) );
  NOR2_X1 U1062 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1063 ( .A(KEYINPUT50), .B(n960), .ZN(n965) );
  XOR2_X1 U1064 ( .A(G2090), .B(G162), .Z(n961) );
  NOR2_X1 U1065 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1066 ( .A(KEYINPUT51), .B(n963), .Z(n964) );
  NAND2_X1 U1067 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1068 ( .A1(n967), .A2(n966), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(G160), .B(G2084), .ZN(n971) );
  NOR2_X1 U1070 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1071 ( .A1(n971), .A2(n970), .ZN(n975) );
  NAND2_X1 U1072 ( .A1(n973), .A2(n972), .ZN(n974) );
  NOR2_X1 U1073 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1074 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1075 ( .A(KEYINPUT52), .B(n978), .ZN(n979) );
  XOR2_X1 U1076 ( .A(KEYINPUT120), .B(n979), .Z(n980) );
  NAND2_X1 U1077 ( .A1(n1058), .A2(n980), .ZN(n981) );
  NAND2_X1 U1078 ( .A1(n981), .A2(G29), .ZN(n1038) );
  XNOR2_X1 U1079 ( .A(KEYINPUT125), .B(G1966), .ZN(n982) );
  XNOR2_X1 U1080 ( .A(n982), .B(G21), .ZN(n995) );
  XNOR2_X1 U1081 ( .A(G20), .B(n983), .ZN(n987) );
  XNOR2_X1 U1082 ( .A(G1981), .B(G6), .ZN(n985) );
  XNOR2_X1 U1083 ( .A(G1341), .B(G19), .ZN(n984) );
  NOR2_X1 U1084 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1085 ( .A1(n987), .A2(n986), .ZN(n990) );
  XOR2_X1 U1086 ( .A(KEYINPUT59), .B(G1348), .Z(n988) );
  XNOR2_X1 U1087 ( .A(G4), .B(n988), .ZN(n989) );
  NOR2_X1 U1088 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1089 ( .A(KEYINPUT60), .B(n991), .Z(n993) );
  XNOR2_X1 U1090 ( .A(G1961), .B(G5), .ZN(n992) );
  NOR2_X1 U1091 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1092 ( .A1(n995), .A2(n994), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(G1986), .B(G24), .ZN(n997) );
  XNOR2_X1 U1094 ( .A(G23), .B(G1976), .ZN(n996) );
  NOR2_X1 U1095 ( .A1(n997), .A2(n996), .ZN(n1000) );
  XOR2_X1 U1096 ( .A(G1971), .B(KEYINPUT126), .Z(n998) );
  XNOR2_X1 U1097 ( .A(G22), .B(n998), .ZN(n999) );
  NAND2_X1 U1098 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1099 ( .A(KEYINPUT58), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1100 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1101 ( .A(n1004), .B(KEYINPUT61), .ZN(n1005) );
  XNOR2_X1 U1102 ( .A(n1005), .B(KEYINPUT127), .ZN(n1007) );
  XNOR2_X1 U1103 ( .A(G16), .B(KEYINPUT124), .ZN(n1006) );
  NOR2_X1 U1104 ( .A1(n1007), .A2(n1006), .ZN(n1036) );
  XNOR2_X1 U1105 ( .A(G16), .B(KEYINPUT56), .ZN(n1008) );
  XNOR2_X1 U1106 ( .A(n1008), .B(KEYINPUT121), .ZN(n1033) );
  XOR2_X1 U1107 ( .A(G168), .B(G1966), .Z(n1009) );
  NOR2_X1 U1108 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1109 ( .A(KEYINPUT57), .B(n1011), .Z(n1021) );
  XNOR2_X1 U1110 ( .A(n1012), .B(G1956), .ZN(n1016) );
  XNOR2_X1 U1111 ( .A(G1961), .B(G301), .ZN(n1013) );
  NOR2_X1 U1112 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1113 ( .A1(n1016), .A2(n1015), .ZN(n1019) );
  XNOR2_X1 U1114 ( .A(G1348), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1115 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1116 ( .A1(n1021), .A2(n1020), .ZN(n1031) );
  XNOR2_X1 U1117 ( .A(G1341), .B(KEYINPUT122), .ZN(n1023) );
  XNOR2_X1 U1118 ( .A(n1023), .B(n1022), .ZN(n1027) );
  NAND2_X1 U1119 ( .A1(G1971), .A2(G303), .ZN(n1024) );
  NAND2_X1 U1120 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1121 ( .A1(n1027), .A2(n1026), .ZN(n1029) );
  NAND2_X1 U1122 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1123 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1124 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XOR2_X1 U1125 ( .A(KEYINPUT123), .B(n1034), .Z(n1035) );
  NOR2_X1 U1126 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1127 ( .A1(n1038), .A2(n1037), .ZN(n1063) );
  XNOR2_X1 U1128 ( .A(G2090), .B(G35), .ZN(n1053) );
  XNOR2_X1 U1129 ( .A(G32), .B(n1039), .ZN(n1040) );
  NAND2_X1 U1130 ( .A1(n1040), .A2(G28), .ZN(n1050) );
  XNOR2_X1 U1131 ( .A(G2067), .B(G26), .ZN(n1042) );
  XNOR2_X1 U1132 ( .A(G33), .B(G2072), .ZN(n1041) );
  NOR2_X1 U1133 ( .A1(n1042), .A2(n1041), .ZN(n1048) );
  XOR2_X1 U1134 ( .A(n1043), .B(G25), .Z(n1046) );
  XNOR2_X1 U1135 ( .A(G27), .B(n1044), .ZN(n1045) );
  NOR2_X1 U1136 ( .A1(n1046), .A2(n1045), .ZN(n1047) );
  NAND2_X1 U1137 ( .A1(n1048), .A2(n1047), .ZN(n1049) );
  NOR2_X1 U1138 ( .A1(n1050), .A2(n1049), .ZN(n1051) );
  XNOR2_X1 U1139 ( .A(KEYINPUT53), .B(n1051), .ZN(n1052) );
  NOR2_X1 U1140 ( .A1(n1053), .A2(n1052), .ZN(n1056) );
  XOR2_X1 U1141 ( .A(G2084), .B(G34), .Z(n1054) );
  XNOR2_X1 U1142 ( .A(KEYINPUT54), .B(n1054), .ZN(n1055) );
  NAND2_X1 U1143 ( .A1(n1056), .A2(n1055), .ZN(n1057) );
  XNOR2_X1 U1144 ( .A(n1058), .B(n1057), .ZN(n1060) );
  INV_X1 U1145 ( .A(G29), .ZN(n1059) );
  NAND2_X1 U1146 ( .A1(n1060), .A2(n1059), .ZN(n1061) );
  NAND2_X1 U1147 ( .A1(G11), .A2(n1061), .ZN(n1062) );
  NOR2_X1 U1148 ( .A1(n1063), .A2(n1062), .ZN(n1064) );
  XNOR2_X1 U1149 ( .A(n1064), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1150 ( .A(G311), .ZN(G150) );
endmodule

