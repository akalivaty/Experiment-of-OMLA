//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 0 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 1 0 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1297,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(new_n203), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT64), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n208), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G107), .ZN(new_n222));
  INV_X1    g0022(.A(G264), .ZN(new_n223));
  OAI22_X1  g0023(.A1(new_n220), .A2(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(G87), .B2(G250), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT66), .B(G68), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT67), .B(G238), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n225), .B(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT65), .Z(new_n231));
  OAI21_X1  g0031(.A(new_n210), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n213), .B(new_n219), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT69), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT68), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n238), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT70), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G41), .ZN(new_n253));
  INV_X1    g0053(.A(G45), .ZN(new_n254));
  AOI21_X1  g0054(.A(G1), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G1), .A3(G13), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n255), .A2(new_n257), .A3(G274), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT71), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G274), .ZN(new_n261));
  INV_X1    g0061(.A(new_n217), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n261), .B1(new_n262), .B2(new_n256), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(KEYINPUT71), .A3(new_n255), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n255), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n260), .A2(new_n264), .B1(G238), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G97), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT78), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT78), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(G33), .A3(G97), .ZN(new_n271));
  AND2_X1   g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G33), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n274), .A2(new_n276), .A3(G226), .A4(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n274), .A2(new_n276), .ZN(new_n280));
  INV_X1    g0080(.A(G232), .ZN(new_n281));
  NOR3_X1   g0081(.A1(new_n280), .A2(new_n281), .A3(new_n277), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n265), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT13), .ZN(new_n284));
  AND3_X1   g0084(.A1(new_n267), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n284), .B1(new_n267), .B2(new_n283), .ZN(new_n286));
  OAI21_X1  g0086(.A(G169), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT14), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT14), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n289), .B(G169), .C1(new_n285), .C2(new_n286), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n267), .A2(new_n283), .A3(new_n284), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(KEYINPUT79), .ZN(new_n292));
  INV_X1    g0092(.A(new_n286), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT79), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n267), .A2(new_n283), .A3(new_n294), .A4(new_n284), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n292), .A2(new_n293), .A3(G179), .A4(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n288), .A2(new_n290), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n227), .A2(G20), .ZN(new_n298));
  INV_X1    g0098(.A(G13), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(G1), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT12), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n299), .A2(new_n208), .A3(G1), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(KEYINPUT12), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT12), .ZN(new_n306));
  NAND3_X1  g0106(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n217), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  OR3_X1    g0109(.A1(new_n208), .A2(KEYINPUT74), .A3(G1), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT74), .B1(new_n208), .B2(G1), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n306), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n305), .B1(new_n203), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT80), .ZN(new_n315));
  INV_X1    g0115(.A(new_n308), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n273), .A2(G20), .ZN(new_n317));
  NOR2_X1   g0117(.A1(G20), .A2(G33), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n317), .A2(G77), .B1(new_n318), .B2(G50), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n316), .B1(new_n298), .B2(new_n319), .ZN(new_n320));
  XOR2_X1   g0120(.A(new_n320), .B(KEYINPUT11), .Z(new_n321));
  INV_X1    g0121(.A(KEYINPUT80), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n305), .B(new_n322), .C1(new_n203), .C2(new_n313), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n315), .A2(new_n321), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n297), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G200), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(new_n293), .B2(new_n291), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(new_n324), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n292), .A2(new_n293), .A3(G190), .A4(new_n295), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT3), .B(G33), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(G222), .A3(new_n277), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(G223), .A3(G1698), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n280), .A2(G77), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n265), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n260), .A2(new_n264), .B1(G226), .B2(new_n266), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n338), .B1(new_n339), .B2(KEYINPUT72), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n260), .A2(new_n264), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n266), .A2(G226), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n341), .A2(KEYINPUT72), .A3(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT73), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n341), .A2(new_n342), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT72), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n339), .A2(KEYINPUT72), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT73), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n347), .A2(new_n348), .A3(new_n349), .A4(new_n338), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G179), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n309), .A2(new_n312), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G50), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n204), .A2(G20), .ZN(new_n357));
  INV_X1    g0157(.A(G150), .ZN(new_n358));
  INV_X1    g0158(.A(new_n318), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n208), .A2(G33), .ZN(new_n360));
  XNOR2_X1  g0160(.A(KEYINPUT8), .B(G58), .ZN(new_n361));
  OAI221_X1 g0161(.A(new_n357), .B1(new_n358), .B2(new_n359), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n362), .A2(new_n308), .B1(new_n201), .B2(new_n303), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n354), .A2(KEYINPUT75), .B1(new_n356), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(KEYINPUT75), .B1(new_n351), .B2(G169), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n353), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n344), .A2(new_n350), .A3(G200), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n363), .A2(new_n356), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n369), .B(KEYINPUT9), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G190), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(new_n344), .B2(new_n350), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT10), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n351), .A2(G190), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT10), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n375), .A2(new_n376), .A3(new_n368), .A4(new_n370), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G20), .A2(G77), .ZN(new_n379));
  XNOR2_X1  g0179(.A(KEYINPUT15), .B(G87), .ZN(new_n380));
  OAI221_X1 g0180(.A(new_n379), .B1(new_n380), .B2(new_n360), .C1(new_n359), .C2(new_n361), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n308), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n355), .A2(G77), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n303), .A2(new_n220), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT77), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n381), .A2(new_n308), .B1(new_n220), .B2(new_n303), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n388), .A2(KEYINPUT77), .A3(new_n383), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n333), .A2(G1698), .ZN(new_n391));
  OAI22_X1  g0191(.A1(new_n391), .A2(new_n228), .B1(new_n222), .B2(new_n333), .ZN(new_n392));
  NOR3_X1   g0192(.A1(new_n280), .A2(new_n281), .A3(G1698), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n265), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n260), .A2(new_n264), .B1(G244), .B2(new_n266), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G169), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n394), .A2(new_n352), .A3(new_n395), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n390), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n396), .A2(G200), .ZN(new_n402));
  INV_X1    g0202(.A(new_n396), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n402), .A2(KEYINPUT76), .B1(new_n403), .B2(G190), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n394), .A2(KEYINPUT76), .A3(G190), .A4(new_n395), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n387), .A2(new_n389), .A3(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n332), .A2(new_n367), .A3(new_n378), .A4(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n361), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n410), .A2(new_n303), .ZN(new_n411));
  INV_X1    g0211(.A(new_n355), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n411), .B1(new_n412), .B2(new_n410), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(KEYINPUT7), .B1(new_n280), .B2(new_n208), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT7), .ZN(new_n416));
  AOI211_X1 g0216(.A(new_n416), .B(G20), .C1(new_n274), .C2(new_n276), .ZN(new_n417));
  OAI21_X1  g0217(.A(G68), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(G159), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n359), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n214), .B1(new_n227), .B2(new_n202), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n420), .B1(new_n421), .B2(G20), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n418), .A2(KEYINPUT16), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n227), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n415), .B2(new_n417), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT16), .B1(new_n425), .B2(new_n422), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT81), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n308), .B(new_n423), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT16), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n421), .A2(G20), .ZN(new_n430));
  INV_X1    g0230(.A(new_n420), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n416), .B1(new_n333), .B2(G20), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n280), .A2(KEYINPUT7), .A3(new_n208), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n227), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n429), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n436), .A2(KEYINPUT81), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n414), .B1(new_n428), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT82), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n436), .A2(KEYINPUT81), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n426), .A2(new_n427), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n441), .A2(new_n442), .A3(new_n308), .A4(new_n423), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(KEYINPUT82), .A3(new_n414), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n274), .A2(new_n276), .A3(G226), .A4(G1698), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n274), .A2(new_n276), .A3(G223), .A4(new_n277), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G87), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT83), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT83), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n445), .A2(new_n446), .A3(new_n450), .A4(new_n447), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n265), .A3(new_n451), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n260), .A2(new_n264), .B1(G232), .B2(new_n266), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G169), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n452), .A2(G179), .A3(new_n453), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n440), .A2(new_n444), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(KEYINPUT18), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT17), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n452), .A2(G190), .A3(new_n453), .ZN(new_n461));
  INV_X1    g0261(.A(new_n454), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n461), .B1(new_n462), .B2(new_n327), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n460), .B1(new_n438), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n327), .B1(new_n452), .B2(new_n453), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n465), .B1(new_n462), .B2(G190), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n466), .A2(new_n443), .A3(KEYINPUT17), .A4(new_n414), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT18), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n440), .A2(new_n444), .A3(new_n469), .A4(new_n457), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n459), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n409), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n309), .B1(G1), .B2(new_n273), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n303), .ZN(new_n475));
  OR3_X1    g0275(.A1(new_n475), .A2(KEYINPUT85), .A3(G97), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT85), .B1(new_n475), .B2(G97), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n474), .A2(G97), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(G107), .B1(new_n415), .B2(new_n417), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT6), .ZN(new_n480));
  AND2_X1   g0280(.A1(G97), .A2(G107), .ZN(new_n481));
  NOR2_X1   g0281(.A1(G97), .A2(G107), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n222), .A2(KEYINPUT6), .A3(G97), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n485), .A2(G20), .B1(G77), .B2(new_n318), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n316), .B1(new_n479), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(KEYINPUT84), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT84), .ZN(new_n489));
  AOI211_X1 g0289(.A(new_n489), .B(new_n316), .C1(new_n479), .C2(new_n486), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n478), .B1(new_n488), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n274), .A2(new_n276), .A3(G244), .A4(new_n277), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT86), .ZN(new_n495));
  OR2_X1    g0295(.A1(new_n492), .A2(new_n493), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT86), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n492), .A2(new_n497), .A3(new_n493), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n274), .A2(new_n276), .A3(G250), .A4(G1698), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G283), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n495), .A2(new_n496), .A3(new_n498), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n265), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n207), .A2(G45), .ZN(new_n504));
  NOR2_X1   g0304(.A1(KEYINPUT5), .A2(G41), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(KEYINPUT5), .A2(G41), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n263), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n254), .A2(G1), .ZN(new_n510));
  INV_X1    g0310(.A(new_n507), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n510), .B1(new_n511), .B2(new_n505), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n257), .ZN(new_n513));
  INV_X1    g0313(.A(G257), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n509), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n503), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n397), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n515), .B1(new_n502), .B2(new_n265), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n352), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n491), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n485), .A2(G20), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n318), .A2(G77), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n222), .B1(new_n433), .B2(new_n434), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n308), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n489), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n487), .A2(KEYINPUT84), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n519), .A2(G200), .ZN(new_n530));
  AOI211_X1 g0330(.A(G190), .B(new_n515), .C1(new_n502), .C2(new_n265), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n529), .B(new_n478), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n274), .A2(new_n276), .A3(G244), .A4(G1698), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n274), .A2(new_n276), .A3(G238), .A4(new_n277), .ZN(new_n534));
  INV_X1    g0334(.A(G116), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n533), .B(new_n534), .C1(new_n273), .C2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n265), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n257), .A2(G274), .A3(new_n510), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n257), .A2(G250), .A3(new_n504), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n327), .B1(new_n537), .B2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(G87), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n482), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT19), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n545), .B1(new_n269), .B2(new_n271), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n544), .B1(new_n546), .B2(G20), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n274), .A2(new_n276), .A3(new_n208), .A4(G68), .ZN(new_n548));
  INV_X1    g0348(.A(G97), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n545), .B1(new_n360), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n316), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n380), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(new_n475), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n473), .A2(new_n543), .ZN(new_n555));
  NOR4_X1   g0355(.A1(new_n542), .A2(new_n552), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT87), .ZN(new_n557));
  AND4_X1   g0357(.A1(new_n557), .A2(new_n537), .A3(G190), .A4(new_n541), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n540), .B1(new_n536), .B2(new_n265), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n557), .B1(new_n559), .B2(G190), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n552), .A2(new_n554), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n473), .B2(new_n380), .ZN(new_n563));
  AOI211_X1 g0363(.A(G179), .B(new_n540), .C1(new_n265), .C2(new_n536), .ZN(new_n564));
  AOI21_X1  g0364(.A(G169), .B1(new_n537), .B2(new_n541), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n556), .A2(new_n561), .B1(new_n563), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n521), .A2(new_n532), .A3(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT21), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n303), .A2(G116), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n570), .B1(new_n473), .B2(G116), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT90), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n500), .B(new_n208), .C1(G33), .C2(new_n549), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n535), .A2(G20), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n308), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(KEYINPUT88), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT88), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n308), .A2(new_n578), .A3(new_n575), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n574), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n572), .B1(new_n580), .B2(KEYINPUT20), .ZN(new_n581));
  INV_X1    g0381(.A(new_n579), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n578), .B1(new_n308), .B2(new_n575), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n573), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT20), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(KEYINPUT90), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n581), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(KEYINPUT20), .B(new_n573), .C1(new_n582), .C2(new_n583), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT89), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n580), .A2(KEYINPUT89), .A3(KEYINPUT20), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n571), .B1(new_n587), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n508), .A2(new_n265), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n594), .A2(G270), .B1(new_n263), .B2(new_n508), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n274), .A2(new_n276), .A3(G264), .A4(G1698), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n274), .A2(new_n276), .A3(G257), .A4(new_n277), .ZN(new_n597));
  INV_X1    g0397(.A(G303), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n596), .B(new_n597), .C1(new_n598), .C2(new_n333), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n265), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n595), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(G169), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n569), .B1(new_n593), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n595), .A2(G179), .A3(new_n600), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(new_n602), .B2(new_n569), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n581), .A2(new_n586), .B1(new_n590), .B2(new_n591), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n605), .B1(new_n606), .B2(new_n571), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n601), .A2(G200), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n595), .A2(G190), .A3(new_n600), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n593), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n603), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(KEYINPUT92), .B1(new_n513), .B2(new_n223), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT92), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n512), .A2(new_n613), .A3(G264), .A4(new_n257), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n333), .A2(G257), .A3(G1698), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n333), .A2(G250), .A3(new_n277), .ZN(new_n616));
  NAND2_X1  g0416(.A1(G33), .A2(G294), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n612), .A2(new_n614), .B1(new_n618), .B2(new_n265), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n619), .A2(new_n352), .A3(new_n509), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n509), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n397), .ZN(new_n622));
  XNOR2_X1  g0422(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n333), .A2(new_n208), .A3(G87), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(KEYINPUT22), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT22), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n333), .A2(new_n627), .A3(new_n208), .A4(G87), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n273), .A2(new_n535), .A3(G20), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT23), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n631), .B1(new_n208), .B2(G107), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n222), .A2(KEYINPUT23), .A3(G20), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n624), .B1(new_n629), .B2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n629), .A2(new_n634), .A3(new_n624), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n316), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(KEYINPUT25), .B1(new_n303), .B2(new_n222), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n303), .A2(KEYINPUT25), .A3(new_n222), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n474), .A2(G107), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n620), .B(new_n622), .C1(new_n638), .C2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n637), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n308), .B1(new_n645), .B2(new_n635), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n619), .A2(new_n372), .A3(new_n509), .ZN(new_n647));
  AOI21_X1  g0447(.A(G200), .B1(new_n619), .B2(new_n509), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n646), .B(new_n642), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  NOR3_X1   g0450(.A1(new_n568), .A2(new_n611), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n472), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n652), .B(KEYINPUT93), .ZN(G372));
  NAND2_X1  g0453(.A1(new_n563), .A2(new_n566), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n644), .A2(new_n603), .A3(new_n607), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n521), .A2(new_n532), .A3(new_n567), .A4(new_n649), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  INV_X1    g0458(.A(new_n560), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n552), .A2(new_n555), .A3(new_n554), .ZN(new_n660));
  INV_X1    g0460(.A(new_n542), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n559), .A2(new_n557), .A3(G190), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n659), .A2(new_n660), .A3(new_n661), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n663), .A2(new_n654), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n658), .B1(new_n521), .B2(new_n664), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n529), .A2(new_n478), .B1(new_n352), .B2(new_n519), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n567), .A2(new_n666), .A3(KEYINPUT26), .A4(new_n518), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g0468(.A1(new_n657), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n472), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n438), .A2(new_n457), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT18), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n438), .A2(new_n469), .A3(new_n457), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT94), .ZN(new_n675));
  AND3_X1   g0475(.A1(new_n388), .A2(KEYINPUT77), .A3(new_n383), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT77), .B1(new_n388), .B2(new_n383), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n398), .A2(new_n399), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n675), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n390), .A2(KEYINPUT94), .A3(new_n398), .A4(new_n399), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n329), .A2(new_n330), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n326), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n464), .A2(new_n467), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n674), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT95), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n378), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n374), .A2(KEYINPUT95), .A3(new_n377), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI22_X1  g0490(.A1(new_n686), .A2(new_n690), .B1(new_n366), .B2(new_n364), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n670), .A2(new_n691), .ZN(G369));
  AND2_X1   g0492(.A1(new_n603), .A2(new_n607), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n300), .A2(new_n208), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(KEYINPUT27), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G213), .A3(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G343), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n606), .B2(new_n571), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n693), .A2(new_n700), .ZN(new_n701));
  AND3_X1   g0501(.A1(new_n603), .A2(new_n607), .A3(new_n610), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n700), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT96), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g0506(.A(KEYINPUT97), .B(G330), .ZN(new_n707));
  INV_X1    g0507(.A(new_n650), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n699), .B1(new_n638), .B2(new_n643), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n644), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n699), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n706), .A2(new_n707), .A3(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n693), .A2(new_n699), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n708), .ZN(new_n716));
  INV_X1    g0516(.A(new_n699), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n711), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n714), .A2(new_n720), .ZN(G399));
  INV_X1    g0521(.A(new_n211), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G41), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n544), .A2(G116), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n724), .A2(G1), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n216), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n726), .B1(new_n727), .B2(new_n724), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT28), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT29), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n521), .A2(new_n532), .A3(new_n567), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n603), .A2(new_n607), .ZN(new_n732));
  OAI211_X1 g0532(.A(new_n731), .B(new_n649), .C1(new_n732), .C2(new_n711), .ZN(new_n733));
  OAI211_X1 g0533(.A(KEYINPUT102), .B(new_n658), .C1(new_n521), .C2(new_n664), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT102), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n665), .A2(new_n667), .A3(new_n735), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n733), .A2(new_n654), .A3(new_n734), .A4(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n730), .B1(new_n737), .B2(new_n717), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n730), .B(new_n717), .C1(new_n657), .C2(new_n668), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT31), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n612), .A2(new_n614), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n618), .A2(new_n265), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n743), .A2(new_n559), .A3(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT98), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n619), .A2(KEYINPUT98), .A3(new_n559), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n604), .A2(KEYINPUT99), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT99), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n595), .A2(new_n600), .A3(new_n751), .A4(G179), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n749), .A2(KEYINPUT30), .A3(new_n753), .A4(new_n519), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n559), .A2(G179), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n517), .A2(new_n755), .A3(new_n601), .A4(new_n621), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n749), .A2(new_n519), .A3(new_n753), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT30), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(KEYINPUT101), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n517), .B1(new_n747), .B2(new_n748), .ZN(new_n762));
  AOI21_X1  g0562(.A(KEYINPUT30), .B1(new_n762), .B2(new_n753), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT101), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n757), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n742), .B1(new_n766), .B2(new_n717), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n731), .A2(new_n702), .A3(new_n708), .A4(new_n717), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n717), .A2(new_n742), .ZN(new_n769));
  OAI211_X1 g0569(.A(KEYINPUT100), .B(new_n769), .C1(new_n757), .C2(new_n763), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n769), .B1(new_n757), .B2(new_n763), .ZN(new_n771));
  INV_X1    g0571(.A(KEYINPUT100), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n767), .A2(new_n768), .A3(new_n770), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n707), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n741), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n729), .B1(new_n777), .B2(G1), .ZN(G364));
  AND2_X1   g0578(.A1(new_n701), .A2(new_n703), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(new_n705), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n704), .A2(KEYINPUT96), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n780), .A2(new_n707), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n299), .A2(G20), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n207), .B1(new_n783), .B2(G45), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n723), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n782), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n706), .A2(new_n707), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n779), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n211), .A2(new_n333), .ZN(new_n795));
  INV_X1    g0595(.A(G355), .ZN(new_n796));
  OAI22_X1  g0596(.A1(new_n795), .A2(new_n796), .B1(G116), .B2(new_n211), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n248), .A2(G45), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n722), .A2(new_n333), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(new_n216), .B2(new_n254), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n797), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n217), .B1(G20), .B2(new_n397), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n793), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n786), .B1(new_n802), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n208), .A2(new_n352), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n807), .A2(G190), .A3(G200), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(KEYINPUT103), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n808), .A2(KEYINPUT103), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(G50), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n372), .A2(G179), .A3(G200), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n208), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G97), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n208), .A2(G179), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n819), .A2(new_n372), .A3(G200), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n818), .B1(new_n222), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n807), .A2(new_n372), .A3(G200), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n819), .A2(G190), .A3(G200), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n822), .A2(new_n203), .B1(new_n823), .B2(new_n543), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(G190), .A2(G200), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n819), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n827), .A2(new_n419), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT32), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n807), .A2(G190), .A3(new_n327), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n333), .B1(new_n830), .B2(new_n202), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n807), .A2(new_n826), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n831), .B1(G77), .B2(new_n833), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n814), .A2(new_n825), .A3(new_n829), .A4(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(G294), .ZN(new_n836));
  INV_X1    g0636(.A(G311), .ZN(new_n837));
  OAI22_X1  g0637(.A1(new_n816), .A2(new_n836), .B1(new_n832), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(new_n813), .B2(G326), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT104), .Z(new_n840));
  INV_X1    g0640(.A(G322), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n280), .B1(new_n830), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n827), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n842), .B1(G329), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n822), .ZN(new_n845));
  INV_X1    g0645(.A(G317), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(KEYINPUT33), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n846), .A2(KEYINPUT33), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n845), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n823), .ZN(new_n850));
  INV_X1    g0650(.A(new_n820), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n850), .A2(G303), .B1(new_n851), .B2(G283), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n844), .A2(new_n849), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n835), .B1(new_n840), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n806), .B1(new_n854), .B2(new_n803), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n790), .B1(new_n794), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(G396));
  NAND2_X1  g0657(.A1(new_n669), .A2(new_n717), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n390), .A2(new_n699), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n680), .A2(new_n860), .A3(new_n681), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n400), .B(new_n859), .C1(new_n404), .C2(new_n406), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n861), .A2(new_n862), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n717), .B(new_n865), .C1(new_n657), .C2(new_n668), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n786), .B1(new_n867), .B2(new_n775), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n775), .B2(new_n867), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n803), .A2(new_n791), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n787), .B1(new_n220), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n830), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n872), .A2(G143), .B1(new_n833), .B2(G159), .ZN(new_n873));
  INV_X1    g0673(.A(G137), .ZN(new_n874));
  OAI221_X1 g0674(.A(new_n873), .B1(new_n358), .B2(new_n822), .C1(new_n812), .C2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n876), .A2(KEYINPUT34), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n876), .A2(KEYINPUT34), .ZN(new_n878));
  INV_X1    g0678(.A(G132), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n333), .B1(new_n827), .B2(new_n879), .C1(new_n203), .C2(new_n820), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n816), .A2(new_n202), .B1(new_n823), .B2(new_n201), .ZN(new_n881));
  NOR4_X1   g0681(.A1(new_n877), .A2(new_n878), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n845), .A2(G283), .B1(new_n833), .B2(G116), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n812), .B2(new_n598), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n884), .B(KEYINPUT105), .Z(new_n885));
  OAI221_X1 g0685(.A(new_n280), .B1(new_n827), .B2(new_n837), .C1(new_n830), .C2(new_n836), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n818), .B1(new_n543), .B2(new_n820), .C1(new_n222), .C2(new_n823), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n882), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n803), .ZN(new_n890));
  OAI221_X1 g0690(.A(new_n871), .B1(new_n865), .B2(new_n792), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n869), .A2(new_n891), .ZN(G384));
  OR2_X1    g0692(.A1(new_n485), .A2(KEYINPUT35), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n485), .A2(KEYINPUT35), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n893), .A2(G116), .A3(new_n218), .A4(new_n894), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT36), .ZN(new_n896));
  OAI21_X1  g0696(.A(G77), .B1(new_n227), .B2(new_n202), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n727), .A2(new_n897), .B1(G50), .B2(new_n203), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n898), .A2(G1), .A3(new_n299), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n899), .B(KEYINPUT106), .Z(new_n900));
  NAND2_X1  g0700(.A1(new_n324), .A2(new_n699), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n325), .A2(new_n683), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n901), .B1(new_n325), .B2(new_n683), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n865), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g0704(.A1(new_n754), .A2(new_n756), .ZN(new_n905));
  AOI211_X1 g0705(.A(KEYINPUT101), .B(KEYINPUT30), .C1(new_n762), .C2(new_n753), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n764), .B1(new_n758), .B2(new_n759), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n651), .A2(new_n717), .B1(new_n908), .B2(new_n769), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n904), .B1(new_n909), .B2(new_n767), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT38), .ZN(new_n911));
  INV_X1    g0711(.A(new_n697), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n440), .A2(new_n444), .A3(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n438), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT37), .B1(new_n914), .B2(new_n466), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n458), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n423), .A2(new_n308), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT16), .B1(new_n418), .B2(new_n422), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n414), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n457), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n912), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n920), .B(new_n921), .C1(new_n438), .C2(new_n463), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT37), .ZN(new_n923));
  INV_X1    g0723(.A(new_n921), .ZN(new_n924));
  AOI221_X4 g0724(.A(new_n911), .B1(new_n916), .B2(new_n923), .C1(new_n471), .C2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n471), .A2(new_n924), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n916), .A2(new_n923), .ZN(new_n927));
  AOI21_X1  g0727(.A(KEYINPUT38), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n910), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT40), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND4_X1  g0731(.A1(new_n672), .A2(new_n464), .A3(new_n467), .A4(new_n673), .ZN(new_n932));
  INV_X1    g0732(.A(new_n913), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n458), .A2(new_n913), .A3(new_n915), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT37), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n438), .A2(new_n463), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n443), .A2(new_n414), .B1(new_n455), .B2(new_n456), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n936), .B1(new_n939), .B2(new_n913), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n934), .B1(new_n935), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n911), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n926), .A2(KEYINPUT38), .A3(new_n927), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n325), .A2(new_n683), .A3(new_n901), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n324), .B(new_n699), .C1(new_n331), .C2(new_n297), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n863), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n769), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n768), .B1(new_n766), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT31), .B1(new_n908), .B2(new_n699), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n947), .B(KEYINPUT40), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n931), .B1(new_n944), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n472), .B1(new_n950), .B2(new_n949), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(new_n953), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n954), .A2(new_n707), .A3(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n325), .A2(new_n699), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT39), .B1(new_n925), .B2(new_n928), .ZN(new_n959));
  XNOR2_X1  g0759(.A(KEYINPUT107), .B(KEYINPUT39), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n942), .A2(new_n943), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n958), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n674), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n697), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n925), .A2(new_n928), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n401), .A2(new_n717), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n866), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n902), .A2(new_n903), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n964), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n962), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n472), .B1(new_n738), .B2(new_n740), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n691), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n972), .B(new_n974), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n956), .A2(new_n975), .B1(new_n207), .B2(new_n783), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n956), .A2(new_n975), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n896), .B(new_n900), .C1(new_n976), .C2(new_n977), .ZN(G367));
  OR2_X1    g0778(.A1(new_n238), .A2(new_n800), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n805), .B1(new_n722), .B2(new_n553), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n787), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n793), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n567), .B1(new_n660), .B2(new_n717), .ZN(new_n983));
  OR3_X1    g0783(.A1(new_n654), .A2(new_n660), .A3(new_n717), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G50), .A2(new_n833), .B1(new_n843), .B2(G137), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n986), .B(new_n333), .C1(new_n358), .C2(new_n830), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G159), .A2(new_n845), .B1(new_n851), .B2(G77), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n202), .B2(new_n823), .C1(new_n203), .C2(new_n816), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n987), .B(new_n989), .C1(G143), .C2(new_n813), .ZN(new_n990));
  AOI22_X1  g0790(.A1(G107), .A2(new_n817), .B1(new_n845), .B2(G294), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n549), .B2(new_n820), .C1(new_n812), .C2(new_n837), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT46), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n823), .A2(new_n993), .A3(new_n535), .ZN(new_n994));
  AOI22_X1  g0794(.A1(G283), .A2(new_n833), .B1(new_n843), .B2(G317), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n333), .B1(new_n872), .B2(G303), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n993), .B1(new_n823), .B2(new_n535), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  NOR3_X1   g0798(.A1(new_n992), .A2(new_n994), .A3(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n990), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT109), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT47), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n981), .B1(new_n982), .B2(new_n985), .C1(new_n1002), .C2(new_n890), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n491), .A2(new_n699), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n521), .A2(new_n532), .A3(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n666), .A2(new_n518), .A3(new_n699), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n719), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT44), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n720), .A2(KEYINPUT45), .A3(new_n1007), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT45), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n719), .B2(new_n1008), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n714), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1011), .A2(new_n714), .A3(new_n1015), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n716), .B1(new_n713), .B2(new_n715), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT108), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1020), .B1(new_n782), .B2(new_n1021), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n706), .A2(KEYINPUT108), .A3(new_n707), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n782), .A2(new_n1021), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1020), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1023), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n777), .B1(new_n1019), .B2(new_n1028), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n723), .B(KEYINPUT41), .Z(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n785), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1005), .A2(new_n644), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n699), .B1(new_n1033), .B2(new_n521), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n715), .A2(new_n708), .A3(new_n1007), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1034), .B1(KEYINPUT42), .B2(new_n1035), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1035), .A2(KEYINPUT42), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1036), .A2(new_n1037), .B1(KEYINPUT43), .B2(new_n985), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1038), .B(new_n1039), .Z(new_n1040));
  NOR2_X1   g0840(.A1(new_n714), .A2(new_n1008), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n1040), .B(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1003), .B1(new_n1032), .B2(new_n1043), .ZN(G387));
  AOI21_X1  g0844(.A(new_n1027), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1045), .A2(new_n1022), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n777), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n776), .B1(new_n1045), .B2(new_n1022), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n723), .B(KEYINPUT111), .Z(new_n1049));
  NAND3_X1  g0849(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n710), .A2(new_n712), .A3(new_n793), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n795), .A2(new_n725), .B1(G107), .B2(new_n211), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n243), .A2(new_n254), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n725), .ZN(new_n1054));
  AOI211_X1 g0854(.A(G45), .B(new_n1054), .C1(G68), .C2(G77), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n361), .A2(G50), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT50), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n800), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1052), .B1(new_n1053), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n786), .B1(new_n1059), .B2(new_n805), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n830), .A2(new_n201), .B1(new_n832), .B2(new_n203), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n280), .B(new_n1061), .C1(G150), .C2(new_n843), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n816), .A2(new_n380), .B1(new_n822), .B2(new_n361), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n220), .A2(new_n823), .B1(new_n820), .B2(new_n549), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT110), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n813), .B2(G159), .ZN(new_n1067));
  NOR3_X1   g0867(.A1(new_n812), .A2(KEYINPUT110), .A3(new_n419), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1062), .B(new_n1065), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n333), .B1(new_n843), .B2(G326), .ZN(new_n1070));
  INV_X1    g0870(.A(G283), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n816), .A2(new_n1071), .B1(new_n823), .B2(new_n836), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n872), .A2(G317), .B1(new_n833), .B2(G303), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n837), .B2(new_n822), .C1(new_n812), .C2(new_n841), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT48), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1072), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n1075), .B2(new_n1074), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT49), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1070), .B1(new_n535), .B2(new_n820), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1069), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1060), .B1(new_n1081), .B2(new_n803), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1046), .A2(new_n785), .B1(new_n1051), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1050), .A2(new_n1083), .ZN(G393));
  NOR2_X1   g0884(.A1(new_n1028), .A2(new_n776), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1018), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1086), .A2(new_n1016), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1047), .A2(new_n1019), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1088), .A2(new_n1049), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1008), .A2(new_n793), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n799), .A2(new_n251), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1092), .B(new_n804), .C1(new_n549), .C2(new_n211), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT112), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n787), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1095), .B1(new_n1094), .B2(new_n1093), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n812), .A2(new_n358), .B1(new_n419), .B2(new_n830), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT51), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n280), .B1(new_n843), .B2(G143), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n361), .B2(new_n832), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n816), .A2(new_n220), .B1(new_n822), .B2(new_n201), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n543), .A2(new_n820), .B1(new_n823), .B2(new_n227), .ZN(new_n1102));
  NOR3_X1   g0902(.A1(new_n1100), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n812), .A2(new_n846), .B1(new_n837), .B2(new_n830), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT52), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n280), .B1(new_n827), .B2(new_n841), .C1(new_n836), .C2(new_n832), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n822), .A2(new_n598), .B1(new_n820), .B2(new_n222), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n816), .A2(new_n535), .B1(new_n823), .B2(new_n1071), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1098), .A2(new_n1103), .B1(new_n1105), .B2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT113), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1096), .B1(new_n1111), .B2(new_n803), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1087), .A2(new_n785), .B1(new_n1091), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1090), .A2(new_n1113), .ZN(G390));
  NAND2_X1  g0914(.A1(new_n970), .A2(new_n958), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1115), .A2(new_n959), .A3(new_n961), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n942), .A2(new_n943), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n736), .A2(new_n734), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n717), .B(new_n865), .C1(new_n1118), .C2(new_n657), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1119), .A2(new_n966), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n958), .B(new_n1117), .C1(new_n1120), .C2(new_n968), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n774), .A2(new_n707), .A3(new_n865), .A4(new_n969), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1116), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(G330), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n909), .B2(new_n767), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n947), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n1116), .B2(new_n1121), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1123), .A2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(G330), .B(new_n865), .C1(new_n949), .C2(new_n950), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n968), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1122), .A2(new_n1130), .A3(new_n1120), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n773), .A2(new_n768), .A3(new_n770), .ZN(new_n1132));
  OAI211_X1 g0932(.A(new_n707), .B(new_n865), .C1(new_n1132), .C2(new_n950), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n968), .A2(new_n1133), .B1(new_n1125), .B2(new_n947), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n967), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1131), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1125), .A2(new_n472), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n973), .A2(new_n1137), .A3(new_n691), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT114), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n973), .A2(new_n1137), .A3(KEYINPUT114), .A4(new_n691), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1136), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1128), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1116), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1116), .A2(new_n1121), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1145), .B1(new_n1146), .B2(new_n1126), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n1142), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1144), .A2(new_n1148), .A3(new_n1049), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n959), .A2(new_n791), .A3(new_n961), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n870), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n786), .B1(new_n410), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n813), .A2(G283), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n830), .A2(new_n535), .B1(new_n827), .B2(new_n836), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n333), .B(new_n1154), .C1(G97), .C2(new_n833), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n850), .A2(G87), .B1(new_n851), .B2(G68), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G77), .A2(new_n817), .B1(new_n845), .B2(G107), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1153), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(G128), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n812), .A2(new_n1159), .B1(new_n879), .B2(new_n830), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT115), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n850), .A2(G150), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT53), .ZN(new_n1163));
  INV_X1    g0963(.A(G125), .ZN(new_n1164));
  XNOR2_X1  g0964(.A(KEYINPUT54), .B(G143), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n333), .B1(new_n827), .B2(new_n1164), .C1(new_n832), .C2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n816), .A2(new_n419), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n822), .A2(new_n874), .B1(new_n820), .B2(new_n201), .ZN(new_n1168));
  OR4_X1    g0968(.A1(new_n1163), .A2(new_n1166), .A3(new_n1167), .A4(new_n1168), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1158), .B1(new_n1161), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1152), .B1(new_n1170), .B2(new_n803), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1150), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n1147), .B2(new_n784), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1149), .A2(new_n1174), .ZN(G378));
  INV_X1    g0975(.A(new_n961), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT39), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n685), .B1(KEYINPUT18), .B2(new_n458), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n921), .B1(new_n1178), .B2(new_n470), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n927), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n911), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1177), .B1(new_n1181), .B2(new_n943), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n957), .B1(new_n1176), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n970), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1181), .A2(new_n943), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1184), .A2(new_n1185), .B1(new_n963), .B2(new_n697), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n951), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1124), .B1(new_n1188), .B2(new_n1117), .ZN(new_n1189));
  XOR2_X1   g0989(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n369), .A2(new_n912), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT55), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n690), .B2(new_n367), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n374), .A2(KEYINPUT95), .A3(new_n377), .ZN(new_n1195));
  AOI21_X1  g0995(.A(KEYINPUT95), .B1(new_n374), .B2(new_n377), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n367), .B(new_n1193), .C1(new_n1195), .C2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1191), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n367), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1193), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1202), .A2(new_n1190), .A3(new_n1197), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1199), .A2(new_n1203), .ZN(new_n1204));
  AND3_X1   g1004(.A1(new_n931), .A2(new_n1189), .A3(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1204), .B1(new_n931), .B2(new_n1189), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1187), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1199), .A2(new_n1203), .ZN(new_n1208));
  OAI21_X1  g1008(.A(G330), .B1(new_n944), .B2(new_n951), .ZN(new_n1209));
  AOI21_X1  g1009(.A(KEYINPUT40), .B1(new_n1185), .B2(new_n910), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1208), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n931), .A2(new_n1189), .A3(new_n1204), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1211), .A2(new_n972), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1207), .A2(new_n1213), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1142), .A2(new_n1123), .A3(new_n1127), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1216));
  OAI211_X1 g1016(.A(KEYINPUT57), .B(new_n1214), .C1(new_n1215), .C2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n1049), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1136), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1140), .B(new_n1141), .C1(new_n1147), .C2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT57), .B1(new_n1220), .B2(new_n1214), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1218), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n784), .B1(new_n1207), .B2(new_n1213), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1208), .A2(new_n791), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n850), .A2(G77), .B1(new_n851), .B2(G58), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n549), .B2(new_n822), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n280), .A2(new_n253), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n830), .A2(new_n222), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n832), .A2(new_n380), .B1(new_n827), .B2(new_n1071), .ZN(new_n1229));
  NOR4_X1   g1029(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n813), .A2(G116), .B1(G68), .B2(new_n817), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1231), .A2(KEYINPUT117), .ZN(new_n1232));
  NOR2_X1   g1032(.A1(new_n1231), .A2(KEYINPUT117), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1230), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT58), .ZN(new_n1235));
  OR2_X1    g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n830), .A2(new_n1159), .B1(new_n832), .B2(new_n874), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(G132), .B2(new_n845), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1165), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n817), .A2(G150), .B1(new_n850), .B2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1239), .B(new_n1241), .C1(new_n1164), .C2(new_n812), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1242), .A2(KEYINPUT59), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(KEYINPUT59), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n851), .A2(G159), .ZN(new_n1245));
  AOI211_X1 g1045(.A(G33), .B(G41), .C1(new_n843), .C2(G124), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1227), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1248));
  XOR2_X1   g1048(.A(new_n1248), .B(KEYINPUT116), .Z(new_n1249));
  NAND4_X1  g1049(.A1(new_n1236), .A2(new_n1237), .A3(new_n1247), .A4(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n803), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n787), .B1(new_n201), .B2(new_n870), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1224), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1223), .A2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1222), .A2(new_n1255), .ZN(G375));
  NAND2_X1  g1056(.A1(new_n1216), .A2(new_n1219), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1257), .A2(new_n1031), .A3(new_n1142), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n968), .A2(new_n791), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n786), .B1(G68), .B2(new_n1151), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n830), .A2(new_n874), .B1(new_n827), .B2(new_n1159), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n280), .B(new_n1261), .C1(G150), .C2(new_n833), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n850), .A2(G159), .B1(new_n851), .B2(G58), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(G50), .A2(new_n817), .B1(new_n845), .B2(new_n1240), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1262), .A2(new_n1263), .A3(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n812), .A2(new_n879), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n812), .A2(new_n836), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n817), .A2(new_n553), .B1(new_n851), .B2(G77), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(G116), .A2(new_n845), .B1(new_n850), .B2(G97), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n872), .A2(G283), .B1(new_n833), .B2(G107), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n333), .B1(new_n843), .B2(G303), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .A4(new_n1271), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n1265), .A2(new_n1266), .B1(new_n1267), .B2(new_n1272), .ZN(new_n1273));
  OR2_X1    g1073(.A1(new_n1273), .A2(KEYINPUT119), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n890), .B1(new_n1273), .B2(KEYINPUT119), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1260), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n1136), .A2(new_n785), .B1(new_n1259), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1258), .A2(new_n1277), .ZN(G381));
  NAND3_X1  g1078(.A1(new_n1050), .A2(new_n856), .A3(new_n1083), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(G384), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT120), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1282), .A2(G381), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n776), .B1(new_n1087), .B2(new_n1046), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n784), .B1(new_n1284), .B2(new_n1030), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1042), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1286), .A2(new_n1003), .A3(new_n1090), .A4(new_n1113), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1280), .A2(KEYINPUT120), .A3(new_n1281), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1283), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT121), .ZN(new_n1291));
  AND2_X1   g1091(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1290), .A2(new_n1291), .ZN(new_n1293));
  AND2_X1   g1093(.A1(new_n1149), .A2(new_n1174), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1222), .A2(new_n1294), .A3(new_n1255), .ZN(new_n1295));
  OR3_X1    g1095(.A1(new_n1292), .A2(new_n1293), .A3(new_n1295), .ZN(G407));
  NAND2_X1  g1096(.A1(new_n698), .A2(G213), .ZN(new_n1297));
  OAI211_X1 g1097(.A(G407), .B(G213), .C1(new_n1295), .C2(new_n1297), .ZN(G409));
  AND3_X1   g1098(.A1(new_n1211), .A2(new_n972), .A3(new_n1212), .ZN(new_n1299));
  AOI22_X1  g1099(.A1(new_n1211), .A2(new_n1212), .B1(new_n1183), .B2(new_n1186), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n785), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1301), .A2(KEYINPUT122), .A3(new_n1253), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT122), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1303), .B1(new_n1223), .B2(new_n1254), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1031), .B(new_n1214), .C1(new_n1215), .C2(new_n1216), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1302), .A2(new_n1304), .A3(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT123), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1306), .A2(new_n1307), .A3(new_n1294), .ZN(new_n1308));
  OAI211_X1 g1108(.A(G378), .B(new_n1255), .C1(new_n1218), .C2(new_n1221), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1307), .B1(new_n1306), .B2(new_n1294), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1297), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT60), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1257), .A2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1216), .A2(new_n1219), .A3(KEYINPUT60), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1314), .A2(new_n1049), .A3(new_n1142), .A4(new_n1315), .ZN(new_n1316));
  AOI21_X1  g1116(.A(G384), .B1(new_n1316), .B2(new_n1277), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1316), .A2(G384), .A3(new_n1277), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n698), .A2(G213), .A3(G2897), .ZN(new_n1320));
  AND3_X1   g1120(.A1(new_n1318), .A2(new_n1319), .A3(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1320), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1321), .A2(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(KEYINPUT61), .B1(new_n1312), .B2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1319), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1325), .A2(new_n1317), .ZN(new_n1326));
  OAI211_X1 g1126(.A(new_n1326), .B(new_n1297), .C1(new_n1310), .C2(new_n1311), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1311), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1330), .A2(new_n1309), .A3(new_n1308), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT62), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1331), .A2(new_n1332), .A3(new_n1297), .A4(new_n1326), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1324), .A2(new_n1329), .A3(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(G387), .A2(G390), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT125), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1335), .A2(new_n1287), .A3(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n856), .B1(new_n1050), .B2(new_n1083), .ZN(new_n1338));
  OAI21_X1  g1138(.A(KEYINPUT124), .B1(new_n1280), .B2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(G393), .A2(G396), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT124), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1340), .A2(new_n1341), .A3(new_n1279), .ZN(new_n1342));
  AND2_X1   g1142(.A1(new_n1339), .A2(new_n1342), .ZN(new_n1343));
  AND3_X1   g1143(.A1(new_n1337), .A2(new_n1343), .A3(KEYINPUT126), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1337), .A2(KEYINPUT126), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT126), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1335), .A2(new_n1287), .A3(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1339), .A2(new_n1342), .ZN(new_n1348));
  AND2_X1   g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n1344), .B1(new_n1345), .B2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1334), .A2(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT63), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1327), .A2(new_n1353), .ZN(new_n1354));
  NAND4_X1  g1154(.A1(new_n1331), .A2(KEYINPUT63), .A3(new_n1297), .A4(new_n1326), .ZN(new_n1355));
  NAND4_X1  g1155(.A1(new_n1350), .A2(new_n1324), .A3(new_n1354), .A4(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1352), .A2(new_n1356), .ZN(G405));
  NAND2_X1  g1157(.A1(G375), .A2(G378), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1358), .A2(new_n1295), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1359), .A2(new_n1326), .ZN(new_n1360));
  OAI211_X1 g1160(.A(new_n1358), .B(new_n1295), .C1(new_n1317), .C2(new_n1325), .ZN(new_n1361));
  AND3_X1   g1161(.A1(new_n1350), .A2(new_n1360), .A3(new_n1361), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1350), .B1(new_n1360), .B2(new_n1361), .ZN(new_n1363));
  NOR2_X1   g1163(.A1(new_n1362), .A2(new_n1363), .ZN(G402));
endmodule


