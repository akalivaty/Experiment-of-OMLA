//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1278, new_n1279,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  INV_X1    g0012(.A(new_n201), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n207), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n212), .B(new_n218), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XNOR2_X1  g0039(.A(G68), .B(G77), .ZN(new_n240));
  INV_X1    g0040(.A(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(KEYINPUT65), .B(G50), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G97), .B(G107), .Z(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  INV_X1    g0048(.A(KEYINPUT10), .ZN(new_n249));
  XOR2_X1   g0049(.A(KEYINPUT8), .B(G58), .Z(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G20), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n207), .A2(new_n251), .A3(KEYINPUT68), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT68), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n255), .B1(G20), .B2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G150), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT69), .ZN(new_n259));
  NOR3_X1   g0059(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n259), .B1(new_n260), .B2(new_n207), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n203), .A2(KEYINPUT69), .A3(G20), .ZN(new_n262));
  NAND4_X1  g0062(.A1(new_n253), .A2(new_n258), .A3(new_n261), .A4(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n216), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n263), .A2(new_n265), .B1(new_n202), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT73), .ZN(new_n269));
  INV_X1    g0069(.A(new_n265), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n266), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT70), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n270), .A2(KEYINPUT70), .A3(new_n266), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n206), .A2(G20), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n273), .A2(new_n274), .A3(G50), .A4(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n268), .A2(new_n269), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n269), .B1(new_n268), .B2(new_n276), .ZN(new_n279));
  OAI21_X1  g0079(.A(KEYINPUT9), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n279), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT9), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(new_n282), .A3(new_n277), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G190), .ZN(new_n285));
  INV_X1    g0085(.A(G200), .ZN(new_n286));
  OR2_X1    g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  AOI21_X1  g0088(.A(G1698), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G222), .ZN(new_n290));
  INV_X1    g0090(.A(G77), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT3), .B(G33), .ZN(new_n292));
  INV_X1    g0092(.A(G223), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(G1698), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n290), .B1(new_n291), .B2(new_n292), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  AND2_X1   g0095(.A1(G1), .A2(G13), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G41), .ZN(new_n297));
  AND3_X1   g0097(.A1(new_n296), .A2(KEYINPUT67), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(KEYINPUT67), .B1(new_n296), .B2(new_n297), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n295), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G274), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n302), .B1(new_n296), .B2(new_n297), .ZN(new_n303));
  NOR2_X1   g0103(.A1(G41), .A2(G45), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(G1), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT66), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(new_n304), .B2(G1), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n296), .A2(new_n297), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n206), .B(KEYINPUT66), .C1(G41), .C2(G45), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n307), .B1(new_n312), .B2(G226), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n301), .A2(new_n313), .ZN(new_n314));
  MUX2_X1   g0114(.A(new_n285), .B(new_n286), .S(new_n314), .Z(new_n315));
  AOI21_X1  g0115(.A(new_n249), .B1(new_n284), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n284), .A2(new_n249), .A3(new_n315), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G169), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n314), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n268), .A2(new_n276), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n321), .B(new_n322), .C1(G179), .C2(new_n314), .ZN(new_n323));
  XOR2_X1   g0123(.A(new_n323), .B(KEYINPUT71), .Z(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT15), .B(G87), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  AOI22_X1  g0127(.A1(new_n327), .A2(new_n252), .B1(G20), .B2(G77), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n250), .A2(new_n257), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n270), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n275), .A2(G77), .ZN(new_n331));
  OAI22_X1  g0131(.A1(new_n271), .A2(new_n331), .B1(G77), .B2(new_n266), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G1698), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n292), .A2(G232), .A3(new_n334), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT72), .B(G107), .ZN(new_n336));
  OAI221_X1 g0136(.A(new_n335), .B1(new_n292), .B2(new_n336), .C1(new_n294), .C2(new_n221), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n300), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n307), .B1(new_n312), .B2(G244), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n333), .B1(G200), .B2(new_n340), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n338), .A2(new_n339), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G190), .ZN(new_n343));
  INV_X1    g0143(.A(G179), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n330), .A2(new_n332), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(new_n340), .B2(new_n320), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n341), .A2(new_n343), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n319), .A2(new_n325), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n267), .A2(new_n220), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT12), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n275), .A2(G68), .ZN(new_n352));
  INV_X1    g0152(.A(new_n257), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(new_n202), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n207), .A2(G33), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n355), .A2(new_n291), .B1(new_n207), .B2(G68), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n265), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT11), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n351), .B1(new_n271), .B2(new_n352), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n357), .A2(new_n358), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT14), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n309), .A2(G238), .A3(new_n310), .A4(new_n311), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n306), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT75), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n364), .A2(KEYINPUT75), .A3(new_n306), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G232), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(G1698), .ZN(new_n371));
  AND2_X1   g0171(.A1(KEYINPUT3), .A2(G33), .ZN(new_n372));
  NOR2_X1   g0172(.A1(KEYINPUT3), .A2(G33), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n371), .B1(G226), .B2(G1698), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G33), .A2(G97), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT74), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n374), .A2(KEYINPUT74), .A3(new_n375), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n379), .A3(new_n300), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT13), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n369), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n381), .B1(new_n369), .B2(new_n380), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n363), .B(G169), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n369), .A2(new_n380), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(KEYINPUT13), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n387), .A2(G179), .A3(new_n382), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n382), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n363), .B1(new_n390), .B2(G169), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n362), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(G200), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n393), .B(new_n361), .C1(new_n285), .C2(new_n390), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT16), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n292), .B2(G20), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n372), .A2(new_n373), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n399), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n220), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g0201(.A(G58), .B(G68), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G20), .ZN(new_n403));
  INV_X1    g0203(.A(G159), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n403), .B1(new_n353), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n396), .B1(new_n401), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT7), .B1(new_n399), .B2(new_n207), .ZN(new_n407));
  NOR4_X1   g0207(.A1(new_n372), .A2(new_n373), .A3(new_n397), .A4(G20), .ZN(new_n408));
  OAI21_X1  g0208(.A(G68), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n257), .A2(G159), .B1(new_n402), .B2(G20), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n409), .A2(KEYINPUT16), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n406), .A2(new_n411), .A3(new_n265), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT76), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n406), .A2(new_n411), .A3(KEYINPUT76), .A4(new_n265), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n250), .A2(new_n267), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n273), .A2(new_n275), .A3(new_n274), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n417), .B1(new_n418), .B2(new_n250), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT18), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n309), .A2(G232), .A3(new_n310), .A4(new_n311), .ZN(new_n423));
  OR2_X1    g0223(.A1(new_n298), .A2(new_n299), .ZN(new_n424));
  MUX2_X1   g0224(.A(G223), .B(G226), .S(G1698), .Z(new_n425));
  AOI22_X1  g0225(.A1(new_n425), .A2(new_n292), .B1(G33), .B2(G87), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n306), .B(new_n423), .C1(new_n424), .C2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n427), .A2(new_n344), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n428), .B1(G169), .B2(new_n427), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n421), .A2(new_n422), .A3(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n427), .A2(new_n285), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(G200), .B2(new_n427), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n416), .A2(new_n420), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT17), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n419), .B1(new_n414), .B2(new_n415), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT18), .B1(new_n437), .B2(new_n429), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(KEYINPUT17), .A3(new_n433), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n431), .A2(new_n436), .A3(new_n438), .A4(new_n439), .ZN(new_n440));
  NOR3_X1   g0240(.A1(new_n349), .A2(new_n395), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT81), .ZN(new_n442));
  INV_X1    g0242(.A(G41), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n206), .B(G45), .C1(new_n443), .C2(KEYINPUT5), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT77), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT5), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G41), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT77), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(new_n206), .A4(G45), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n446), .A2(G41), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n445), .A2(new_n449), .A3(new_n303), .A4(new_n451), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n310), .B(G270), .C1(new_n444), .C2(new_n450), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(G264), .B(G1698), .C1(new_n372), .C2(new_n373), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT80), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n292), .A2(KEYINPUT80), .A3(G264), .A4(G1698), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n399), .A2(G303), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n292), .A2(G257), .A3(new_n334), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n457), .A2(new_n458), .A3(new_n459), .A4(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n454), .B1(new_n300), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(G116), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n264), .A2(new_n216), .B1(G20), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  INV_X1    g0265(.A(G97), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n465), .B(new_n207), .C1(G33), .C2(new_n466), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n464), .A2(KEYINPUT20), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(KEYINPUT20), .B1(new_n464), .B2(new_n467), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n267), .A2(G116), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n206), .A2(G33), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n266), .A2(new_n472), .A3(new_n216), .A4(new_n264), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n471), .B1(G116), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(G169), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n462), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n442), .B1(new_n476), .B2(KEYINPUT21), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n461), .A2(new_n300), .ZN(new_n478));
  INV_X1    g0278(.A(new_n454), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n464), .A2(new_n467), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT20), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n464), .A2(KEYINPUT20), .A3(new_n467), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n473), .A2(G116), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(G116), .B2(new_n267), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n320), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n480), .A2(new_n442), .A3(KEYINPUT21), .A4(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n485), .A2(new_n487), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n462), .A2(G179), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(KEYINPUT82), .B1(new_n477), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n480), .A2(KEYINPUT21), .A3(new_n488), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT81), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT82), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n495), .A2(new_n496), .A3(new_n491), .A4(new_n489), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT21), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n462), .B2(new_n475), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n490), .B1(new_n480), .B2(G200), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n462), .A2(G190), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n493), .A2(new_n497), .A3(new_n499), .A4(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(G13), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(G1), .ZN(new_n506));
  INV_X1    g0306(.A(G107), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n506), .A2(G20), .A3(new_n507), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n508), .B(KEYINPUT25), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n473), .A2(new_n507), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT22), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT83), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n207), .B1(new_n372), .B2(new_n373), .ZN(new_n514));
  OAI21_X1  g0314(.A(G87), .B1(new_n512), .B2(KEYINPUT83), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT83), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n222), .B1(new_n517), .B2(KEYINPUT22), .ZN(new_n518));
  INV_X1    g0318(.A(new_n513), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n292), .A2(new_n518), .A3(new_n519), .A4(new_n207), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT23), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n522), .A2(new_n507), .A3(G20), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n463), .B2(new_n355), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n507), .A2(KEYINPUT72), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT72), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G107), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n527), .A3(G20), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n524), .B1(KEYINPUT23), .B2(new_n528), .ZN(new_n529));
  AND3_X1   g0329(.A1(new_n521), .A2(KEYINPUT84), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT84), .B1(new_n521), .B2(new_n529), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT24), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(G20), .B1(new_n287), .B2(new_n288), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n519), .B1(new_n534), .B2(new_n518), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n514), .A2(new_n515), .A3(new_n513), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n529), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT84), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n538), .A3(new_n532), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n265), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n511), .B1(new_n533), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(G257), .B(G1698), .C1(new_n372), .C2(new_n373), .ZN(new_n542));
  OAI211_X1 g0342(.A(G250), .B(new_n334), .C1(new_n372), .C2(new_n373), .ZN(new_n543));
  AND2_X1   g0343(.A1(KEYINPUT85), .A2(G294), .ZN(new_n544));
  NOR2_X1   g0344(.A1(KEYINPUT85), .A2(G294), .ZN(new_n545));
  OAI21_X1  g0345(.A(G33), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n542), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n300), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n310), .B(G264), .C1(new_n444), .C2(new_n450), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(new_n452), .A3(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n550), .A2(G179), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n320), .B2(new_n550), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n541), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n537), .A2(new_n538), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n521), .A2(KEYINPUT84), .A3(new_n529), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(KEYINPUT24), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n270), .B1(new_n531), .B2(new_n532), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT86), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n548), .A2(G190), .A3(new_n452), .A4(new_n549), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n511), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n452), .A2(new_n549), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n286), .B1(new_n562), .B2(new_n548), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AND3_X1   g0364(.A1(new_n558), .A2(new_n559), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n559), .B1(new_n558), .B2(new_n564), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n553), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT87), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT87), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n569), .B(new_n553), .C1(new_n565), .C2(new_n566), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n252), .A2(G97), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT19), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n220), .B2(new_n514), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n525), .A2(new_n527), .A3(new_n466), .ZN(new_n576));
  XNOR2_X1  g0376(.A(KEYINPUT78), .B(G87), .ZN(new_n577));
  NAND3_X1  g0377(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n576), .A2(new_n577), .B1(new_n207), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n265), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  OR2_X1    g0380(.A1(new_n473), .A2(new_n222), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n327), .A2(new_n266), .ZN(new_n582));
  INV_X1    g0382(.A(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n206), .A2(new_n302), .A3(G45), .ZN(new_n585));
  INV_X1    g0385(.A(G45), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n223), .B1(new_n586), .B2(G1), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n310), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(G244), .B(G1698), .C1(new_n372), .C2(new_n373), .ZN(new_n590));
  OAI211_X1 g0390(.A(G238), .B(new_n334), .C1(new_n372), .C2(new_n373), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n590), .B(new_n591), .C1(new_n251), .C2(new_n463), .ZN(new_n592));
  AOI211_X1 g0392(.A(new_n285), .B(new_n589), .C1(new_n592), .C2(new_n300), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n584), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n589), .B1(new_n592), .B2(new_n300), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n595), .A2(new_n286), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n595), .A2(G169), .ZN(new_n598));
  AOI211_X1 g0398(.A(G179), .B(new_n589), .C1(new_n592), .C2(new_n300), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n580), .B(new_n583), .C1(new_n326), .C2(new_n473), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n594), .A2(new_n597), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(G250), .B(G1698), .C1(new_n372), .C2(new_n373), .ZN(new_n603));
  OAI211_X1 g0403(.A(G244), .B(new_n334), .C1(new_n372), .C2(new_n373), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT4), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n465), .B(new_n603), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT4), .B1(new_n289), .B2(G244), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n300), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n310), .B(G257), .C1(new_n444), .C2(new_n450), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n608), .A2(new_n452), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n320), .ZN(new_n611));
  INV_X1    g0411(.A(new_n609), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n604), .A2(new_n605), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n292), .A2(KEYINPUT4), .A3(G244), .A4(new_n334), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n613), .A2(new_n614), .A3(new_n465), .A4(new_n603), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n612), .B1(new_n615), .B2(new_n300), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n616), .A2(new_n344), .A3(new_n452), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT6), .ZN(new_n618));
  NOR3_X1   g0418(.A1(new_n618), .A2(new_n466), .A3(G107), .ZN(new_n619));
  XNOR2_X1  g0419(.A(G97), .B(G107), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n619), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  OAI22_X1  g0421(.A1(new_n621), .A2(new_n207), .B1(new_n291), .B2(new_n353), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n336), .B1(new_n398), .B2(new_n400), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n265), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  MUX2_X1   g0424(.A(new_n266), .B(new_n473), .S(G97), .Z(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n611), .A2(new_n617), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n610), .A2(G200), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n616), .A2(G190), .A3(new_n452), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n628), .A2(new_n629), .A3(new_n624), .A4(new_n625), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n602), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT79), .ZN(new_n632));
  XNOR2_X1  g0432(.A(new_n631), .B(new_n632), .ZN(new_n633));
  AND4_X1   g0433(.A1(new_n441), .A2(new_n504), .A3(new_n571), .A4(new_n633), .ZN(G372));
  NAND2_X1  g0434(.A1(new_n595), .A2(new_n344), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(G169), .B2(new_n595), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n336), .A2(new_n577), .A3(new_n466), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n578), .A2(new_n207), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n534), .A2(G68), .B1(new_n572), .B2(new_n573), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n270), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n473), .A2(new_n326), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n641), .A2(new_n582), .A3(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n636), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n627), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n602), .A2(new_n645), .A3(KEYINPUT26), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n595), .A2(G190), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n648), .A2(new_n580), .A3(new_n583), .A4(new_n581), .ZN(new_n649));
  OAI22_X1  g0449(.A1(new_n649), .A2(new_n596), .B1(new_n636), .B2(new_n643), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n647), .B1(new_n650), .B2(new_n627), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n644), .B1(new_n646), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n558), .A2(new_n564), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(KEYINPUT86), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n558), .A2(new_n559), .A3(new_n564), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n630), .A2(new_n627), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n657), .A2(new_n650), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n553), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n495), .A2(new_n499), .A3(new_n491), .A4(new_n489), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n652), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n441), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n436), .A2(new_n439), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n394), .A2(new_n345), .A3(new_n347), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n665), .B1(new_n666), .B2(new_n392), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n431), .A2(new_n438), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n319), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n669), .A2(new_n325), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n664), .A2(new_n670), .ZN(G369));
  INV_X1    g0471(.A(KEYINPUT88), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n503), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n499), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n495), .A2(new_n491), .A3(new_n489), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n674), .B1(new_n675), .B2(KEYINPUT82), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n676), .A2(KEYINPUT88), .A3(new_n497), .A4(new_n502), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n506), .A2(new_n207), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G213), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n490), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n673), .A2(new_n677), .A3(new_n684), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n661), .A2(new_n684), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n685), .A2(G330), .A3(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n541), .A2(new_n683), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n569), .B1(new_n656), .B2(new_n553), .ZN(new_n690));
  INV_X1    g0490(.A(new_n570), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n683), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n553), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n688), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n553), .A2(new_n683), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n683), .B1(new_n676), .B2(new_n497), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n698), .B1(new_n571), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n697), .A2(new_n700), .ZN(G399));
  INV_X1    g0501(.A(KEYINPUT91), .ZN(new_n702));
  AOI21_X1  g0502(.A(G179), .B1(new_n562), .B2(new_n548), .ZN(new_n703));
  INV_X1    g0503(.A(new_n595), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n480), .A2(new_n703), .A3(new_n610), .A4(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT90), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n704), .A2(new_n550), .A3(new_n344), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n708), .A2(KEYINPUT90), .A3(new_n480), .A4(new_n610), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n616), .A2(new_n548), .A3(new_n562), .A4(new_n595), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n462), .A2(G179), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n478), .A2(G179), .A3(new_n479), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n704), .A2(new_n550), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n714), .A2(new_n715), .A3(KEYINPUT30), .A4(new_n616), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n707), .A2(new_n709), .A3(new_n713), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(new_n683), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT31), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n713), .A2(new_n716), .A3(new_n705), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n702), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(KEYINPUT31), .B1(new_n717), .B2(new_n683), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n683), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n724), .A2(new_n725), .A3(KEYINPUT91), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n571), .A2(new_n633), .A3(new_n504), .A4(new_n693), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(G330), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n663), .A2(new_n693), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT29), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n731), .A2(KEYINPUT92), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT92), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n656), .B(new_n658), .C1(new_n660), .C2(new_n661), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n683), .B1(new_n735), .B2(new_n652), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n734), .B1(new_n736), .B2(KEYINPUT29), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n493), .A2(new_n497), .A3(new_n499), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n656), .B(new_n658), .C1(new_n738), .C2(new_n660), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n652), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n740), .A2(KEYINPUT29), .A3(new_n693), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n733), .A2(new_n737), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n730), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n206), .ZN(new_n744));
  INV_X1    g0544(.A(new_n210), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G41), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G1), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n576), .A2(new_n463), .A3(new_n577), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n748), .A2(new_n749), .B1(new_n214), .B2(new_n747), .ZN(new_n750));
  XOR2_X1   g0550(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n751));
  XNOR2_X1  g0551(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n744), .A2(new_n752), .ZN(G364));
  NOR2_X1   g0553(.A1(new_n505), .A2(G20), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G45), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G1), .ZN(new_n756));
  OR3_X1    g0556(.A1(new_n746), .A2(KEYINPUT93), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(KEYINPUT93), .B1(new_n746), .B2(new_n756), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n745), .A2(new_n399), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT94), .ZN(new_n762));
  NAND2_X1  g0562(.A1(G355), .A2(new_n762), .ZN(new_n763));
  OR2_X1    g0563(.A1(G355), .A2(new_n762), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n761), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n765), .B1(G116), .B2(new_n210), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n244), .A2(G45), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n745), .A2(new_n292), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(new_n586), .B2(new_n215), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n766), .B1(new_n767), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G13), .A2(G33), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n216), .B1(G20), .B2(new_n320), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n760), .B1(new_n771), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n286), .A2(G179), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT97), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n207), .A2(new_n285), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT99), .Z(new_n783));
  NAND3_X1  g0583(.A1(new_n781), .A2(G179), .A3(new_n286), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(KEYINPUT95), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n784), .A2(KEYINPUT95), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G322), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n207), .A2(new_n344), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G200), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G190), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  XOR2_X1   g0593(.A(KEYINPUT33), .B(G317), .Z(new_n794));
  OAI22_X1  g0594(.A1(new_n788), .A2(new_n789), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n783), .A2(G303), .B1(new_n795), .B2(KEYINPUT101), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(KEYINPUT101), .B2(new_n795), .ZN(new_n797));
  NOR2_X1   g0597(.A1(G179), .A2(G200), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n207), .B1(new_n798), .B2(G190), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n544), .A2(new_n545), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n790), .A2(new_n285), .A3(new_n286), .ZN(new_n802));
  INV_X1    g0602(.A(G311), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n399), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n791), .A2(new_n285), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n801), .B(new_n804), .C1(G326), .C2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G283), .ZN(new_n807));
  OAI21_X1  g0607(.A(KEYINPUT96), .B1(new_n207), .B2(G190), .ZN(new_n808));
  OR3_X1    g0608(.A1(new_n207), .A2(KEYINPUT96), .A3(G190), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n780), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n809), .A2(new_n798), .A3(new_n808), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n812), .A2(KEYINPUT100), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(KEYINPUT100), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G329), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n806), .B1(new_n807), .B2(new_n810), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n292), .B1(new_n782), .B2(new_n577), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT98), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n812), .A2(G159), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT32), .Z(new_n821));
  INV_X1    g0621(.A(new_n802), .ZN(new_n822));
  INV_X1    g0622(.A(new_n799), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n822), .A2(G77), .B1(new_n823), .B2(G97), .ZN(new_n824));
  INV_X1    g0624(.A(new_n788), .ZN(new_n825));
  INV_X1    g0625(.A(new_n810), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n825), .A2(G58), .B1(G107), .B2(new_n826), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n792), .A2(G68), .B1(new_n805), .B2(G50), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n821), .A2(new_n824), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n797), .A2(new_n817), .B1(new_n819), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n778), .B1(new_n830), .B2(new_n775), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n685), .A2(new_n686), .ZN(new_n832));
  INV_X1    g0632(.A(new_n774), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n832), .A2(G330), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n687), .A2(new_n759), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g0637(.A(new_n837), .B(KEYINPUT102), .ZN(G396));
  INV_X1    g0638(.A(G294), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n788), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g0640(.A(KEYINPUT103), .B(G283), .Z(new_n841));
  INV_X1    g0641(.A(new_n805), .ZN(new_n842));
  INV_X1    g0642(.A(G303), .ZN(new_n843));
  OAI22_X1  g0643(.A1(new_n793), .A2(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n810), .A2(new_n222), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n399), .B1(new_n799), .B2(new_n466), .C1(new_n802), .C2(new_n463), .ZN(new_n846));
  NOR4_X1   g0646(.A1(new_n840), .A2(new_n844), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n783), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n847), .B1(new_n803), .B2(new_n815), .C1(new_n507), .C2(new_n848), .ZN(new_n849));
  AOI22_X1  g0649(.A1(G137), .A2(new_n805), .B1(new_n822), .B2(G159), .ZN(new_n850));
  INV_X1    g0650(.A(G150), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n850), .B1(new_n851), .B2(new_n793), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(G143), .B2(new_n825), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT34), .ZN(new_n854));
  INV_X1    g0654(.A(new_n815), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(G132), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n292), .B1(new_n799), .B2(new_n241), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(new_n826), .B2(G68), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n856), .B(new_n858), .C1(new_n848), .C2(new_n202), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n849), .B1(new_n854), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n775), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n775), .A2(new_n772), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n759), .B1(new_n291), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n345), .A2(new_n347), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT104), .B1(new_n864), .B2(new_n693), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT104), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n345), .A2(new_n347), .A3(new_n866), .A4(new_n683), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n333), .A2(new_n683), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n865), .A2(new_n867), .B1(new_n348), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n861), .B(new_n863), .C1(new_n870), .C2(new_n773), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n736), .A2(new_n870), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n683), .B(new_n869), .C1(new_n735), .C2(new_n652), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n760), .B1(new_n875), .B2(new_n730), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n875), .A2(new_n730), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n871), .B1(new_n877), .B2(new_n878), .ZN(G384));
  NOR2_X1   g0679(.A1(new_n754), .A2(new_n206), .ZN(new_n880));
  INV_X1    g0680(.A(G330), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n409), .A2(new_n410), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT16), .B1(new_n882), .B2(KEYINPUT106), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(KEYINPUT106), .B2(new_n882), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(new_n265), .A3(new_n411), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n681), .B1(new_n885), .B2(new_n420), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n440), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n421), .A2(new_n430), .ZN(new_n888));
  INV_X1    g0688(.A(new_n681), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n421), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT37), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n888), .A2(new_n890), .A3(new_n891), .A4(new_n434), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n885), .A2(new_n420), .B1(new_n429), .B2(new_n681), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n416), .A2(new_n420), .A3(new_n433), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT37), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n887), .A2(KEYINPUT38), .A3(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n434), .B1(new_n437), .B2(new_n429), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n437), .A2(new_n681), .ZN(new_n899));
  OAI21_X1  g0699(.A(KEYINPUT37), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n892), .A2(new_n900), .B1(new_n440), .B2(new_n899), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n897), .B1(new_n901), .B2(KEYINPUT38), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n392), .A2(KEYINPUT105), .A3(new_n394), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n362), .A2(new_n683), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT105), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n392), .A2(new_n906), .A3(new_n394), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n389), .A2(new_n904), .A3(new_n391), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n905), .A2(new_n909), .A3(new_n870), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n718), .A2(new_n719), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n911), .A2(new_n724), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n728), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n902), .A2(new_n910), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n905), .A2(new_n909), .A3(new_n870), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n728), .B2(new_n912), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n887), .A2(new_n896), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT38), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT40), .B1(new_n919), .B2(new_n897), .ZN(new_n920));
  AOI22_X1  g0720(.A1(KEYINPUT40), .A2(new_n914), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  AND2_X1   g0722(.A1(new_n441), .A2(new_n913), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n881), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n924), .B1(new_n923), .B2(new_n922), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n864), .A2(new_n683), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n736), .B2(new_n870), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n905), .A2(new_n909), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n919), .A2(new_n897), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n929), .A2(new_n930), .B1(new_n668), .B2(new_n681), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT39), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n902), .A2(new_n932), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n392), .A2(new_n683), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n919), .A2(KEYINPUT39), .A3(new_n897), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n933), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n931), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n441), .A2(new_n741), .A3(new_n733), .A4(new_n737), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n939), .A2(new_n670), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n938), .B(new_n940), .Z(new_n941));
  AOI21_X1  g0741(.A(new_n880), .B1(new_n925), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n941), .B2(new_n925), .ZN(new_n943));
  INV_X1    g0743(.A(new_n621), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n944), .A2(KEYINPUT35), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(KEYINPUT35), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n945), .A2(G116), .A3(new_n217), .A4(new_n946), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT36), .ZN(new_n948));
  OAI21_X1  g0748(.A(G77), .B1(new_n241), .B2(new_n220), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n214), .A2(new_n949), .B1(G50), .B2(new_n220), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n950), .A2(G1), .A3(new_n505), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n943), .A2(new_n948), .A3(new_n951), .ZN(G367));
  AOI21_X1  g0752(.A(new_n777), .B1(new_n745), .B2(new_n327), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n768), .A2(new_n238), .ZN(new_n954));
  AND2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n799), .A2(new_n220), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n292), .B1(new_n202), .B2(new_n802), .C1(new_n793), .C2(new_n404), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n956), .B(new_n957), .C1(G143), .C2(new_n805), .ZN(new_n958));
  INV_X1    g0758(.A(new_n782), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n959), .A2(G58), .B1(G137), .B2(new_n812), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n826), .A2(G77), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n825), .A2(G150), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n958), .A2(new_n960), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n783), .A2(KEYINPUT46), .A3(G116), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n399), .B1(new_n802), .B2(new_n841), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n793), .A2(new_n800), .B1(new_n336), .B2(new_n799), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n965), .B(new_n966), .C1(G311), .C2(new_n805), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n826), .A2(G97), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n825), .A2(G303), .B1(new_n812), .B2(G317), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n964), .A2(new_n967), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT46), .B1(new_n959), .B2(G116), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT111), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n963), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n973), .B(new_n974), .Z(new_n975));
  AOI211_X1 g0775(.A(new_n759), .B(new_n955), .C1(new_n975), .C2(new_n775), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n976), .A2(KEYINPUT113), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(KEYINPUT113), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n584), .A2(new_n683), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n602), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n644), .A2(new_n584), .A3(new_n683), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n977), .B(new_n978), .C1(new_n833), .C2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT109), .ZN(new_n985));
  INV_X1    g0785(.A(new_n699), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n692), .A2(new_n695), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n699), .B1(new_n690), .B2(new_n691), .ZN(new_n988));
  AND3_X1   g0788(.A1(new_n987), .A2(new_n687), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n687), .B1(new_n988), .B2(new_n987), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(KEYINPUT108), .B1(new_n991), .B2(new_n743), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n987), .A2(new_n988), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n688), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n987), .A2(new_n687), .A3(new_n988), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT108), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n996), .A2(new_n997), .A3(new_n730), .A4(new_n742), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n992), .A2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n697), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n645), .A2(new_n683), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n626), .A2(new_n683), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n630), .A2(new_n627), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(KEYINPUT45), .B1(new_n700), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n698), .ZN(new_n1006));
  AND4_X1   g0806(.A1(KEYINPUT45), .A2(new_n988), .A3(new_n1006), .A4(new_n1004), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n988), .A2(new_n1006), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1004), .ZN(new_n1010));
  XOR2_X1   g0810(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n1011));
  NAND3_X1  g0811(.A1(new_n1009), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n1011), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n700), .B2(new_n1004), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1000), .B1(new_n1008), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT45), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n700), .A2(KEYINPUT45), .A3(new_n1004), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1020), .A2(new_n697), .A3(new_n1012), .A4(new_n1014), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1016), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n743), .B1(new_n999), .B2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n746), .B(KEYINPUT41), .Z(new_n1024));
  OAI21_X1  g0824(.A(new_n985), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1024), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1016), .A2(new_n1021), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n992), .B2(new_n998), .ZN(new_n1028));
  OAI211_X1 g0828(.A(KEYINPUT109), .B(new_n1026), .C1(new_n1028), .C2(new_n743), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n756), .B(KEYINPUT110), .Z(new_n1030));
  NAND3_X1  g0830(.A1(new_n1025), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n571), .A2(new_n699), .A3(new_n1004), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1032), .A2(KEYINPUT42), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n627), .B1(new_n1003), .B2(new_n553), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n1032), .A2(KEYINPUT42), .B1(new_n693), .B2(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1033), .A2(new_n1035), .B1(KEYINPUT43), .B2(new_n982), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1036), .B(new_n1037), .Z(new_n1038));
  NOR2_X1   g0838(.A1(new_n697), .A2(new_n1010), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1038), .B(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n984), .B1(new_n1031), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(G387));
  OR2_X1    g0842(.A1(new_n235), .A2(new_n586), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1043), .A2(new_n768), .B1(new_n749), .B2(new_n761), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n250), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1045), .A2(G50), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT50), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n586), .B1(new_n220), .B2(new_n291), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n749), .B(new_n1048), .C1(new_n1047), .C2(new_n1046), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n1044), .A2(new_n1049), .B1(G107), .B2(new_n210), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n759), .B1(new_n1050), .B2(new_n776), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n782), .A2(new_n291), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n825), .B2(G50), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1053), .B(new_n968), .C1(new_n851), .C2(new_n811), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n292), .B1(new_n220), .B2(new_n802), .C1(new_n842), .C2(new_n404), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n793), .A2(new_n1045), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n799), .A2(new_n326), .ZN(new_n1057));
  NOR4_X1   g0857(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G311), .A2(new_n792), .B1(new_n822), .B2(G303), .ZN(new_n1059));
  INV_X1    g0859(.A(G317), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1059), .B1(new_n789), .B2(new_n842), .C1(new_n788), .C2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT48), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n782), .A2(new_n800), .B1(new_n799), .B2(new_n841), .ZN(new_n1065));
  OR3_X1    g0865(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1067), .A2(KEYINPUT49), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n292), .B1(new_n812), .B2(G326), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n463), .B2(new_n810), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT114), .Z(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(new_n1067), .B2(KEYINPUT49), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1058), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n775), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1051), .B1(new_n1073), .B2(new_n1074), .C1(new_n696), .C2(new_n833), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n991), .A2(new_n743), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n746), .B1(new_n991), .B2(new_n743), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1075), .B1(new_n991), .B2(new_n1030), .C1(new_n1076), .C2(new_n1077), .ZN(G393));
  NOR2_X1   g0878(.A1(new_n1028), .A2(new_n747), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n991), .A2(new_n743), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT115), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1021), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(KEYINPUT115), .B2(new_n1027), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1079), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1030), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1010), .A2(new_n774), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n782), .A2(new_n841), .B1(new_n789), .B2(new_n811), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n292), .B(new_n1087), .C1(G107), .C2(new_n826), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1088), .B(KEYINPUT117), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n788), .A2(new_n803), .B1(new_n1060), .B2(new_n842), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT52), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n792), .A2(G303), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n822), .A2(G294), .B1(new_n823), .B2(G116), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1089), .A2(new_n1091), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n788), .A2(new_n404), .B1(new_n851), .B2(new_n842), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1095), .B(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n799), .A2(new_n291), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n292), .B1(new_n1045), .B2(new_n802), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1098), .B(new_n1099), .C1(G50), .C2(new_n792), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n782), .A2(new_n220), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1101), .B(new_n845), .C1(G143), .C2(new_n812), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1097), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1074), .B1(new_n1094), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n769), .A2(new_n247), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n777), .B(new_n1105), .C1(G97), .C2(new_n745), .ZN(new_n1106));
  NOR3_X1   g0906(.A1(new_n1104), .A2(new_n759), .A3(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1083), .A2(new_n1085), .B1(new_n1086), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1084), .A2(new_n1108), .ZN(G390));
  NAND3_X1  g0909(.A1(new_n441), .A2(G330), .A3(new_n913), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n939), .A2(new_n670), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n927), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n904), .A2(new_n903), .B1(new_n907), .B2(new_n908), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n881), .B1(new_n727), .B2(new_n728), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1113), .B1(new_n1114), .B2(new_n870), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n913), .A2(G330), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1116), .A2(new_n915), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1112), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n928), .B1(new_n1116), .B2(new_n869), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n683), .B1(new_n739), .B2(new_n652), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n926), .B1(new_n1120), .B2(new_n870), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1114), .A2(new_n870), .A3(new_n1113), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1119), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1111), .B1(new_n1118), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1113), .B1(new_n873), .B2(new_n926), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n933), .A2(new_n936), .B1(new_n934), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n902), .A2(new_n934), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n740), .A2(new_n693), .A3(new_n870), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n926), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n928), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1117), .B1(new_n1127), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n900), .A2(new_n892), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n440), .A2(new_n899), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n918), .ZN(new_n1137));
  AOI21_X1  g0937(.A(KEYINPUT39), .B1(new_n1137), .B2(new_n897), .ZN(new_n1138));
  AND3_X1   g0938(.A1(new_n887), .A2(KEYINPUT38), .A3(new_n896), .ZN(new_n1139));
  AOI21_X1  g0939(.A(KEYINPUT38), .B1(new_n887), .B2(new_n896), .ZN(new_n1140));
  NOR3_X1   g0940(.A1(new_n1139), .A2(new_n1140), .A3(new_n932), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n1138), .A2(new_n1141), .B1(new_n929), .B2(new_n935), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n934), .B(new_n902), .C1(new_n1121), .C2(new_n928), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n1143), .A3(new_n1122), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1133), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1125), .A2(new_n1145), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n1133), .A2(new_n1144), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1147), .A2(new_n1124), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1146), .A2(new_n1148), .A3(new_n746), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n772), .B1(new_n1138), .B2(new_n1141), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n788), .A2(new_n463), .B1(new_n810), .B2(new_n220), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n807), .A2(new_n842), .B1(new_n793), .B2(new_n336), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n399), .B1(new_n802), .B2(new_n466), .ZN(new_n1153));
  NOR4_X1   g0953(.A1(new_n1151), .A2(new_n1098), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  OAI221_X1 g0954(.A(new_n1154), .B1(new_n839), .B2(new_n815), .C1(new_n222), .C2(new_n848), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(KEYINPUT54), .B(G143), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n292), .B1(new_n802), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(G128), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n842), .A2(new_n1158), .B1(new_n799), .B2(new_n404), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1157), .B(new_n1159), .C1(G137), .C2(new_n792), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n855), .A2(G125), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n782), .A2(new_n851), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT53), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n825), .A2(G132), .B1(G50), .B2(new_n826), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1160), .A2(new_n1161), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1074), .B1(new_n1155), .B2(new_n1165), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n759), .B(new_n1166), .C1(new_n1045), .C2(new_n862), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT118), .Z(new_n1168));
  AOI22_X1  g0968(.A1(new_n1147), .A2(new_n1085), .B1(new_n1150), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1149), .A2(new_n1169), .ZN(G378));
  INV_X1    g0970(.A(KEYINPUT121), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n284), .A2(new_n249), .A3(new_n315), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n323), .B1(new_n1172), .B2(new_n316), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n281), .A2(new_n277), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n889), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n323), .B(new_n1175), .C1(new_n1172), .C2(new_n316), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1179), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n921), .A2(new_n881), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT119), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1179), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1177), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1187), .A2(KEYINPUT119), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1184), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT40), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(new_n916), .B2(new_n902), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n910), .A2(new_n913), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1191), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1190), .B(G330), .C1(new_n1192), .C2(new_n1195), .ZN(new_n1196));
  AND3_X1   g0996(.A1(new_n1182), .A2(new_n1196), .A3(new_n938), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n938), .B1(new_n1182), .B2(new_n1196), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1171), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1182), .A2(new_n1196), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n938), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1182), .A2(new_n1196), .A3(new_n938), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1202), .A2(KEYINPUT121), .A3(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1111), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n881), .B(new_n869), .C1(new_n727), .C2(new_n728), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n1206), .A2(new_n1113), .B1(new_n915), .B2(new_n1116), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1121), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n1206), .B2(new_n1113), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n1112), .A2(new_n1207), .B1(new_n1209), .B2(new_n1119), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1205), .B1(new_n1145), .B2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1199), .A2(new_n1204), .A3(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT57), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1211), .B(KEYINPUT57), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(new_n746), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1214), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1199), .A2(new_n1204), .A3(new_n1085), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n759), .B1(new_n202), .B2(new_n862), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n810), .A2(new_n241), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1052), .B(new_n1221), .C1(G107), .C2(new_n825), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n793), .A2(new_n466), .B1(new_n842), .B2(new_n463), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n399), .A2(new_n443), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n802), .A2(new_n326), .ZN(new_n1225));
  NOR4_X1   g1025(.A1(new_n1223), .A2(new_n956), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1222), .B(new_n1226), .C1(new_n807), .C2(new_n815), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT58), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n792), .A2(G132), .B1(new_n805), .B2(G125), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n822), .A2(G137), .B1(new_n823), .B2(G150), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1232), .B1(new_n782), .B2(new_n1156), .C1(new_n1158), .C2(new_n788), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1233), .A2(KEYINPUT59), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(KEYINPUT59), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n826), .A2(G159), .ZN(new_n1236));
  AOI211_X1 g1036(.A(G33), .B(G41), .C1(new_n812), .C2(G124), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .A4(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1224), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1240));
  AND4_X1   g1040(.A1(new_n1229), .A2(new_n1238), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1220), .B1(new_n1241), .B2(new_n1074), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n1190), .B2(new_n772), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(KEYINPUT120), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1219), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1218), .A2(new_n1246), .ZN(G375));
  AOI22_X1  g1047(.A1(new_n783), .A2(G159), .B1(new_n855), .B2(G128), .ZN(new_n1248));
  XOR2_X1   g1048(.A(new_n1248), .B(KEYINPUT123), .Z(new_n1249));
  AOI22_X1  g1049(.A1(new_n805), .A2(G132), .B1(G50), .B2(new_n823), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n399), .B1(new_n822), .B2(G150), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1250), .B(new_n1251), .C1(new_n793), .C2(new_n1156), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n1221), .B(new_n1252), .C1(G137), .C2(new_n825), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1249), .A2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n961), .B1(new_n807), .B2(new_n788), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n399), .B1(new_n802), .B2(new_n336), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n793), .A2(new_n463), .B1(new_n842), .B2(new_n839), .ZN(new_n1257));
  NOR4_X1   g1057(.A1(new_n1255), .A2(new_n1057), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n1258), .B1(new_n466), .B2(new_n848), .C1(new_n843), .C2(new_n815), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1074), .B1(new_n1254), .B2(new_n1259), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n759), .B(new_n1260), .C1(new_n220), .C2(new_n862), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n1113), .B2(new_n773), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1030), .B1(new_n1118), .B2(new_n1123), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1262), .B1(new_n1263), .B2(KEYINPUT122), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT122), .ZN(new_n1265));
  NOR3_X1   g1065(.A1(new_n1210), .A2(new_n1265), .A3(new_n1030), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1118), .A2(new_n1123), .A3(new_n1111), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1125), .A2(new_n1026), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(G381));
  NOR2_X1   g1070(.A1(G375), .A2(G378), .ZN(new_n1271));
  OR2_X1    g1071(.A1(G393), .A2(G396), .ZN(new_n1272));
  NOR4_X1   g1072(.A1(G390), .A2(G381), .A3(G384), .A4(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(KEYINPUT124), .A3(new_n1041), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1271), .A2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT124), .B1(new_n1273), .B2(new_n1041), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1275), .A2(new_n1276), .ZN(G407));
  INV_X1    g1077(.A(G213), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1278), .B1(new_n1271), .B2(new_n682), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G407), .A2(new_n1279), .ZN(G409));
  INV_X1    g1080(.A(G390), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1040), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1026), .B1(new_n1028), .B2(new_n743), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1085), .B1(new_n1283), .B2(new_n985), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1282), .B1(new_n1284), .B2(new_n1029), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1281), .B1(new_n1285), .B2(new_n984), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1041), .A2(G390), .ZN(new_n1287));
  XNOR2_X1  g1087(.A(G393), .B(G396), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1286), .A2(new_n1287), .A3(KEYINPUT125), .A4(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT125), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1290), .B1(new_n1041), .B2(G390), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1288), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n682), .A2(G213), .A3(G2897), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1295), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1118), .A2(new_n1123), .A3(KEYINPUT60), .A4(new_n1111), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1297), .A2(new_n746), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT60), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1268), .B1(new_n1124), .B2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1267), .A2(new_n1301), .A3(G384), .ZN(new_n1302));
  AOI21_X1  g1102(.A(G384), .B1(new_n1267), .B2(new_n1301), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1296), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(G384), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1298), .A2(new_n1300), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1265), .B1(new_n1210), .B2(new_n1030), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1263), .A2(KEYINPUT122), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1307), .A2(new_n1308), .A3(new_n1262), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1305), .B1(new_n1306), .B2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1267), .A2(new_n1301), .A3(G384), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1310), .A2(new_n1311), .A3(new_n1295), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1304), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(G378), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1315), .B1(new_n1218), .B2(new_n1246), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1085), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1317));
  AND4_X1   g1117(.A1(new_n1149), .A2(new_n1317), .A3(new_n1169), .A4(new_n1244), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1199), .A2(new_n1204), .A3(new_n1026), .A4(new_n1211), .ZN(new_n1319));
  AOI22_X1  g1119(.A1(new_n1318), .A2(new_n1319), .B1(G213), .B2(new_n682), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1314), .B1(new_n1316), .B2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT61), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1216), .B1(new_n1213), .B2(new_n1212), .ZN(new_n1324));
  OAI21_X1  g1124(.A(G378), .B1(new_n1324), .B2(new_n1245), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT62), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1325), .A2(new_n1320), .A3(new_n1326), .A4(new_n1327), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1322), .A2(new_n1323), .A3(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1325), .A2(new_n1320), .A3(new_n1327), .ZN(new_n1330));
  AND2_X1   g1130(.A1(new_n1330), .A2(KEYINPUT62), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1289), .B(new_n1294), .C1(new_n1329), .C2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(KEYINPUT63), .ZN(new_n1333));
  OR2_X1    g1133(.A1(new_n1330), .A2(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1313), .B1(new_n1325), .B2(new_n1320), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1330), .B1(new_n1335), .B2(new_n1333), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT61), .B1(new_n1294), .B2(new_n1289), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT126), .ZN(new_n1338));
  OAI211_X1 g1138(.A(new_n1334), .B(new_n1336), .C1(new_n1337), .C2(new_n1338), .ZN(new_n1339));
  AOI211_X1 g1139(.A(KEYINPUT126), .B(KEYINPUT61), .C1(new_n1294), .C2(new_n1289), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1332), .B1(new_n1339), .B2(new_n1340), .ZN(G405));
  INV_X1    g1141(.A(KEYINPUT127), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1327), .A2(new_n1342), .ZN(new_n1343));
  NOR3_X1   g1143(.A1(new_n1271), .A2(new_n1316), .A3(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1327), .A2(new_n1342), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1294), .A2(new_n1289), .A3(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1346), .B1(new_n1294), .B2(new_n1289), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1345), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1349), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1351), .A2(new_n1344), .A3(new_n1347), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1350), .A2(new_n1352), .ZN(G402));
endmodule


