

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587;

  OR2_X1 U322 ( .A1(n570), .A2(n454), .ZN(n456) );
  XNOR2_X1 U323 ( .A(n339), .B(n338), .ZN(n347) );
  NOR2_X1 U324 ( .A1(n466), .A2(n457), .ZN(n458) );
  XNOR2_X1 U325 ( .A(n388), .B(KEYINPUT47), .ZN(n389) );
  XNOR2_X1 U326 ( .A(n337), .B(KEYINPUT74), .ZN(n338) );
  XNOR2_X1 U327 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U328 ( .A(n347), .B(n346), .ZN(n393) );
  XNOR2_X1 U329 ( .A(n349), .B(KEYINPUT41), .ZN(n550) );
  XNOR2_X1 U330 ( .A(n459), .B(n458), .ZN(n568) );
  INV_X1 U331 ( .A(n550), .ZN(n564) );
  XOR2_X1 U332 ( .A(n329), .B(n328), .Z(n531) );
  XOR2_X1 U333 ( .A(KEYINPUT28), .B(n472), .Z(n526) );
  XNOR2_X1 U334 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n460) );
  XOR2_X1 U335 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n291) );
  XNOR2_X1 U336 ( .A(G162GAT), .B(G106GAT), .ZN(n290) );
  XNOR2_X1 U337 ( .A(n291), .B(n290), .ZN(n308) );
  XOR2_X1 U338 ( .A(KEYINPUT68), .B(KEYINPUT10), .Z(n293) );
  XNOR2_X1 U339 ( .A(G92GAT), .B(G218GAT), .ZN(n292) );
  XNOR2_X1 U340 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U341 ( .A(KEYINPUT67), .B(KEYINPUT66), .Z(n295) );
  XNOR2_X1 U342 ( .A(G43GAT), .B(G99GAT), .ZN(n294) );
  XNOR2_X1 U343 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U344 ( .A(n297), .B(n296), .Z(n306) );
  XOR2_X1 U345 ( .A(KEYINPUT7), .B(G50GAT), .Z(n299) );
  XNOR2_X1 U346 ( .A(G36GAT), .B(G29GAT), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U348 ( .A(KEYINPUT8), .B(n300), .Z(n363) );
  XNOR2_X1 U349 ( .A(G85GAT), .B(KEYINPUT75), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n301), .B(KEYINPUT76), .ZN(n341) );
  XOR2_X1 U351 ( .A(G190GAT), .B(G134GAT), .Z(n312) );
  XOR2_X1 U352 ( .A(n341), .B(n312), .Z(n303) );
  NAND2_X1 U353 ( .A1(G232GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U354 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n363), .B(n304), .ZN(n305) );
  XNOR2_X1 U356 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n555) );
  INV_X1 U358 ( .A(KEYINPUT123), .ZN(n459) );
  XOR2_X1 U359 ( .A(KEYINPUT65), .B(KEYINPUT20), .Z(n310) );
  XNOR2_X1 U360 ( .A(KEYINPUT86), .B(KEYINPUT87), .ZN(n309) );
  XNOR2_X1 U361 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U362 ( .A(n312), .B(n311), .Z(n314) );
  NAND2_X1 U363 ( .A1(G227GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U364 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U365 ( .A(n315), .B(KEYINPUT85), .Z(n318) );
  XNOR2_X1 U366 ( .A(G43GAT), .B(G15GAT), .ZN(n316) );
  XNOR2_X1 U367 ( .A(n316), .B(G113GAT), .ZN(n359) );
  XNOR2_X1 U368 ( .A(n359), .B(KEYINPUT84), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n321) );
  XOR2_X1 U370 ( .A(KEYINPUT0), .B(KEYINPUT83), .Z(n320) );
  XNOR2_X1 U371 ( .A(G127GAT), .B(KEYINPUT82), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n320), .B(n319), .ZN(n432) );
  XOR2_X1 U373 ( .A(n321), .B(n432), .Z(n329) );
  XOR2_X1 U374 ( .A(KEYINPUT88), .B(KEYINPUT19), .Z(n323) );
  XNOR2_X1 U375 ( .A(G176GAT), .B(KEYINPUT18), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U377 ( .A(n324), .B(G183GAT), .Z(n326) );
  XNOR2_X1 U378 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n325) );
  XNOR2_X1 U379 ( .A(n326), .B(n325), .ZN(n403) );
  XNOR2_X1 U380 ( .A(G99GAT), .B(G71GAT), .ZN(n327) );
  XNOR2_X1 U381 ( .A(n327), .B(G120GAT), .ZN(n330) );
  XNOR2_X1 U382 ( .A(n403), .B(n330), .ZN(n328) );
  INV_X1 U383 ( .A(n531), .ZN(n466) );
  XOR2_X1 U384 ( .A(G57GAT), .B(KEYINPUT13), .Z(n371) );
  XNOR2_X1 U385 ( .A(n330), .B(n371), .ZN(n334) );
  INV_X1 U386 ( .A(n334), .ZN(n332) );
  AND2_X1 U387 ( .A1(G230GAT), .A2(G233GAT), .ZN(n333) );
  INV_X1 U388 ( .A(n333), .ZN(n331) );
  NAND2_X1 U389 ( .A1(n332), .A2(n331), .ZN(n336) );
  NAND2_X1 U390 ( .A1(n334), .A2(n333), .ZN(n335) );
  NAND2_X1 U391 ( .A1(n336), .A2(n335), .ZN(n339) );
  XOR2_X1 U392 ( .A(G92GAT), .B(G64GAT), .Z(n400) );
  XOR2_X1 U393 ( .A(n400), .B(KEYINPUT31), .Z(n337) );
  XNOR2_X1 U394 ( .A(G148GAT), .B(G106GAT), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n340), .B(G78GAT), .ZN(n441) );
  XNOR2_X1 U396 ( .A(n341), .B(n441), .ZN(n345) );
  XOR2_X1 U397 ( .A(KEYINPUT32), .B(G204GAT), .Z(n343) );
  XNOR2_X1 U398 ( .A(G176GAT), .B(KEYINPUT33), .ZN(n342) );
  XOR2_X1 U399 ( .A(n343), .B(n342), .Z(n344) );
  INV_X1 U400 ( .A(KEYINPUT64), .ZN(n348) );
  XNOR2_X1 U401 ( .A(n393), .B(n348), .ZN(n349) );
  XOR2_X1 U402 ( .A(KEYINPUT29), .B(KEYINPUT72), .Z(n351) );
  XNOR2_X1 U403 ( .A(KEYINPUT30), .B(KEYINPUT70), .ZN(n350) );
  XNOR2_X1 U404 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U405 ( .A(KEYINPUT69), .B(KEYINPUT71), .Z(n353) );
  XOR2_X1 U406 ( .A(G141GAT), .B(G22GAT), .Z(n439) );
  XOR2_X1 U407 ( .A(G197GAT), .B(G8GAT), .Z(n402) );
  XNOR2_X1 U408 ( .A(n439), .B(n402), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U410 ( .A(n355), .B(n354), .Z(n357) );
  NAND2_X1 U411 ( .A1(G229GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U413 ( .A(n358), .B(G1GAT), .Z(n361) );
  XNOR2_X1 U414 ( .A(G169GAT), .B(n359), .ZN(n360) );
  XNOR2_X1 U415 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U416 ( .A(n363), .B(n362), .ZN(n574) );
  NOR2_X1 U417 ( .A1(n550), .A2(n574), .ZN(n364) );
  XNOR2_X1 U418 ( .A(n364), .B(KEYINPUT46), .ZN(n385) );
  XOR2_X1 U419 ( .A(G8GAT), .B(G22GAT), .Z(n366) );
  XNOR2_X1 U420 ( .A(G15GAT), .B(G1GAT), .ZN(n365) );
  XNOR2_X1 U421 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U422 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n368) );
  XNOR2_X1 U423 ( .A(G71GAT), .B(G78GAT), .ZN(n367) );
  XNOR2_X1 U424 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U425 ( .A(n370), .B(n369), .Z(n376) );
  XOR2_X1 U426 ( .A(n371), .B(G155GAT), .Z(n373) );
  NAND2_X1 U427 ( .A1(G231GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U429 ( .A(G127GAT), .B(n374), .ZN(n375) );
  XNOR2_X1 U430 ( .A(n376), .B(n375), .ZN(n384) );
  XOR2_X1 U431 ( .A(KEYINPUT81), .B(KEYINPUT78), .Z(n378) );
  XNOR2_X1 U432 ( .A(KEYINPUT80), .B(KEYINPUT15), .ZN(n377) );
  XNOR2_X1 U433 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U434 ( .A(G211GAT), .B(KEYINPUT79), .Z(n380) );
  XNOR2_X1 U435 ( .A(G183GAT), .B(G64GAT), .ZN(n379) );
  XNOR2_X1 U436 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U437 ( .A(n382), .B(n381), .Z(n383) );
  XOR2_X1 U438 ( .A(n384), .B(n383), .Z(n567) );
  NOR2_X1 U439 ( .A1(n385), .A2(n567), .ZN(n386) );
  XNOR2_X1 U440 ( .A(n386), .B(KEYINPUT113), .ZN(n387) );
  NOR2_X1 U441 ( .A1(n555), .A2(n387), .ZN(n390) );
  INV_X1 U442 ( .A(KEYINPUT114), .ZN(n388) );
  XNOR2_X1 U443 ( .A(n390), .B(n389), .ZN(n398) );
  XNOR2_X1 U444 ( .A(KEYINPUT73), .B(n574), .ZN(n559) );
  XOR2_X1 U445 ( .A(n555), .B(KEYINPUT106), .Z(n391) );
  XNOR2_X1 U446 ( .A(n391), .B(KEYINPUT36), .ZN(n585) );
  INV_X1 U447 ( .A(n567), .ZN(n581) );
  NOR2_X1 U448 ( .A1(n585), .A2(n581), .ZN(n392) );
  XNOR2_X1 U449 ( .A(KEYINPUT45), .B(n392), .ZN(n394) );
  NAND2_X1 U450 ( .A1(n394), .A2(n393), .ZN(n395) );
  XOR2_X1 U451 ( .A(KEYINPUT115), .B(n395), .Z(n396) );
  NOR2_X1 U452 ( .A1(n559), .A2(n396), .ZN(n397) );
  NOR2_X1 U453 ( .A1(n398), .A2(n397), .ZN(n399) );
  XNOR2_X1 U454 ( .A(n399), .B(KEYINPUT48), .ZN(n530) );
  XNOR2_X1 U455 ( .A(G36GAT), .B(G190GAT), .ZN(n401) );
  XOR2_X1 U456 ( .A(n401), .B(n400), .Z(n412) );
  XOR2_X1 U457 ( .A(n403), .B(n402), .Z(n405) );
  NAND2_X1 U458 ( .A1(G226GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U459 ( .A(n405), .B(n404), .ZN(n408) );
  XOR2_X1 U460 ( .A(KEYINPUT21), .B(G211GAT), .Z(n407) );
  XNOR2_X1 U461 ( .A(G204GAT), .B(G218GAT), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n448) );
  XOR2_X1 U463 ( .A(n408), .B(n448), .Z(n410) );
  XNOR2_X1 U464 ( .A(KEYINPUT98), .B(KEYINPUT97), .ZN(n409) );
  XNOR2_X1 U465 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U466 ( .A(n412), .B(n411), .Z(n521) );
  INV_X1 U467 ( .A(n521), .ZN(n413) );
  NOR2_X1 U468 ( .A1(n530), .A2(n413), .ZN(n415) );
  INV_X1 U469 ( .A(KEYINPUT54), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n415), .B(n414), .ZN(n570) );
  NAND2_X1 U471 ( .A1(G225GAT), .A2(G233GAT), .ZN(n421) );
  XOR2_X1 U472 ( .A(G85GAT), .B(G141GAT), .Z(n417) );
  XNOR2_X1 U473 ( .A(G113GAT), .B(G1GAT), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n417), .B(n416), .ZN(n419) );
  XOR2_X1 U475 ( .A(G29GAT), .B(G134GAT), .Z(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n438) );
  XOR2_X1 U478 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n423) );
  XNOR2_X1 U479 ( .A(KEYINPUT1), .B(KEYINPUT92), .ZN(n422) );
  XNOR2_X1 U480 ( .A(n423), .B(n422), .ZN(n436) );
  XOR2_X1 U481 ( .A(KEYINPUT4), .B(G148GAT), .Z(n425) );
  XNOR2_X1 U482 ( .A(G120GAT), .B(G57GAT), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U484 ( .A(KEYINPUT95), .B(KEYINPUT6), .Z(n427) );
  XNOR2_X1 U485 ( .A(KEYINPUT93), .B(KEYINPUT94), .ZN(n426) );
  XNOR2_X1 U486 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U487 ( .A(n429), .B(n428), .Z(n434) );
  XOR2_X1 U488 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n431) );
  XNOR2_X1 U489 ( .A(G162GAT), .B(G155GAT), .ZN(n430) );
  XNOR2_X1 U490 ( .A(n431), .B(n430), .ZN(n449) );
  XNOR2_X1 U491 ( .A(n432), .B(n449), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U493 ( .A(n436), .B(n435), .Z(n437) );
  XOR2_X1 U494 ( .A(n438), .B(n437), .Z(n479) );
  XNOR2_X1 U495 ( .A(G50GAT), .B(n439), .ZN(n440) );
  XNOR2_X1 U496 ( .A(n440), .B(G197GAT), .ZN(n453) );
  XOR2_X1 U497 ( .A(KEYINPUT91), .B(n441), .Z(n443) );
  NAND2_X1 U498 ( .A1(G228GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n447) );
  XOR2_X1 U500 ( .A(KEYINPUT90), .B(KEYINPUT22), .Z(n445) );
  XNOR2_X1 U501 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n444) );
  XNOR2_X1 U502 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U503 ( .A(n447), .B(n446), .Z(n451) );
  XNOR2_X1 U504 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U505 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U506 ( .A(n453), .B(n452), .ZN(n472) );
  NAND2_X1 U507 ( .A1(n479), .A2(n472), .ZN(n454) );
  XOR2_X1 U508 ( .A(KEYINPUT122), .B(KEYINPUT55), .Z(n455) );
  XNOR2_X1 U509 ( .A(n456), .B(n455), .ZN(n457) );
  NAND2_X1 U510 ( .A1(n555), .A2(n568), .ZN(n461) );
  XNOR2_X1 U511 ( .A(n461), .B(n460), .ZN(G1351GAT) );
  XNOR2_X1 U512 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n462) );
  XNOR2_X1 U513 ( .A(n462), .B(KEYINPUT101), .ZN(n463) );
  XOR2_X1 U514 ( .A(KEYINPUT102), .B(n463), .Z(n484) );
  NAND2_X1 U515 ( .A1(n393), .A2(n559), .ZN(n464) );
  XOR2_X1 U516 ( .A(KEYINPUT77), .B(n464), .Z(n496) );
  NOR2_X1 U517 ( .A1(n555), .A2(n581), .ZN(n465) );
  XNOR2_X1 U518 ( .A(n465), .B(KEYINPUT16), .ZN(n482) );
  INV_X1 U519 ( .A(n479), .ZN(n571) );
  XNOR2_X1 U520 ( .A(n521), .B(KEYINPUT27), .ZN(n475) );
  NAND2_X1 U521 ( .A1(n571), .A2(n475), .ZN(n529) );
  XOR2_X1 U522 ( .A(KEYINPUT89), .B(n466), .Z(n467) );
  INV_X1 U523 ( .A(n526), .ZN(n533) );
  NAND2_X1 U524 ( .A1(n467), .A2(n533), .ZN(n468) );
  NOR2_X1 U525 ( .A1(n529), .A2(n468), .ZN(n469) );
  XNOR2_X1 U526 ( .A(KEYINPUT99), .B(n469), .ZN(n481) );
  NAND2_X1 U527 ( .A1(n531), .A2(n521), .ZN(n470) );
  NAND2_X1 U528 ( .A1(n472), .A2(n470), .ZN(n471) );
  XOR2_X1 U529 ( .A(KEYINPUT25), .B(n471), .Z(n477) );
  NOR2_X1 U530 ( .A1(n531), .A2(n472), .ZN(n474) );
  XNOR2_X1 U531 ( .A(KEYINPUT100), .B(KEYINPUT26), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n474), .B(n473), .ZN(n572) );
  NAND2_X1 U533 ( .A1(n475), .A2(n572), .ZN(n476) );
  NAND2_X1 U534 ( .A1(n477), .A2(n476), .ZN(n478) );
  NAND2_X1 U535 ( .A1(n479), .A2(n478), .ZN(n480) );
  NAND2_X1 U536 ( .A1(n481), .A2(n480), .ZN(n493) );
  NAND2_X1 U537 ( .A1(n482), .A2(n493), .ZN(n508) );
  NOR2_X1 U538 ( .A1(n496), .A2(n508), .ZN(n491) );
  NAND2_X1 U539 ( .A1(n491), .A2(n571), .ZN(n483) );
  XNOR2_X1 U540 ( .A(n484), .B(n483), .ZN(G1324GAT) );
  XOR2_X1 U541 ( .A(G8GAT), .B(KEYINPUT103), .Z(n486) );
  NAND2_X1 U542 ( .A1(n491), .A2(n521), .ZN(n485) );
  XNOR2_X1 U543 ( .A(n486), .B(n485), .ZN(G1325GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT105), .B(KEYINPUT35), .Z(n488) );
  NAND2_X1 U545 ( .A1(n491), .A2(n531), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n488), .B(n487), .ZN(n490) );
  XOR2_X1 U547 ( .A(G15GAT), .B(KEYINPUT104), .Z(n489) );
  XNOR2_X1 U548 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  NAND2_X1 U549 ( .A1(n526), .A2(n491), .ZN(n492) );
  XNOR2_X1 U550 ( .A(n492), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U551 ( .A1(n581), .A2(n493), .ZN(n494) );
  NOR2_X1 U552 ( .A1(n585), .A2(n494), .ZN(n495) );
  XNOR2_X1 U553 ( .A(KEYINPUT37), .B(n495), .ZN(n519) );
  NOR2_X1 U554 ( .A1(n519), .A2(n496), .ZN(n497) );
  XNOR2_X1 U555 ( .A(KEYINPUT38), .B(n497), .ZN(n504) );
  NAND2_X1 U556 ( .A1(n571), .A2(n504), .ZN(n499) );
  XOR2_X1 U557 ( .A(G29GAT), .B(KEYINPUT39), .Z(n498) );
  XNOR2_X1 U558 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  XOR2_X1 U559 ( .A(G36GAT), .B(KEYINPUT107), .Z(n501) );
  NAND2_X1 U560 ( .A1(n504), .A2(n521), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n501), .B(n500), .ZN(G1329GAT) );
  NAND2_X1 U562 ( .A1(n504), .A2(n531), .ZN(n502) );
  XNOR2_X1 U563 ( .A(n502), .B(KEYINPUT40), .ZN(n503) );
  XNOR2_X1 U564 ( .A(G43GAT), .B(n503), .ZN(G1330GAT) );
  XNOR2_X1 U565 ( .A(G50GAT), .B(KEYINPUT108), .ZN(n506) );
  NAND2_X1 U566 ( .A1(n526), .A2(n504), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n506), .B(n505), .ZN(G1331GAT) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n510) );
  NAND2_X1 U569 ( .A1(n574), .A2(n564), .ZN(n507) );
  XOR2_X1 U570 ( .A(KEYINPUT109), .B(n507), .Z(n518) );
  NOR2_X1 U571 ( .A1(n518), .A2(n508), .ZN(n515) );
  NAND2_X1 U572 ( .A1(n571), .A2(n515), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(G1332GAT) );
  NAND2_X1 U574 ( .A1(n521), .A2(n515), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n511), .B(KEYINPUT110), .ZN(n512) );
  XNOR2_X1 U576 ( .A(G64GAT), .B(n512), .ZN(G1333GAT) );
  XOR2_X1 U577 ( .A(G71GAT), .B(KEYINPUT111), .Z(n514) );
  NAND2_X1 U578 ( .A1(n515), .A2(n531), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .Z(n517) );
  NAND2_X1 U581 ( .A1(n515), .A2(n526), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NOR2_X1 U583 ( .A1(n519), .A2(n518), .ZN(n525) );
  NAND2_X1 U584 ( .A1(n571), .A2(n525), .ZN(n520) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(n520), .ZN(G1336GAT) );
  NAND2_X1 U586 ( .A1(n521), .A2(n525), .ZN(n522) );
  XNOR2_X1 U587 ( .A(n522), .B(KEYINPUT112), .ZN(n523) );
  XNOR2_X1 U588 ( .A(G92GAT), .B(n523), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n531), .A2(n525), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n524), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n527), .B(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  NOR2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n545) );
  NAND2_X1 U595 ( .A1(n545), .A2(n531), .ZN(n532) );
  XOR2_X1 U596 ( .A(KEYINPUT116), .B(n532), .Z(n534) );
  NAND2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U598 ( .A(n535), .B(KEYINPUT117), .ZN(n542) );
  NAND2_X1 U599 ( .A1(n542), .A2(n559), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n536), .B(KEYINPUT118), .ZN(n537) );
  XNOR2_X1 U601 ( .A(G113GAT), .B(n537), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(G120GAT), .B(KEYINPUT49), .Z(n539) );
  NAND2_X1 U603 ( .A1(n542), .A2(n564), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  NAND2_X1 U605 ( .A1(n542), .A2(n567), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n540), .B(KEYINPUT50), .ZN(n541) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U609 ( .A1(n542), .A2(n555), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NAND2_X1 U611 ( .A1(n545), .A2(n572), .ZN(n556) );
  NOR2_X1 U612 ( .A1(n574), .A2(n556), .ZN(n547) );
  XNOR2_X1 U613 ( .A(G141GAT), .B(KEYINPUT119), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT120), .B(KEYINPUT52), .Z(n549) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n548) );
  XNOR2_X1 U617 ( .A(n549), .B(n548), .ZN(n552) );
  NOR2_X1 U618 ( .A1(n550), .A2(n556), .ZN(n551) );
  XOR2_X1 U619 ( .A(n552), .B(n551), .Z(G1345GAT) );
  NOR2_X1 U620 ( .A1(n581), .A2(n556), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(KEYINPUT121), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(G1346GAT) );
  INV_X1 U623 ( .A(n555), .ZN(n557) );
  NOR2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U625 ( .A(G162GAT), .B(n558), .Z(G1347GAT) );
  NAND2_X1 U626 ( .A1(n568), .A2(n559), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n560), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n562) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(n563) );
  XOR2_X1 U631 ( .A(KEYINPUT56), .B(n563), .Z(n566) );
  NAND2_X1 U632 ( .A1(n568), .A2(n564), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(G1349GAT) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U636 ( .A(KEYINPUT126), .B(KEYINPUT59), .ZN(n578) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n584) );
  NOR2_X1 U639 ( .A1(n574), .A2(n584), .ZN(n576) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n578), .B(n577), .ZN(G1352GAT) );
  NOR2_X1 U643 ( .A1(n393), .A2(n584), .ZN(n580) );
  XNOR2_X1 U644 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n584), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(n586), .Z(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

