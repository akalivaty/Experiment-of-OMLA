//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G128), .ZN(new_n188));
  OR2_X1    g002(.A1(new_n188), .A2(KEYINPUT23), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(KEYINPUT23), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  OAI211_X1 g005(.A(new_n189), .B(new_n190), .C1(G119), .C2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G119), .B(G128), .ZN(new_n193));
  XOR2_X1   g007(.A(KEYINPUT24), .B(G110), .Z(new_n194));
  OAI22_X1  g008(.A1(new_n192), .A2(G110), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G125), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n196), .A2(KEYINPUT16), .A3(G140), .ZN(new_n197));
  OR2_X1    g011(.A1(G125), .A2(G140), .ZN(new_n198));
  NAND2_X1  g012(.A1(G125), .A2(G140), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n197), .B1(new_n200), .B2(KEYINPUT16), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  AND2_X1   g017(.A1(G125), .A2(G140), .ZN(new_n204));
  NOR2_X1   g018(.A1(G125), .A2(G140), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n195), .A2(new_n202), .A3(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(new_n201), .B(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n192), .A2(G110), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n194), .A2(new_n193), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT73), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n207), .A2(new_n211), .A3(KEYINPUT73), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT22), .B(G137), .ZN(new_n216));
  INV_X1    g030(.A(G953), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(G221), .A3(G234), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n216), .B(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n214), .A2(new_n215), .A3(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n212), .A2(new_n213), .A3(new_n219), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G217), .ZN(new_n224));
  INV_X1    g038(.A(G902), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n224), .B1(G234), .B2(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(G902), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT74), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n228), .B(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT25), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n231), .B1(new_n223), .B2(new_n225), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n223), .A2(new_n231), .A3(new_n225), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n226), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(G472), .A2(G902), .ZN(new_n237));
  INV_X1    g051(.A(G137), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT67), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G137), .ZN(new_n241));
  INV_X1    g055(.A(G134), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n239), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n238), .A2(G134), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G131), .ZN(new_n246));
  NAND2_X1  g060(.A1(KEYINPUT11), .A2(G134), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n240), .A2(G137), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n238), .A2(KEYINPUT67), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n238), .A2(G134), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n254), .B1(new_n242), .B2(G137), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT66), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI211_X1 g071(.A(KEYINPUT66), .B(new_n254), .C1(new_n242), .C2(G137), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n251), .A2(new_n253), .A3(new_n257), .A4(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n246), .B1(new_n259), .B2(G131), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n203), .A2(G143), .ZN(new_n261));
  INV_X1    g075(.A(G143), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT64), .B1(new_n262), .B2(G146), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT64), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(new_n203), .A3(G143), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n261), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT1), .B1(new_n262), .B2(G146), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT68), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n203), .A2(G143), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n271), .A3(KEYINPUT1), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n269), .A2(G128), .A3(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT65), .B1(new_n203), .B2(G143), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT65), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n262), .A3(G146), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n274), .A2(new_n276), .B1(G143), .B2(new_n203), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT1), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n278), .B1(G143), .B2(new_n203), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n279), .A2(new_n191), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n267), .A2(new_n273), .B1(new_n277), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n260), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n275), .B1(new_n262), .B2(G146), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n203), .A2(KEYINPUT65), .A3(G143), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n270), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(KEYINPUT0), .A2(G128), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(KEYINPUT0), .A2(G128), .ZN(new_n288));
  OR2_X1    g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI22_X1  g103(.A1(new_n285), .A2(new_n286), .B1(new_n266), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT67), .B(G137), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n253), .B1(new_n291), .B2(new_n247), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n257), .A2(new_n258), .ZN(new_n293));
  OAI21_X1  g107(.A(G131), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n258), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT66), .B1(new_n244), .B2(new_n254), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G131), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n239), .A2(new_n241), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n252), .B1(new_n299), .B2(new_n248), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n290), .B1(new_n294), .B2(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(KEYINPUT70), .B(KEYINPUT30), .C1(new_n282), .C2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n290), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n292), .A2(new_n293), .A3(G131), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n298), .B1(new_n297), .B2(new_n300), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n277), .A2(new_n280), .ZN(new_n308));
  OAI21_X1  g122(.A(G128), .B1(new_n268), .B2(KEYINPUT68), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n271), .B1(new_n270), .B2(KEYINPUT1), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n308), .B1(new_n311), .B2(new_n266), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(new_n301), .A3(new_n246), .ZN(new_n313));
  OR2_X1    g127(.A1(KEYINPUT70), .A2(KEYINPUT30), .ZN(new_n314));
  NAND2_X1  g128(.A1(KEYINPUT70), .A2(KEYINPUT30), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n307), .A2(new_n313), .A3(new_n314), .A4(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n303), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n187), .A2(G116), .ZN(new_n318));
  INV_X1    g132(.A(G116), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G119), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT2), .B(G113), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n321), .B(KEYINPUT69), .ZN(new_n325));
  INV_X1    g139(.A(new_n322), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n317), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT31), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n318), .A2(new_n320), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n330), .B(KEYINPUT69), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n323), .B1(new_n331), .B2(new_n322), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n307), .A2(new_n313), .A3(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(G237), .A2(G953), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G210), .ZN(new_n335));
  INV_X1    g149(.A(G101), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n335), .B(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n337), .B(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n328), .A2(new_n329), .A3(new_n333), .A4(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n341), .A2(KEYINPUT71), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT71), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n332), .B1(new_n303), .B2(new_n316), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n282), .A2(new_n302), .A3(new_n327), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n344), .A2(new_n345), .A3(new_n339), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n343), .B1(new_n346), .B2(new_n329), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n342), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n328), .A2(new_n333), .A3(new_n340), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT31), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT72), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT28), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n327), .B1(new_n282), .B2(new_n302), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n352), .B1(new_n353), .B2(new_n333), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n333), .A2(new_n352), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n351), .B1(new_n357), .B2(new_n340), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n332), .B1(new_n307), .B2(new_n313), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT28), .B1(new_n345), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n340), .B1(new_n360), .B2(new_n355), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT72), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n350), .A2(new_n358), .A3(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n237), .B1(new_n348), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(KEYINPUT32), .ZN(new_n365));
  AOI22_X1  g179(.A1(new_n349), .A2(KEYINPUT31), .B1(new_n361), .B2(KEYINPUT72), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n366), .B(new_n358), .C1(new_n342), .C2(new_n347), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT32), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n368), .A3(new_n237), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n365), .A2(new_n369), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n354), .A2(new_n356), .A3(new_n339), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT29), .ZN(new_n372));
  OR2_X1    g186(.A1(new_n371), .A2(KEYINPUT29), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n344), .A2(new_n345), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(new_n340), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n225), .B(new_n372), .C1(new_n373), .C2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G472), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n236), .B1(new_n370), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G237), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n217), .A3(G214), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n262), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n334), .A2(G143), .A3(G214), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G131), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n381), .A2(new_n298), .A3(new_n382), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(KEYINPUT17), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n383), .A2(KEYINPUT17), .A3(G131), .ZN(new_n388));
  OR3_X1    g202(.A1(new_n387), .A2(new_n208), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(KEYINPUT18), .A2(G131), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n381), .A2(new_n382), .A3(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n198), .A2(G146), .A3(new_n199), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n206), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT84), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n334), .A2(G143), .A3(G214), .ZN(new_n396));
  AOI21_X1  g210(.A(G143), .B1(new_n334), .B2(G214), .ZN(new_n397));
  OAI211_X1 g211(.A(KEYINPUT18), .B(G131), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n394), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n398), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n391), .A2(new_n393), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT84), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G113), .B(G122), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(G104), .ZN(new_n405));
  XOR2_X1   g219(.A(new_n405), .B(KEYINPUT88), .Z(new_n406));
  NAND3_X1  g220(.A1(new_n389), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n405), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n409), .B1(new_n389), .B2(new_n403), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n225), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G475), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT20), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT85), .ZN(new_n414));
  AOI21_X1  g228(.A(KEYINPUT19), .B1(new_n200), .B2(new_n414), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n414), .B(KEYINPUT19), .C1(new_n204), .C2(new_n205), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n203), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n386), .A2(new_n202), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n395), .B1(new_n394), .B2(new_n398), .ZN(new_n420));
  AND4_X1   g234(.A1(new_n395), .A2(new_n398), .A3(new_n391), .A4(new_n393), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT86), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n403), .A2(KEYINPUT86), .A3(new_n419), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n405), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT87), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n424), .A2(new_n425), .A3(KEYINPUT87), .A4(new_n405), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(G475), .B1(new_n430), .B2(new_n407), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n413), .B1(new_n431), .B2(new_n225), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n408), .B1(new_n428), .B2(new_n429), .ZN(new_n433));
  NOR4_X1   g247(.A1(new_n433), .A2(KEYINPUT20), .A3(G475), .A4(G902), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n412), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT89), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT89), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n437), .B(new_n412), .C1(new_n432), .C2(new_n434), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT93), .ZN(new_n439));
  INV_X1    g253(.A(G122), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(G116), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n440), .A2(G116), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT14), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n444), .B(KEYINPUT91), .ZN(new_n445));
  INV_X1    g259(.A(new_n442), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n446), .A2(KEYINPUT14), .ZN(new_n447));
  OAI21_X1  g261(.A(G107), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n446), .A2(new_n441), .ZN(new_n449));
  INV_X1    g263(.A(G107), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n191), .A2(G143), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n191), .A2(G143), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(new_n242), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n448), .A2(new_n451), .A3(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n449), .B(new_n450), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n455), .A2(new_n242), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n452), .B1(new_n454), .B2(KEYINPUT13), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT90), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n460), .A2(new_n461), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n454), .A2(KEYINPUT13), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n458), .B(new_n459), .C1(new_n465), .C2(new_n242), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n457), .A2(new_n466), .ZN(new_n467));
  XOR2_X1   g281(.A(KEYINPUT9), .B(G234), .Z(new_n468));
  NAND3_X1  g282(.A1(new_n468), .A2(G217), .A3(new_n217), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n469), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n457), .A2(new_n466), .A3(new_n471), .ZN(new_n472));
  AOI211_X1 g286(.A(new_n439), .B(G902), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n470), .A2(new_n472), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n225), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT92), .ZN(new_n476));
  AOI21_X1  g290(.A(G902), .B1(new_n470), .B2(new_n472), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT92), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n473), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G478), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n481), .A2(KEYINPUT15), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n482), .B1(new_n477), .B2(new_n439), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n436), .A2(new_n438), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n468), .ZN(new_n488));
  OAI21_X1  g302(.A(G221), .B1(new_n488), .B2(G902), .ZN(new_n489));
  XOR2_X1   g303(.A(new_n489), .B(KEYINPUT75), .Z(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G469), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n305), .A2(new_n306), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT78), .ZN(new_n495));
  INV_X1    g309(.A(G104), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n496), .A2(KEYINPUT77), .A3(G107), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT3), .B1(new_n497), .B2(KEYINPUT76), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT77), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(new_n450), .A3(G104), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT76), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT3), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n450), .A2(KEYINPUT76), .A3(G104), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n496), .A2(G107), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n504), .A2(new_n336), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n450), .A2(G104), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n506), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(G101), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n191), .B1(new_n279), .B2(new_n271), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n266), .B1(new_n512), .B2(new_n269), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n277), .A2(new_n280), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT10), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n495), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT10), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n267), .A2(new_n273), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n517), .B1(new_n518), .B2(new_n308), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n519), .A2(KEYINPUT78), .A3(new_n507), .A4(new_n510), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n502), .B1(new_n500), .B2(new_n501), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n505), .B(new_n506), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(G101), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(KEYINPUT4), .A3(new_n507), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT4), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n524), .A2(new_n527), .A3(G101), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n304), .A3(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n277), .B(new_n280), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n530), .A2(new_n507), .A3(new_n510), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n517), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n494), .B1(new_n521), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n516), .A2(new_n520), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n535), .A2(new_n493), .A3(new_n529), .A4(new_n532), .ZN(new_n536));
  XNOR2_X1  g350(.A(G110), .B(G140), .ZN(new_n537));
  INV_X1    g351(.A(G227), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(G953), .ZN(new_n539));
  XOR2_X1   g353(.A(new_n537), .B(new_n539), .Z(new_n540));
  AND3_X1   g354(.A1(new_n534), .A2(new_n536), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n531), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n312), .B1(new_n507), .B2(new_n510), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n494), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT12), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n511), .A2(new_n281), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n493), .B1(new_n547), .B2(new_n531), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT12), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n540), .B1(new_n550), .B2(new_n536), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT79), .B1(new_n541), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n544), .A2(new_n545), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n548), .A2(KEYINPUT12), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n536), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n540), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT79), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n534), .A2(new_n536), .A3(new_n540), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n492), .B1(new_n552), .B2(new_n560), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n550), .A2(new_n536), .A3(new_n540), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n540), .B1(new_n534), .B2(new_n536), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n492), .B(new_n225), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n492), .A2(new_n225), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n491), .B1(new_n561), .B2(new_n567), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n217), .A2(G952), .ZN(new_n569));
  NAND2_X1  g383(.A1(G234), .A2(G237), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  XOR2_X1   g386(.A(KEYINPUT21), .B(G898), .Z(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n570), .A2(G902), .A3(G953), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n572), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(G214), .B1(G237), .B2(G902), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n526), .A2(new_n327), .A3(new_n528), .ZN(new_n580));
  INV_X1    g394(.A(new_n511), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n325), .A2(KEYINPUT5), .ZN(new_n582));
  OAI21_X1  g396(.A(G113), .B1(new_n318), .B2(KEYINPUT5), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n323), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n580), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(G110), .B(G122), .Z(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n588), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n580), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n589), .A2(KEYINPUT6), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT80), .B1(new_n290), .B2(G125), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n281), .A2(new_n196), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n290), .A2(G125), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n593), .B1(new_n596), .B2(KEYINPUT80), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n217), .A2(G224), .ZN(new_n598));
  XOR2_X1   g412(.A(new_n598), .B(KEYINPUT81), .Z(new_n599));
  XNOR2_X1  g413(.A(new_n597), .B(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT6), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n587), .A2(new_n601), .A3(new_n588), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n592), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(G210), .B1(G237), .B2(G902), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT83), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n598), .A2(KEYINPUT7), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n607), .B1(new_n597), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT80), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n594), .B2(new_n595), .ZN(new_n612));
  OAI211_X1 g426(.A(KEYINPUT83), .B(new_n608), .C1(new_n612), .C2(new_n593), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n583), .A2(KEYINPUT82), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n583), .A2(KEYINPUT82), .ZN(new_n615));
  AOI211_X1 g429(.A(new_n614), .B(new_n615), .C1(KEYINPUT5), .C2(new_n330), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n581), .B1(new_n323), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n585), .A2(new_n511), .ZN(new_n618));
  XOR2_X1   g432(.A(new_n588), .B(KEYINPUT8), .Z(new_n619));
  NAND3_X1  g433(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n610), .A2(new_n613), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n597), .A2(new_n609), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n591), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n225), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n604), .A2(new_n606), .A3(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n610), .A2(new_n613), .A3(new_n620), .ZN(new_n626));
  INV_X1    g440(.A(new_n623), .ZN(new_n627));
  AOI21_X1  g441(.A(G902), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n605), .B1(new_n628), .B2(new_n603), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n578), .B(new_n579), .C1(new_n625), .C2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n568), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n378), .A2(new_n487), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(G101), .ZN(G3));
  NAND2_X1  g447(.A1(new_n436), .A2(new_n438), .ZN(new_n634));
  INV_X1    g448(.A(G472), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n635), .B1(new_n367), .B2(new_n225), .ZN(new_n636));
  INV_X1    g450(.A(new_n237), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n350), .A2(new_n358), .A3(new_n362), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n341), .B(KEYINPUT71), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n636), .A2(new_n640), .A3(new_n236), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n474), .B(KEYINPUT33), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n642), .A2(G478), .A3(new_n225), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n476), .A2(new_n481), .A3(new_n479), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n634), .A2(new_n631), .A3(new_n641), .A4(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  AND2_X1   g462(.A1(new_n631), .A2(new_n641), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n484), .B1(new_n480), .B2(new_n482), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT94), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n412), .B(new_n651), .ZN(new_n652));
  OAI211_X1 g466(.A(new_n650), .B(new_n652), .C1(new_n432), .C2(new_n434), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n649), .A2(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT35), .B(G107), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G9));
  NAND3_X1  g471(.A1(new_n436), .A2(new_n438), .A3(new_n486), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n564), .A2(new_n566), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n541), .A2(new_n551), .A3(KEYINPUT79), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n558), .B1(new_n557), .B2(new_n559), .ZN(new_n661));
  OAI21_X1  g475(.A(G469), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n490), .B1(new_n659), .B2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n579), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n606), .B1(new_n604), .B2(new_n624), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n628), .A2(new_n605), .A3(new_n603), .ZN(new_n666));
  AOI211_X1 g480(.A(new_n577), .B(new_n664), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n636), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n364), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n658), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n220), .A2(KEYINPUT36), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n212), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n227), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n235), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT37), .B(G110), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G12));
  INV_X1    g492(.A(G900), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n572), .B1(new_n576), .B2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n653), .A2(new_n680), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n367), .A2(new_n368), .A3(new_n237), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n368), .B1(new_n367), .B2(new_n237), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n377), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n665), .A2(new_n666), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n675), .A2(new_n685), .A3(new_n579), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n681), .A2(new_n684), .A3(new_n663), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  NAND2_X1  g503(.A1(new_n634), .A2(new_n650), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n685), .B(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n690), .A2(new_n693), .A3(new_n664), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n680), .B(KEYINPUT39), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n663), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n675), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n339), .B1(new_n345), .B2(new_n359), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT96), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n635), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n349), .B(new_n703), .C1(new_n702), .C2(new_n701), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n635), .A2(new_n225), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(new_n707), .B(KEYINPUT97), .Z(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n365), .B2(new_n369), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n694), .A2(new_n699), .A3(new_n700), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G143), .ZN(G45));
  NAND3_X1  g526(.A1(new_n684), .A2(new_n663), .A3(new_n687), .ZN(new_n713));
  INV_X1    g527(.A(new_n680), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n430), .A2(new_n407), .ZN(new_n715));
  INV_X1    g529(.A(G475), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n715), .A2(new_n716), .A3(new_n225), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT20), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n431), .A2(new_n413), .A3(new_n225), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n437), .B1(new_n720), .B2(new_n412), .ZN(new_n721));
  INV_X1    g535(.A(new_n438), .ZN(new_n722));
  OAI211_X1 g536(.A(new_n645), .B(new_n714), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n713), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n203), .ZN(G48));
  INV_X1    g539(.A(new_n236), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n534), .A2(new_n536), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n556), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n550), .A2(new_n536), .A3(new_n540), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n225), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(G469), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n491), .A3(new_n564), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n684), .A2(new_n726), .A3(new_n667), .A4(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n645), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n736), .B1(new_n436), .B2(new_n438), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g553(.A(KEYINPUT41), .B(G113), .Z(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G15));
  AND4_X1   g555(.A1(new_n684), .A2(new_n726), .A3(new_n667), .A4(new_n734), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT99), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n743), .A3(new_n654), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT99), .B1(new_n735), .B2(new_n653), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G116), .ZN(G18));
  NOR3_X1   g561(.A1(new_n686), .A2(new_n733), .A3(new_n577), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n487), .A2(new_n748), .A3(new_n684), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G119), .ZN(G21));
  NAND2_X1  g564(.A1(new_n690), .A2(KEYINPUT101), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n340), .B1(new_n357), .B2(KEYINPUT100), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n752), .B1(KEYINPUT100), .B2(new_n357), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n639), .A2(new_n350), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(new_n237), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n669), .A2(new_n755), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n756), .A2(new_n236), .A3(new_n733), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT101), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n634), .A2(new_n758), .A3(new_n650), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n751), .A2(new_n667), .A3(new_n757), .A4(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT102), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n758), .B1(new_n634), .B2(new_n650), .ZN(new_n762));
  AOI211_X1 g576(.A(KEYINPUT101), .B(new_n486), .C1(new_n436), .C2(new_n438), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT102), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n764), .A2(new_n765), .A3(new_n667), .A4(new_n757), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n761), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G122), .ZN(G24));
  AOI21_X1  g582(.A(new_n636), .B1(new_n237), .B2(new_n754), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n686), .A2(new_n733), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n737), .A2(new_n769), .A3(new_n714), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT103), .ZN(new_n772));
  AOI211_X1 g586(.A(new_n736), .B(new_n680), .C1(new_n436), .C2(new_n438), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT103), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n773), .A2(new_n774), .A3(new_n770), .A4(new_n769), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G125), .ZN(G27));
  INV_X1    g591(.A(KEYINPUT42), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n685), .A2(new_n664), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n737), .A2(new_n714), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n559), .A2(KEYINPUT104), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n541), .A2(new_n551), .ZN(new_n782));
  OAI211_X1 g596(.A(G469), .B(new_n781), .C1(new_n782), .C2(KEYINPUT104), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n490), .B1(new_n659), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n684), .A2(new_n726), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n778), .B1(new_n780), .B2(new_n785), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n684), .A2(new_n726), .A3(new_n784), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(KEYINPUT42), .A3(new_n773), .A4(new_n779), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G131), .ZN(G33));
  AND4_X1   g604(.A1(new_n684), .A2(new_n681), .A3(new_n726), .A4(new_n784), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n791), .A2(new_n779), .ZN(new_n792));
  XOR2_X1   g606(.A(KEYINPUT105), .B(G134), .Z(new_n793));
  XNOR2_X1  g607(.A(new_n792), .B(new_n793), .ZN(G36));
  NAND3_X1  g608(.A1(new_n436), .A2(new_n438), .A3(new_n645), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT43), .Z(new_n796));
  OR2_X1    g610(.A1(new_n796), .A2(KEYINPUT106), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(KEYINPUT106), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n797), .A2(new_n670), .A3(new_n675), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(KEYINPUT44), .ZN(new_n800));
  OAI211_X1 g614(.A(KEYINPUT45), .B(new_n781), .C1(new_n782), .C2(KEYINPUT104), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n552), .A2(new_n560), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n801), .B(G469), .C1(KEYINPUT45), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n566), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT46), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n804), .A2(new_n805), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n807), .A2(new_n564), .A3(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(new_n490), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n695), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n779), .B(KEYINPUT107), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n800), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G137), .ZN(G39));
  NOR2_X1   g629(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n810), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT108), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT47), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  MUX2_X1   g635(.A(new_n810), .B(new_n817), .S(new_n821), .Z(new_n822));
  AOI22_X1  g636(.A1(new_n365), .A2(new_n369), .B1(G472), .B2(new_n376), .ZN(new_n823));
  INV_X1    g637(.A(new_n780), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n822), .A2(new_n823), .A3(new_n236), .A4(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(G140), .ZN(G42));
  NAND2_X1  g640(.A1(new_n732), .A2(new_n564), .ZN(new_n827));
  XOR2_X1   g641(.A(new_n827), .B(KEYINPUT49), .Z(new_n828));
  NAND4_X1  g642(.A1(new_n828), .A2(new_n726), .A3(new_n579), .A4(new_n693), .ZN(new_n829));
  OR4_X1    g643(.A1(new_n490), .A2(new_n829), .A3(new_n710), .A4(new_n795), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT109), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n631), .A2(new_n438), .A3(new_n436), .A4(new_n486), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n684), .A2(new_n726), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n646), .B(new_n831), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n831), .B1(new_n632), .B2(new_n646), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AND4_X1   g651(.A1(new_n720), .A2(new_n486), .A3(new_n652), .A4(new_n714), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n684), .A2(new_n838), .A3(new_n663), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n769), .A2(new_n784), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n839), .B1(new_n723), .B2(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n700), .A2(new_n664), .A3(new_n685), .ZN(new_n842));
  AOI22_X1  g656(.A1(new_n841), .A2(new_n842), .B1(new_n791), .B2(new_n779), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n634), .A2(new_n486), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n671), .A2(new_n675), .B1(new_n649), .B2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n837), .A2(new_n789), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n749), .B1(new_n738), .B2(new_n735), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(new_n744), .B2(new_n745), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n767), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT110), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n846), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n658), .A2(new_n823), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n742), .A2(new_n737), .B1(new_n852), .B2(new_n748), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n743), .B1(new_n742), .B2(new_n654), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n735), .A2(KEYINPUT99), .A3(new_n653), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n766), .B2(new_n761), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n789), .A2(new_n843), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n646), .B1(new_n832), .B2(new_n833), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT109), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n845), .A3(new_n834), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT110), .B1(new_n857), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n688), .B1(new_n713), .B2(new_n723), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n864), .B1(new_n775), .B2(new_n772), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n685), .A2(new_n579), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n700), .A2(KEYINPUT111), .A3(new_n714), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT111), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n869), .B1(new_n675), .B2(new_n680), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n868), .A2(new_n784), .A3(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n764), .A2(new_n867), .A3(new_n710), .A4(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT52), .B1(new_n865), .B2(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n865), .A2(KEYINPUT52), .A3(new_n872), .ZN(new_n874));
  OAI22_X1  g688(.A1(new_n851), .A2(new_n863), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT113), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n846), .A2(new_n849), .ZN(new_n880));
  INV_X1    g694(.A(new_n864), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n872), .A2(new_n776), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT52), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT112), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n865), .A2(KEYINPUT52), .A3(new_n872), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n873), .A2(KEYINPUT112), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n880), .A2(new_n887), .A3(KEYINPUT53), .A4(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n874), .A2(new_n873), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n850), .B1(new_n846), .B2(new_n849), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n857), .A2(new_n862), .A3(KEYINPUT110), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI211_X1 g708(.A(new_n879), .B(new_n889), .C1(new_n894), .C2(KEYINPUT53), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT113), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n892), .A2(new_n893), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n897), .A2(new_n876), .A3(new_n888), .A4(new_n887), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n898), .B(KEYINPUT54), .C1(new_n876), .C2(new_n894), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT114), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n890), .A2(new_n896), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n827), .B(KEYINPUT115), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n490), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(new_n904));
  OR3_X1    g718(.A1(new_n822), .A2(KEYINPUT116), .A3(new_n904), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n796), .A2(new_n572), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n906), .A2(new_n726), .A3(new_n769), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n907), .A2(new_n813), .ZN(new_n908));
  OAI21_X1  g722(.A(KEYINPUT116), .B1(new_n822), .B2(new_n904), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n905), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n907), .A2(new_n734), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n911), .A2(KEYINPUT50), .A3(new_n664), .A4(new_n693), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT50), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n907), .A2(new_n664), .A3(new_n734), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n913), .B1(new_n914), .B2(new_n692), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n733), .A2(new_n664), .A3(new_n685), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n906), .A2(new_n917), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n918), .A2(new_n700), .A3(new_n756), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n709), .A2(new_n726), .A3(new_n572), .A4(new_n917), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n921), .A2(new_n634), .A3(new_n645), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n916), .A2(KEYINPUT51), .A3(new_n920), .A4(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(KEYINPUT117), .B1(new_n910), .B2(new_n924), .ZN(new_n925));
  AOI211_X1 g739(.A(new_n919), .B(new_n922), .C1(new_n912), .C2(new_n915), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT117), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n905), .A2(new_n908), .A3(new_n909), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n926), .A2(new_n927), .A3(new_n928), .A4(KEYINPUT51), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n908), .B1(new_n822), .B2(new_n904), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n916), .A2(new_n920), .A3(new_n923), .A4(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT51), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n925), .A2(new_n929), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n890), .A2(new_n896), .A3(new_n899), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(KEYINPUT114), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n918), .A2(new_n833), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT48), .Z(new_n938));
  OR2_X1    g752(.A1(new_n921), .A2(new_n738), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n911), .A2(new_n867), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n938), .A2(new_n569), .A3(new_n939), .A4(new_n940), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT118), .Z(new_n942));
  AND4_X1   g756(.A1(new_n901), .A2(new_n934), .A3(new_n936), .A4(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(G952), .A2(G953), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n830), .B1(new_n943), .B2(new_n944), .ZN(G75));
  AND2_X1   g759(.A1(new_n592), .A2(new_n602), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(new_n600), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT55), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n877), .A2(new_n889), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(G902), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT119), .ZN(new_n951));
  AOI211_X1 g765(.A(KEYINPUT56), .B(new_n948), .C1(new_n951), .C2(new_n606), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n217), .A2(G952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT56), .ZN(new_n954));
  INV_X1    g768(.A(G210), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n954), .B1(new_n950), .B2(new_n955), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n956), .A2(new_n948), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n952), .A2(new_n953), .A3(new_n957), .ZN(G51));
  INV_X1    g772(.A(new_n951), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n959), .A2(new_n803), .ZN(new_n960));
  XOR2_X1   g774(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n961));
  OR2_X1    g775(.A1(new_n961), .A2(new_n565), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n565), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n879), .B1(new_n877), .B2(new_n889), .ZN(new_n964));
  INV_X1    g778(.A(new_n895), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n962), .B(new_n963), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT121), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n966), .A2(new_n967), .A3(new_n730), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n967), .B1(new_n966), .B2(new_n730), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n953), .B1(new_n960), .B2(new_n970), .ZN(G54));
  NAND2_X1  g785(.A1(KEYINPUT58), .A2(G475), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n433), .B1(new_n959), .B2(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n951), .A2(KEYINPUT58), .A3(G475), .A4(new_n715), .ZN(new_n974));
  INV_X1    g788(.A(new_n953), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(G60));
  OR2_X1    g790(.A1(new_n964), .A2(new_n965), .ZN(new_n977));
  INV_X1    g791(.A(new_n642), .ZN(new_n978));
  NAND2_X1  g792(.A1(G478), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT59), .Z(new_n980));
  NOR2_X1   g794(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n953), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n980), .B1(new_n936), .B2(new_n901), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n982), .B1(new_n983), .B2(new_n642), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(KEYINPUT122), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT122), .ZN(new_n986));
  OAI211_X1 g800(.A(new_n986), .B(new_n982), .C1(new_n983), .C2(new_n642), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(G63));
  NAND2_X1  g802(.A1(G217), .A2(G902), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT124), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT60), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n949), .A2(new_n673), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n975), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n223), .B1(new_n949), .B2(new_n991), .ZN(new_n994));
  OAI21_X1  g808(.A(KEYINPUT123), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT61), .ZN(G66));
  AOI21_X1  g810(.A(new_n217), .B1(new_n573), .B2(G224), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n857), .A2(new_n845), .A3(new_n837), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n997), .B1(new_n998), .B2(new_n217), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT125), .ZN(new_n1000));
  INV_X1    g814(.A(G898), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n946), .B1(new_n1001), .B2(G953), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1000), .B(new_n1002), .ZN(G69));
  OAI21_X1  g817(.A(G953), .B1(new_n538), .B2(new_n679), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT126), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n865), .A2(new_n711), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT62), .Z(new_n1007));
  OAI21_X1  g821(.A(new_n738), .B1(new_n634), .B2(new_n486), .ZN(new_n1008));
  INV_X1    g822(.A(new_n697), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n1008), .A2(new_n378), .A3(new_n1009), .A4(new_n779), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n814), .A2(new_n825), .A3(new_n1007), .A4(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n415), .A2(new_n417), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n317), .B(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1011), .A2(new_n217), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n792), .B1(new_n786), .B2(new_n788), .ZN(new_n1016));
  INV_X1    g830(.A(new_n865), .ZN(new_n1017));
  NOR4_X1   g831(.A1(new_n762), .A2(new_n763), .A3(new_n833), .A4(new_n866), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1017), .B1(new_n812), .B2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n814), .A2(new_n825), .A3(new_n1016), .A4(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1013), .B1(new_n1020), .B2(new_n217), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1005), .B1(new_n1015), .B2(new_n1021), .ZN(new_n1022));
  AND2_X1   g836(.A1(new_n1013), .A2(new_n538), .ZN(new_n1023));
  OAI21_X1  g837(.A(G953), .B1(new_n1023), .B2(new_n679), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1022), .A2(new_n1024), .ZN(G72));
  XNOR2_X1  g839(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n706), .B(new_n1026), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1027), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1028), .B1(new_n1011), .B2(new_n998), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n374), .A2(new_n339), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n953), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1028), .B1(new_n1020), .B2(new_n998), .ZN(new_n1032));
  NOR3_X1   g846(.A1(new_n344), .A2(new_n345), .A3(new_n340), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NOR3_X1   g848(.A1(new_n1030), .A2(new_n1027), .A3(new_n1033), .ZN(new_n1035));
  OAI211_X1 g849(.A(new_n898), .B(new_n1035), .C1(new_n876), .C2(new_n894), .ZN(new_n1036));
  AND3_X1   g850(.A1(new_n1031), .A2(new_n1034), .A3(new_n1036), .ZN(G57));
endmodule


