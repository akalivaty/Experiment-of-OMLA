//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 0 0 0 1 0 1 0 1 0 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G119), .ZN(new_n188));
  INV_X1    g002(.A(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G128), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT24), .B(G110), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n194), .B1(new_n189), .B2(G128), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n187), .A2(KEYINPUT23), .A3(G119), .ZN(new_n196));
  INV_X1    g010(.A(G110), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n195), .A2(new_n196), .A3(new_n197), .A4(new_n190), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n193), .A2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(G125), .B(G140), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G125), .ZN(new_n204));
  INV_X1    g018(.A(G125), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G140), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT16), .ZN(new_n207));
  OR3_X1    g021(.A1(new_n205), .A2(KEYINPUT16), .A3(G140), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G146), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n199), .A2(new_n202), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT77), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n199), .A2(KEYINPUT77), .A3(new_n202), .A4(new_n209), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n207), .A2(new_n208), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(new_n201), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(new_n209), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n195), .A2(new_n196), .A3(new_n190), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G110), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n217), .B(new_n219), .C1(new_n191), .C2(new_n192), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G953), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(G221), .A3(G234), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n223), .B(KEYINPUT79), .ZN(new_n224));
  XOR2_X1   g038(.A(KEYINPUT22), .B(G137), .Z(new_n225));
  XNOR2_X1  g039(.A(new_n224), .B(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n221), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT78), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n221), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n214), .A2(KEYINPUT78), .A3(new_n220), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(new_n226), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT80), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT80), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n229), .A2(new_n233), .A3(new_n230), .A4(new_n226), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n227), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT76), .B(G217), .ZN(new_n236));
  INV_X1    g050(.A(G902), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n236), .B1(G234), .B2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(G902), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n237), .B1(new_n221), .B2(new_n226), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n241), .B1(new_n232), .B2(new_n234), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT25), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n238), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AOI211_X1 g058(.A(KEYINPUT25), .B(new_n241), .C1(new_n232), .C2(new_n234), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n240), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n247));
  INV_X1    g061(.A(G116), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT68), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT68), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G116), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n249), .A2(new_n251), .A3(G119), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n248), .A2(G119), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT2), .A2(G113), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  NOR3_X1   g072(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n256), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n247), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT68), .B(G116), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n253), .B1(new_n262), .B2(G119), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT2), .ZN(new_n265));
  INV_X1    g079(.A(G113), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n267), .A2(new_n257), .B1(KEYINPUT2), .B2(G113), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n263), .A2(KEYINPUT69), .A3(new_n268), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n261), .A2(new_n269), .B1(new_n260), .B2(new_n255), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT11), .ZN(new_n271));
  INV_X1    g085(.A(G134), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n271), .B1(new_n272), .B2(G137), .ZN(new_n273));
  INV_X1    g087(.A(G137), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(KEYINPUT11), .A3(G134), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n272), .A2(G137), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G131), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT66), .ZN(new_n279));
  INV_X1    g093(.A(G131), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n273), .A2(new_n275), .A3(new_n280), .A4(new_n276), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n278), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G143), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(G146), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT65), .B1(new_n201), .B2(G143), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT65), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(new_n283), .A3(G146), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n284), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  AND2_X1   g102(.A1(KEYINPUT0), .A2(G128), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n201), .A2(G143), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n283), .A2(G146), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT64), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT0), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n293), .A2(new_n294), .A3(new_n187), .ZN(new_n295));
  OAI21_X1  g109(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n288), .A2(new_n289), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n277), .A2(KEYINPUT66), .A3(G131), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n282), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT1), .ZN(new_n301));
  OAI21_X1  g115(.A(G128), .B1(new_n284), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n290), .A2(new_n291), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n187), .A2(KEYINPUT1), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n286), .B1(new_n283), .B2(G146), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n201), .A2(KEYINPUT65), .A3(G143), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n290), .B(new_n305), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n276), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n272), .A2(G137), .ZN(new_n311));
  OAI21_X1  g125(.A(G131), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n281), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n270), .A2(new_n300), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT28), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n314), .A2(KEYINPUT70), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n300), .A2(new_n313), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n261), .A2(new_n269), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n255), .A2(new_n260), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT70), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n270), .A2(new_n324), .A3(new_n300), .A4(new_n313), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n318), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n317), .B1(new_n326), .B2(KEYINPUT28), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT26), .B(G101), .ZN(new_n329));
  NOR2_X1   g143(.A1(G237), .A2(G953), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G210), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n329), .B(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n332), .B(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n318), .A2(new_n325), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT30), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n300), .A2(new_n337), .A3(new_n313), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n337), .B1(new_n300), .B2(new_n313), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n322), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n336), .A2(KEYINPUT31), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT31), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n318), .A2(new_n325), .A3(new_n335), .ZN(new_n343));
  INV_X1    g157(.A(new_n339), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n300), .A2(new_n313), .A3(new_n337), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n270), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n342), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n328), .A2(new_n334), .B1(new_n341), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(G472), .A2(G902), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT72), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT32), .ZN(new_n352));
  AOI21_X1  g166(.A(KEYINPUT31), .B1(new_n336), .B2(new_n340), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n343), .A2(new_n346), .A3(new_n342), .ZN(new_n354));
  OAI22_X1  g168(.A1(new_n353), .A2(new_n354), .B1(new_n327), .B2(new_n335), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT72), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n356), .A3(new_n349), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n351), .A2(new_n352), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n348), .A2(new_n350), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(KEYINPUT32), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n326), .A2(KEYINPUT28), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(new_n316), .A3(new_n335), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n340), .A2(new_n318), .A3(new_n325), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT29), .B1(new_n364), .B2(new_n334), .ZN(new_n365));
  AOI21_X1  g179(.A(G902), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT73), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n323), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n319), .A2(KEYINPUT73), .A3(new_n322), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n368), .A2(new_n318), .A3(new_n325), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT28), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n316), .A2(KEYINPUT29), .A3(new_n335), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT74), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT74), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n375), .A3(new_n372), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n366), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G472), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT75), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n377), .A2(KEYINPUT75), .A3(G472), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n246), .B1(new_n361), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G104), .ZN(new_n384));
  OAI211_X1 g198(.A(KEYINPUT81), .B(KEYINPUT3), .C1(new_n384), .C2(G107), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT3), .ZN(new_n386));
  INV_X1    g200(.A(G107), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n387), .A3(G104), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n384), .A2(G107), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n385), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n387), .A2(G104), .ZN(new_n391));
  AOI21_X1  g205(.A(KEYINPUT81), .B1(new_n391), .B2(KEYINPUT3), .ZN(new_n392));
  OAI21_X1  g206(.A(G101), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT82), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT82), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n395), .B(G101), .C1(new_n390), .C2(new_n392), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n388), .A2(new_n389), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT81), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n384), .A2(G107), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n398), .B1(new_n399), .B2(new_n386), .ZN(new_n400));
  INV_X1    g214(.A(G101), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n397), .A2(new_n400), .A3(new_n401), .A4(new_n385), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n394), .A2(KEYINPUT4), .A3(new_n396), .A4(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT4), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n404), .B(G101), .C1(new_n390), .C2(new_n392), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(new_n322), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT87), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n391), .A2(new_n389), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G101), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n402), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n263), .A2(KEYINPUT5), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT5), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n266), .B1(new_n253), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  AND4_X1   g228(.A1(new_n407), .A2(new_n410), .A3(new_n320), .A4(new_n414), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n261), .A2(new_n269), .B1(new_n411), .B2(new_n413), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n407), .B1(new_n416), .B2(new_n410), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n406), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(G110), .B(G122), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n419), .B(new_n406), .C1(new_n415), .C2(new_n417), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n421), .A2(KEYINPUT6), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT6), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n418), .A2(new_n424), .A3(new_n420), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n309), .A2(G125), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n288), .A2(new_n289), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n292), .A2(new_n297), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n205), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n222), .A2(G224), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(KEYINPUT88), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n430), .B(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n423), .A2(new_n425), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G210), .B1(G237), .B2(G902), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n320), .A2(new_n414), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n402), .A2(new_n409), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n416), .A2(new_n410), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n419), .B(KEYINPUT8), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT89), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n432), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n443), .B1(new_n426), .B2(new_n429), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n432), .A2(KEYINPUT7), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n445), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n443), .B(new_n447), .C1(new_n426), .C2(new_n429), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n440), .A2(new_n441), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n422), .ZN(new_n450));
  AOI21_X1  g264(.A(KEYINPUT90), .B1(new_n450), .B2(new_n237), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT90), .ZN(new_n452));
  AOI211_X1 g266(.A(new_n452), .B(G902), .C1(new_n449), .C2(new_n422), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n434), .B(new_n435), .C1(new_n451), .C2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n435), .B(KEYINPUT92), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n434), .B1(new_n451), .B2(new_n453), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n457), .B1(new_n458), .B2(KEYINPUT91), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT91), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n434), .B(new_n460), .C1(new_n451), .C2(new_n453), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n455), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G469), .ZN(new_n463));
  XNOR2_X1  g277(.A(G110), .B(G140), .ZN(new_n464));
  INV_X1    g278(.A(G227), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(G953), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n464), .B(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n282), .A2(new_n299), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n405), .A2(new_n298), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n396), .A2(KEYINPUT4), .A3(new_n402), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n397), .A2(new_n400), .A3(new_n385), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n395), .B1(new_n473), .B2(G101), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n471), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n410), .A2(KEYINPUT10), .A3(new_n309), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n290), .B1(new_n306), .B2(new_n307), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT84), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n479), .B1(new_n290), .B2(KEYINPUT1), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n479), .B(KEYINPUT1), .C1(new_n283), .C2(G146), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G128), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n478), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n308), .A2(KEYINPUT83), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT83), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n288), .A2(new_n485), .A3(new_n305), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT10), .B1(new_n487), .B2(new_n410), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n470), .B1(new_n477), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT86), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n487), .A2(new_n410), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT10), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(new_n475), .A3(new_n476), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(KEYINPUT86), .A3(new_n470), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n494), .A2(new_n469), .A3(new_n475), .A4(new_n476), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n468), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n468), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n437), .A2(new_n304), .A3(new_n308), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n469), .B1(new_n492), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT12), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT85), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n503), .B1(new_n469), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  OR2_X1    g320(.A1(new_n502), .A2(new_n505), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n500), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n463), .B(new_n237), .C1(new_n499), .C2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n500), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n495), .A2(KEYINPUT86), .A3(new_n470), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT86), .B1(new_n495), .B2(new_n470), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n492), .A2(new_n501), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n514), .A2(new_n470), .A3(new_n505), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n502), .A2(new_n505), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n498), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n467), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n513), .A2(new_n518), .A3(G469), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n463), .A2(new_n237), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n509), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT9), .B(G234), .ZN(new_n523));
  OAI21_X1  g337(.A(G221), .B1(new_n523), .B2(G902), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(G214), .B1(G237), .B2(G902), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n462), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n330), .A2(G143), .A3(G214), .ZN(new_n529));
  AOI21_X1  g343(.A(G143), .B1(new_n330), .B2(G214), .ZN(new_n530));
  OAI21_X1  g344(.A(G131), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n532));
  INV_X1    g346(.A(G237), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n222), .A3(G214), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n283), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n330), .A2(G143), .A3(G214), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n280), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n531), .A2(new_n532), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT94), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n217), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n531), .A2(new_n537), .A3(KEYINPUT94), .A4(new_n532), .ZN(new_n542));
  OR2_X1    g356(.A1(new_n531), .A2(new_n532), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n540), .A2(new_n541), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(G113), .B(G122), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(new_n384), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n529), .A2(new_n530), .ZN(new_n547));
  NAND2_X1  g361(.A1(KEYINPUT18), .A2(G131), .ZN(new_n548));
  OR2_X1    g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n204), .A2(new_n206), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(G146), .ZN(new_n551));
  AOI22_X1  g365(.A1(new_n547), .A2(new_n548), .B1(new_n202), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n544), .A2(new_n546), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n546), .B1(new_n544), .B2(new_n553), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n237), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(G475), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT19), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n550), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n200), .A2(KEYINPUT19), .ZN(new_n561));
  AOI21_X1  g375(.A(G146), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n209), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n531), .A2(new_n537), .ZN(new_n565));
  AOI22_X1  g379(.A1(new_n564), .A2(new_n565), .B1(new_n549), .B2(new_n552), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT93), .B1(new_n566), .B2(new_n546), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n560), .A2(new_n561), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n565), .B(new_n209), .C1(new_n568), .C2(G146), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n553), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT93), .ZN(new_n571));
  INV_X1    g385(.A(new_n546), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n554), .A2(new_n567), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT20), .ZN(new_n575));
  NOR2_X1   g389(.A1(G475), .A2(G902), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n575), .B1(new_n574), .B2(new_n576), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n558), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n187), .A2(G143), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT13), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n272), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(G128), .B(G143), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(KEYINPUT95), .B(G122), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(G116), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n249), .A2(new_n251), .A3(G122), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n586), .A2(new_n387), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n387), .B1(new_n586), .B2(new_n587), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n584), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n587), .A2(KEYINPUT14), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n587), .A2(KEYINPUT14), .B1(new_n585), .B2(G116), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n387), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n583), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT96), .B(G134), .ZN(new_n595));
  OR2_X1    g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n586), .A2(new_n387), .A3(new_n587), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n594), .A2(new_n595), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n590), .B1(new_n593), .B2(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n236), .A2(new_n523), .A3(G953), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n590), .B(new_n601), .C1(new_n593), .C2(new_n599), .ZN(new_n604));
  AOI21_X1  g418(.A(G902), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(G478), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n606), .A2(KEYINPUT15), .ZN(new_n607));
  XOR2_X1   g421(.A(new_n605), .B(new_n607), .Z(new_n608));
  OR2_X1    g422(.A1(new_n579), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n222), .A2(G952), .ZN(new_n610));
  INV_X1    g424(.A(G234), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n610), .B1(new_n611), .B2(new_n533), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  AOI211_X1 g427(.A(new_n237), .B(new_n222), .C1(G234), .C2(G237), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT21), .B(G898), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n609), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n383), .A2(new_n528), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  INV_X1    g433(.A(new_n525), .ZN(new_n620));
  OAI21_X1  g434(.A(G472), .B1(new_n348), .B2(G902), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n621), .A2(new_n351), .A3(new_n357), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n622), .A2(new_n246), .ZN(new_n623));
  INV_X1    g437(.A(new_n435), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n458), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n527), .B1(new_n625), .B2(new_n454), .ZN(new_n626));
  AND3_X1   g440(.A1(new_n620), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n616), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n603), .A2(new_n604), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n600), .A2(KEYINPUT97), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(KEYINPUT33), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n603), .A2(new_n630), .A3(KEYINPUT33), .A4(new_n604), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n606), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n605), .A2(new_n606), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n606), .A2(new_n237), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n579), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n627), .A2(new_n628), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT34), .B(G104), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  OAI211_X1 g458(.A(new_n608), .B(new_n558), .C1(new_n578), .C2(new_n577), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n627), .A2(new_n628), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT35), .B(G107), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  NAND2_X1  g463(.A1(new_n229), .A2(new_n230), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n226), .A2(KEYINPUT36), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n650), .A2(new_n651), .ZN(new_n653));
  OR2_X1    g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n239), .ZN(new_n655));
  OAI22_X1  g469(.A1(new_n244), .A2(new_n245), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n617), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n622), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n462), .A2(new_n527), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n658), .A2(new_n659), .A3(new_n620), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT37), .B(G110), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G12));
  AND3_X1   g476(.A1(new_n377), .A2(KEYINPUT75), .A3(G472), .ZN(new_n663));
  AOI21_X1  g477(.A(KEYINPUT75), .B1(new_n377), .B2(G472), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n358), .B(new_n360), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n626), .A2(new_n656), .ZN(new_n666));
  INV_X1    g480(.A(G900), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n614), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n645), .B1(new_n612), .B2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n665), .A2(new_n666), .A3(new_n620), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G128), .ZN(G30));
  NAND2_X1  g485(.A1(new_n668), .A2(new_n612), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(KEYINPUT39), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n620), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT99), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT99), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n674), .B(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT40), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n462), .B(KEYINPUT38), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n579), .A2(new_n608), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n526), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n238), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n232), .A2(new_n234), .ZN(new_n686));
  INV_X1    g500(.A(new_n241), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n685), .B1(new_n688), .B2(KEYINPUT25), .ZN(new_n689));
  INV_X1    g503(.A(new_n245), .ZN(new_n690));
  INV_X1    g504(.A(new_n654), .ZN(new_n691));
  AOI22_X1  g505(.A1(new_n689), .A2(new_n690), .B1(new_n239), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n343), .A2(new_n346), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n370), .A2(new_n334), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n694), .B1(new_n695), .B2(KEYINPUT98), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n696), .B1(KEYINPUT98), .B2(new_n695), .ZN(new_n697));
  OAI21_X1  g511(.A(G472), .B1(new_n697), .B2(G902), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n358), .A3(new_n360), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n684), .A2(new_n692), .A3(new_n699), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n676), .A2(new_n680), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n283), .ZN(G45));
  NAND3_X1  g516(.A1(new_n579), .A2(new_n639), .A3(new_n672), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT100), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT100), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n579), .A2(new_n639), .A3(new_n705), .A4(new_n672), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n665), .A2(new_n666), .A3(new_n620), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  NAND2_X1  g523(.A1(new_n625), .A2(new_n454), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n526), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n498), .B1(new_n511), .B2(new_n512), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n508), .B1(new_n712), .B2(new_n467), .ZN(new_n713));
  OAI21_X1  g527(.A(G469), .B1(new_n713), .B2(G902), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n524), .A3(new_n509), .ZN(new_n715));
  NOR4_X1   g529(.A1(new_n711), .A2(new_n715), .A3(new_n616), .A4(new_n640), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n383), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XOR2_X1   g532(.A(new_n718), .B(KEYINPUT101), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n717), .B(new_n719), .ZN(G15));
  NAND2_X1  g534(.A1(new_n646), .A2(new_n628), .ZN(new_n721));
  NOR3_X1   g535(.A1(new_n711), .A2(new_n721), .A3(new_n715), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n383), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT102), .B(G116), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G18));
  NOR2_X1   g539(.A1(new_n711), .A2(new_n715), .ZN(new_n726));
  INV_X1    g540(.A(new_n657), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n665), .A3(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT103), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n657), .B1(new_n361), .B2(new_n382), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(KEYINPUT103), .A3(new_n726), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G119), .ZN(G21));
  INV_X1    g548(.A(KEYINPUT104), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n317), .B1(new_n370), .B2(KEYINPUT28), .ZN(new_n736));
  OAI22_X1  g550(.A1(new_n353), .A2(new_n354), .B1(new_n736), .B2(new_n335), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n349), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n621), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n739), .A2(new_n246), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n714), .A2(new_n524), .A3(new_n509), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n741), .A3(new_n628), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n626), .A2(new_n682), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n735), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n626), .A2(new_n682), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n739), .A2(new_n246), .A3(new_n616), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n745), .A2(new_n746), .A3(KEYINPUT104), .A4(new_n741), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G122), .ZN(G24));
  OAI21_X1  g563(.A(KEYINPUT105), .B1(new_n692), .B2(new_n739), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT105), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n656), .A2(new_n751), .A3(new_n621), .A4(new_n738), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n707), .A3(new_n726), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G125), .ZN(G27));
  NAND2_X1  g569(.A1(new_n458), .A2(KEYINPUT91), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n461), .A3(new_n456), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT106), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n519), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n513), .A2(new_n518), .A3(KEYINPUT106), .A4(G469), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n509), .A2(new_n521), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n524), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n527), .ZN(new_n763));
  AND4_X1   g577(.A1(new_n454), .A2(new_n757), .A3(new_n761), .A4(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n246), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n764), .A2(new_n665), .A3(new_n765), .A4(new_n707), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT42), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n359), .B(new_n352), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n246), .B1(new_n382), .B2(new_n768), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n704), .A2(KEYINPUT42), .A3(new_n706), .ZN(new_n770));
  AND4_X1   g584(.A1(new_n462), .A2(new_n770), .A3(new_n761), .A4(new_n763), .ZN(new_n771));
  AOI22_X1  g585(.A1(new_n766), .A2(new_n767), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  XOR2_X1   g586(.A(KEYINPUT107), .B(G131), .Z(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(G33));
  NAND4_X1  g588(.A1(new_n764), .A2(new_n665), .A3(new_n765), .A4(new_n669), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G134), .ZN(G36));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n777));
  INV_X1    g591(.A(new_n513), .ZN(new_n778));
  INV_X1    g592(.A(new_n518), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n777), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n513), .A2(new_n518), .A3(KEYINPUT45), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(G469), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(KEYINPUT46), .A3(new_n521), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n783), .A2(KEYINPUT108), .A3(new_n509), .ZN(new_n784));
  INV_X1    g598(.A(new_n782), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n520), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n784), .B1(KEYINPUT46), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT108), .B1(new_n783), .B2(new_n509), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n524), .B(new_n673), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n791));
  XNOR2_X1  g605(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n792));
  INV_X1    g606(.A(new_n633), .ZN(new_n793));
  AOI22_X1  g607(.A1(KEYINPUT33), .A2(new_n630), .B1(new_n603), .B2(new_n604), .ZN(new_n794));
  OAI21_X1  g608(.A(G478), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n636), .B1(new_n605), .B2(new_n606), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n579), .A2(new_n797), .ZN(new_n798));
  MUX2_X1   g612(.A(new_n791), .B(new_n792), .S(new_n798), .Z(new_n799));
  NAND4_X1  g613(.A1(new_n799), .A2(KEYINPUT44), .A3(new_n622), .A4(new_n656), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT110), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n462), .A2(new_n526), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n799), .A2(new_n622), .A3(new_n656), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT44), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n790), .A2(new_n802), .A3(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G137), .ZN(G39));
  OAI21_X1  g622(.A(new_n524), .B1(new_n787), .B2(new_n788), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT47), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(KEYINPUT111), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n810), .A2(KEYINPUT111), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n809), .B1(new_n813), .B2(new_n811), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n707), .A2(new_n246), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n665), .A2(new_n803), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n812), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G140), .ZN(G42));
  NAND2_X1  g632(.A1(new_n714), .A2(new_n509), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n819), .A2(KEYINPUT49), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n765), .A2(new_n763), .A3(new_n798), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n819), .A2(KEYINPUT49), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n820), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n699), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n681), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n383), .B1(new_n716), .B2(new_n722), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT103), .B1(new_n731), .B2(new_n726), .ZN(new_n827));
  AND4_X1   g641(.A1(KEYINPUT103), .A2(new_n726), .A3(new_n665), .A4(new_n727), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n748), .B(new_n826), .C1(new_n827), .C2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n616), .B1(new_n645), .B2(new_n640), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n659), .A2(new_n620), .A3(new_n623), .A4(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n659), .A2(new_n617), .A3(new_n620), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n665), .A2(new_n765), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n831), .B(new_n660), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  AND4_X1   g649(.A1(new_n524), .A2(new_n626), .A3(new_n672), .A4(new_n682), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(new_n692), .A3(new_n699), .A4(new_n761), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n837), .A2(new_n754), .A3(new_n670), .A4(new_n708), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n711), .A2(new_n525), .A3(new_n692), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n841), .B(new_n665), .C1(new_n669), .C2(new_n707), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(KEYINPUT52), .A3(new_n754), .A4(new_n837), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n803), .ZN(new_n845));
  INV_X1    g659(.A(new_n609), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n656), .A3(new_n672), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n847), .A2(new_n525), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n845), .A2(new_n848), .A3(new_n665), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n753), .A2(new_n764), .A3(new_n707), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n775), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n772), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n835), .A2(new_n844), .A3(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT53), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n618), .A2(KEYINPUT53), .A3(new_n660), .A4(new_n831), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n857), .A2(new_n772), .A3(new_n851), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT112), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n829), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n733), .A2(KEYINPUT112), .A3(new_n748), .A4(new_n826), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n844), .A2(new_n858), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n855), .A2(new_n856), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n853), .B(new_n854), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n864), .B1(KEYINPUT54), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT51), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n799), .A2(new_n613), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(new_n740), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n869), .A2(new_n526), .A3(new_n715), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n681), .ZN(new_n871));
  XOR2_X1   g685(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n803), .A2(new_n715), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n868), .A2(new_n874), .A3(new_n753), .ZN(new_n875));
  NOR2_X1   g689(.A1(KEYINPUT114), .A2(KEYINPUT50), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n870), .A2(new_n681), .A3(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n874), .A2(new_n824), .A3(new_n765), .A4(new_n613), .ZN(new_n878));
  OR3_X1    g692(.A1(new_n878), .A2(new_n579), .A3(new_n639), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n873), .A2(new_n875), .A3(new_n877), .A4(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n868), .A2(new_n740), .A3(new_n845), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n812), .A2(new_n814), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n714), .A2(new_n762), .A3(new_n509), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n883), .B(KEYINPUT113), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n881), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n867), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT115), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n888));
  OR3_X1    g702(.A1(new_n880), .A2(new_n888), .A3(new_n867), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n868), .A2(new_n874), .A3(new_n769), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT48), .Z(new_n891));
  NAND3_X1  g705(.A1(new_n868), .A2(new_n726), .A3(new_n740), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n610), .B(new_n892), .C1(new_n878), .C2(new_n640), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  AND4_X1   g708(.A1(new_n866), .A2(new_n887), .A3(new_n889), .A4(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(G952), .A2(G953), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n825), .B1(new_n895), .B2(new_n896), .ZN(G75));
  NOR4_X1   g711(.A1(new_n829), .A2(new_n772), .A3(new_n834), .A4(new_n851), .ZN(new_n898));
  AOI21_X1  g712(.A(KEYINPUT53), .B1(new_n898), .B2(new_n844), .ZN(new_n899));
  AND4_X1   g713(.A1(new_n844), .A2(new_n858), .A3(new_n860), .A4(new_n861), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(new_n237), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT56), .B1(new_n902), .B2(G210), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n423), .A2(new_n425), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(new_n433), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT55), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n222), .A2(G952), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n901), .A2(new_n237), .A3(new_n457), .ZN(new_n910));
  XNOR2_X1  g724(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n909), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n907), .A2(new_n913), .ZN(G51));
  OAI21_X1  g728(.A(KEYINPUT54), .B1(new_n899), .B2(new_n900), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n915), .A2(KEYINPUT117), .A3(new_n863), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n855), .A2(new_n862), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT117), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n917), .A2(new_n918), .A3(KEYINPUT54), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n520), .B(KEYINPUT57), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(KEYINPUT118), .ZN(new_n922));
  INV_X1    g736(.A(new_n713), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT118), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n916), .A2(new_n924), .A3(new_n919), .A4(new_n920), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n902), .A2(new_n785), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n908), .B1(new_n926), .B2(new_n927), .ZN(G54));
  NAND2_X1  g742(.A1(KEYINPUT58), .A2(G475), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT119), .Z(new_n930));
  NAND3_X1  g744(.A1(new_n902), .A2(new_n574), .A3(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n931), .A2(KEYINPUT120), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(KEYINPUT120), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n574), .B1(new_n902), .B2(new_n930), .ZN(new_n934));
  NOR4_X1   g748(.A1(new_n932), .A2(new_n933), .A3(new_n908), .A4(new_n934), .ZN(G60));
  NOR2_X1   g749(.A1(new_n793), .A2(new_n794), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  XNOR2_X1  g751(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n637), .B(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n937), .B1(new_n866), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n937), .A2(new_n939), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n916), .A2(new_n919), .A3(new_n941), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n940), .A2(new_n909), .A3(new_n942), .ZN(G63));
  NAND2_X1  g757(.A1(G217), .A2(G902), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT60), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n917), .A2(new_n691), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n909), .ZN(new_n948));
  OAI21_X1  g762(.A(KEYINPUT61), .B1(new_n948), .B2(KEYINPUT122), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n901), .A2(new_n945), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n909), .B(new_n947), .C1(new_n950), .C2(new_n235), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n949), .B(new_n951), .ZN(G66));
  INV_X1    g766(.A(new_n615), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n222), .B1(new_n953), .B2(G224), .ZN(new_n954));
  INV_X1    g768(.A(new_n835), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n954), .B1(new_n955), .B2(new_n222), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n904), .B1(G898), .B2(new_n222), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n956), .B(new_n957), .Z(G69));
  OAI21_X1  g772(.A(G953), .B1(new_n465), .B2(new_n667), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT124), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n344), .A2(new_n345), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(new_n568), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(G900), .B2(G953), .ZN(new_n963));
  INV_X1    g777(.A(new_n775), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n772), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT126), .Z(new_n966));
  NAND3_X1  g780(.A1(new_n790), .A2(new_n745), .A3(new_n769), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n817), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n842), .A2(new_n754), .ZN(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(KEYINPUT125), .B1(new_n807), .B2(new_n970), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n807), .A2(KEYINPUT125), .A3(new_n970), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n966), .B(new_n968), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n963), .B1(new_n973), .B2(G953), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n383), .B(new_n845), .C1(new_n641), .C2(new_n646), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n675), .A2(new_n975), .ZN(new_n976));
  OR2_X1    g790(.A1(new_n976), .A2(KEYINPUT123), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(KEYINPUT123), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n977), .A2(new_n817), .A3(new_n807), .A4(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT62), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(new_n701), .B2(new_n969), .ZN(new_n981));
  OR2_X1    g795(.A1(new_n680), .A2(new_n700), .ZN(new_n982));
  OAI211_X1 g796(.A(KEYINPUT62), .B(new_n970), .C1(new_n982), .C2(new_n676), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n979), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n962), .B1(new_n984), .B2(G953), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n974), .A2(new_n985), .A3(KEYINPUT127), .ZN(new_n986));
  AOI21_X1  g800(.A(KEYINPUT127), .B1(new_n974), .B2(new_n985), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n960), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OR2_X1    g802(.A1(new_n987), .A2(new_n960), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(G72));
  AND2_X1   g804(.A1(new_n984), .A2(new_n835), .ZN(new_n991));
  NAND2_X1  g805(.A1(G472), .A2(G902), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT63), .Z(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  OAI211_X1 g808(.A(new_n335), .B(new_n364), .C1(new_n991), .C2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n364), .A2(new_n334), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n994), .B1(new_n694), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n908), .B1(new_n865), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n993), .B1(new_n973), .B2(new_n955), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n364), .A2(new_n335), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(G57));
endmodule


