

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590;

  XNOR2_X1 U327 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U328 ( .A(n441), .B(n440), .Z(n295) );
  NOR2_X1 U329 ( .A1(n529), .A2(n522), .ZN(n392) );
  INV_X1 U330 ( .A(KEYINPUT72), .ZN(n434) );
  XNOR2_X1 U331 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U332 ( .A(n319), .B(n430), .ZN(n320) );
  XNOR2_X1 U333 ( .A(n442), .B(n295), .ZN(n443) );
  XNOR2_X1 U334 ( .A(n467), .B(n466), .ZN(n545) );
  XNOR2_X1 U335 ( .A(n321), .B(n320), .ZN(n329) );
  XNOR2_X1 U336 ( .A(n444), .B(n443), .ZN(n448) );
  NOR2_X1 U337 ( .A1(n516), .A2(n485), .ZN(n449) );
  NOR2_X1 U338 ( .A1(n530), .A2(n474), .ZN(n569) );
  NOR2_X1 U339 ( .A1(n515), .A2(n507), .ZN(n512) );
  XOR2_X1 U340 ( .A(n472), .B(KEYINPUT28), .Z(n504) );
  XNOR2_X1 U341 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U342 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U343 ( .A(n478), .B(n477), .ZN(G1351GAT) );
  XNOR2_X1 U344 ( .A(n453), .B(n452), .ZN(G1330GAT) );
  XOR2_X1 U345 ( .A(G155GAT), .B(G211GAT), .Z(n297) );
  XNOR2_X1 U346 ( .A(G127GAT), .B(G183GAT), .ZN(n296) );
  XNOR2_X1 U347 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U348 ( .A(n298), .B(G78GAT), .Z(n300) );
  XOR2_X1 U349 ( .A(G15GAT), .B(G1GAT), .Z(n420) );
  XNOR2_X1 U350 ( .A(G22GAT), .B(n420), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n300), .B(n299), .ZN(n305) );
  XNOR2_X1 U352 ( .A(G71GAT), .B(G57GAT), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n301), .B(KEYINPUT13), .ZN(n446) );
  XOR2_X1 U354 ( .A(G64GAT), .B(n446), .Z(n303) );
  NAND2_X1 U355 ( .A1(G231GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U356 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U357 ( .A(n305), .B(n304), .Z(n313) );
  XOR2_X1 U358 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n307) );
  XNOR2_X1 U359 ( .A(KEYINPUT79), .B(KEYINPUT78), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U361 ( .A(KEYINPUT12), .B(KEYINPUT77), .Z(n309) );
  XNOR2_X1 U362 ( .A(G8GAT), .B(KEYINPUT76), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U364 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n313), .B(n312), .ZN(n584) );
  XOR2_X1 U366 ( .A(G78GAT), .B(G148GAT), .Z(n315) );
  XNOR2_X1 U367 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n315), .B(n314), .ZN(n437) );
  XOR2_X1 U369 ( .A(n437), .B(KEYINPUT85), .Z(n317) );
  NAND2_X1 U370 ( .A1(G228GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n321) );
  XNOR2_X1 U372 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n318) );
  XNOR2_X1 U373 ( .A(n318), .B(KEYINPUT2), .ZN(n368) );
  XOR2_X1 U374 ( .A(G50GAT), .B(G162GAT), .Z(n399) );
  XOR2_X1 U375 ( .A(n368), .B(n399), .Z(n319) );
  XOR2_X1 U376 ( .A(G141GAT), .B(G22GAT), .Z(n430) );
  XOR2_X1 U377 ( .A(KEYINPUT21), .B(G218GAT), .Z(n323) );
  XNOR2_X1 U378 ( .A(KEYINPUT84), .B(G211GAT), .ZN(n322) );
  XNOR2_X1 U379 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U380 ( .A(G197GAT), .B(n324), .ZN(n359) );
  XOR2_X1 U381 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n326) );
  XNOR2_X1 U382 ( .A(KEYINPUT22), .B(G204GAT), .ZN(n325) );
  XNOR2_X1 U383 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U384 ( .A(n359), .B(n327), .Z(n328) );
  XNOR2_X1 U385 ( .A(n329), .B(n328), .ZN(n472) );
  INV_X1 U386 ( .A(KEYINPUT94), .ZN(n362) );
  XOR2_X1 U387 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n331) );
  XNOR2_X1 U388 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U390 ( .A(n332), .B(G127GAT), .Z(n334) );
  XNOR2_X1 U391 ( .A(G113GAT), .B(G120GAT), .ZN(n333) );
  XNOR2_X1 U392 ( .A(n334), .B(n333), .ZN(n379) );
  XOR2_X1 U393 ( .A(G71GAT), .B(G15GAT), .Z(n336) );
  XNOR2_X1 U394 ( .A(G169GAT), .B(G43GAT), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U396 ( .A(G99GAT), .B(G190GAT), .Z(n338) );
  XNOR2_X1 U397 ( .A(KEYINPUT20), .B(G176GAT), .ZN(n337) );
  XNOR2_X1 U398 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U399 ( .A(n340), .B(n339), .Z(n342) );
  NAND2_X1 U400 ( .A1(G227GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U402 ( .A(n379), .B(n343), .ZN(n347) );
  XOR2_X1 U403 ( .A(KEYINPUT18), .B(KEYINPUT83), .Z(n345) );
  XNOR2_X1 U404 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n344) );
  XNOR2_X1 U405 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U406 ( .A(KEYINPUT19), .B(n346), .Z(n358) );
  XOR2_X1 U407 ( .A(n347), .B(n358), .Z(n530) );
  INV_X1 U408 ( .A(n530), .ZN(n522) );
  XOR2_X1 U409 ( .A(G64GAT), .B(G92GAT), .Z(n349) );
  XNOR2_X1 U410 ( .A(G176GAT), .B(G204GAT), .ZN(n348) );
  XNOR2_X1 U411 ( .A(n349), .B(n348), .ZN(n445) );
  XOR2_X1 U412 ( .A(G169GAT), .B(G8GAT), .Z(n418) );
  XOR2_X1 U413 ( .A(n445), .B(n418), .Z(n351) );
  NAND2_X1 U414 ( .A1(G226GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U415 ( .A(n351), .B(n350), .ZN(n353) );
  INV_X1 U416 ( .A(KEYINPUT91), .ZN(n352) );
  XNOR2_X1 U417 ( .A(n353), .B(n352), .ZN(n356) );
  XNOR2_X1 U418 ( .A(G36GAT), .B(G190GAT), .ZN(n354) );
  XNOR2_X1 U419 ( .A(n354), .B(KEYINPUT75), .ZN(n407) );
  XNOR2_X1 U420 ( .A(n407), .B(KEYINPUT92), .ZN(n355) );
  XNOR2_X1 U421 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U422 ( .A(n358), .B(n357), .ZN(n360) );
  XOR2_X1 U423 ( .A(n360), .B(n359), .Z(n500) );
  INV_X1 U424 ( .A(n500), .ZN(n519) );
  NAND2_X1 U425 ( .A1(n522), .A2(n519), .ZN(n361) );
  XNOR2_X1 U426 ( .A(n362), .B(n361), .ZN(n363) );
  NOR2_X1 U427 ( .A1(n472), .A2(n363), .ZN(n364) );
  XOR2_X1 U428 ( .A(KEYINPUT25), .B(n364), .Z(n391) );
  XOR2_X1 U429 ( .A(KEYINPUT93), .B(KEYINPUT26), .Z(n366) );
  NAND2_X1 U430 ( .A1(n472), .A2(n530), .ZN(n365) );
  XNOR2_X1 U431 ( .A(n366), .B(n365), .ZN(n574) );
  XOR2_X1 U432 ( .A(KEYINPUT27), .B(n500), .Z(n389) );
  INV_X1 U433 ( .A(n389), .ZN(n367) );
  NOR2_X1 U434 ( .A1(n574), .A2(n367), .ZN(n546) );
  XNOR2_X1 U435 ( .A(n368), .B(KEYINPUT87), .ZN(n369) );
  XNOR2_X1 U436 ( .A(n369), .B(KEYINPUT89), .ZN(n373) );
  XOR2_X1 U437 ( .A(KEYINPUT88), .B(KEYINPUT5), .Z(n371) );
  XNOR2_X1 U438 ( .A(KEYINPUT6), .B(KEYINPUT90), .ZN(n370) );
  XNOR2_X1 U439 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U440 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U441 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n375) );
  XNOR2_X1 U442 ( .A(G1GAT), .B(KEYINPUT86), .ZN(n374) );
  XNOR2_X1 U443 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U444 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U445 ( .A(n379), .B(n378), .ZN(n387) );
  NAND2_X1 U446 ( .A1(G225GAT), .A2(G233GAT), .ZN(n385) );
  XOR2_X1 U447 ( .A(G57GAT), .B(G148GAT), .Z(n381) );
  XNOR2_X1 U448 ( .A(G29GAT), .B(G141GAT), .ZN(n380) );
  XNOR2_X1 U449 ( .A(n381), .B(n380), .ZN(n383) );
  XOR2_X1 U450 ( .A(G162GAT), .B(G85GAT), .Z(n382) );
  XNOR2_X1 U451 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U452 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U453 ( .A(n387), .B(n386), .Z(n517) );
  INV_X1 U454 ( .A(n517), .ZN(n548) );
  INV_X1 U455 ( .A(n504), .ZN(n524) );
  NOR2_X1 U456 ( .A1(n548), .A2(n524), .ZN(n388) );
  NAND2_X1 U457 ( .A1(n389), .A2(n388), .ZN(n529) );
  OR2_X1 U458 ( .A1(n546), .A2(n392), .ZN(n390) );
  NOR2_X1 U459 ( .A1(n391), .A2(n390), .ZN(n395) );
  INV_X1 U460 ( .A(n392), .ZN(n393) );
  AND2_X1 U461 ( .A1(n393), .A2(n517), .ZN(n394) );
  OR2_X2 U462 ( .A1(n395), .A2(n394), .ZN(n482) );
  NOR2_X1 U463 ( .A1(n584), .A2(n482), .ZN(n396) );
  XNOR2_X1 U464 ( .A(n396), .B(KEYINPUT100), .ZN(n414) );
  XOR2_X1 U465 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n398) );
  XNOR2_X1 U466 ( .A(G106GAT), .B(G92GAT), .ZN(n397) );
  XOR2_X1 U467 ( .A(n398), .B(n397), .Z(n403) );
  XOR2_X1 U468 ( .A(G99GAT), .B(G85GAT), .Z(n439) );
  XOR2_X1 U469 ( .A(n439), .B(n399), .Z(n401) );
  XNOR2_X1 U470 ( .A(G134GAT), .B(G218GAT), .ZN(n400) );
  XNOR2_X1 U471 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U472 ( .A(n403), .B(n402), .ZN(n405) );
  NAND2_X1 U473 ( .A1(G232GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U474 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U475 ( .A(n406), .B(KEYINPUT11), .Z(n409) );
  XNOR2_X1 U476 ( .A(n407), .B(KEYINPUT74), .ZN(n408) );
  XNOR2_X1 U477 ( .A(n409), .B(n408), .ZN(n413) );
  XOR2_X1 U478 ( .A(KEYINPUT8), .B(KEYINPUT67), .Z(n411) );
  XNOR2_X1 U479 ( .A(G43GAT), .B(G29GAT), .ZN(n410) );
  XNOR2_X1 U480 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U481 ( .A(KEYINPUT7), .B(n412), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n413), .B(n421), .ZN(n479) );
  XOR2_X1 U483 ( .A(KEYINPUT36), .B(n479), .Z(n586) );
  NAND2_X1 U484 ( .A1(n414), .A2(n586), .ZN(n415) );
  XOR2_X1 U485 ( .A(KEYINPUT37), .B(n415), .Z(n516) );
  XOR2_X1 U486 ( .A(G197GAT), .B(G113GAT), .Z(n417) );
  XNOR2_X1 U487 ( .A(G36GAT), .B(G50GAT), .ZN(n416) );
  XNOR2_X1 U488 ( .A(n417), .B(n416), .ZN(n419) );
  XOR2_X1 U489 ( .A(n419), .B(n418), .Z(n423) );
  XOR2_X1 U490 ( .A(n421), .B(n420), .Z(n422) );
  XNOR2_X1 U491 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U492 ( .A(KEYINPUT66), .B(KEYINPUT65), .Z(n425) );
  NAND2_X1 U493 ( .A1(G229GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U494 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U495 ( .A(n427), .B(n426), .Z(n433) );
  XOR2_X1 U496 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n429) );
  XNOR2_X1 U497 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n428) );
  XNOR2_X1 U498 ( .A(n429), .B(n428), .ZN(n431) );
  XNOR2_X1 U499 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U500 ( .A(n433), .B(n432), .Z(n506) );
  INV_X1 U501 ( .A(n506), .ZN(n575) );
  NAND2_X1 U502 ( .A1(G230GAT), .A2(G233GAT), .ZN(n435) );
  XOR2_X1 U503 ( .A(n438), .B(KEYINPUT73), .Z(n444) );
  XNOR2_X1 U504 ( .A(G120GAT), .B(n439), .ZN(n442) );
  XOR2_X1 U505 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n441) );
  XNOR2_X1 U506 ( .A(KEYINPUT31), .B(KEYINPUT70), .ZN(n440) );
  XNOR2_X1 U507 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U508 ( .A(n448), .B(n447), .ZN(n578) );
  NAND2_X1 U509 ( .A1(n575), .A2(n578), .ZN(n485) );
  XOR2_X1 U510 ( .A(KEYINPUT38), .B(n449), .Z(n503) );
  NOR2_X1 U511 ( .A1(n503), .A2(n530), .ZN(n453) );
  XNOR2_X1 U512 ( .A(KEYINPUT102), .B(KEYINPUT40), .ZN(n451) );
  INV_X1 U513 ( .A(G43GAT), .ZN(n450) );
  XNOR2_X1 U514 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n467) );
  XNOR2_X1 U515 ( .A(KEYINPUT45), .B(KEYINPUT107), .ZN(n455) );
  AND2_X1 U516 ( .A1(n586), .A2(n584), .ZN(n454) );
  XNOR2_X1 U517 ( .A(n455), .B(n454), .ZN(n456) );
  NOR2_X1 U518 ( .A1(n575), .A2(n456), .ZN(n457) );
  NAND2_X1 U519 ( .A1(n578), .A2(n457), .ZN(n458) );
  XNOR2_X1 U520 ( .A(KEYINPUT108), .B(n458), .ZN(n465) );
  XOR2_X1 U521 ( .A(KEYINPUT106), .B(KEYINPUT47), .Z(n463) );
  XNOR2_X1 U522 ( .A(n578), .B(KEYINPUT41), .ZN(n550) );
  NAND2_X1 U523 ( .A1(n575), .A2(n550), .ZN(n459) );
  XNOR2_X1 U524 ( .A(KEYINPUT46), .B(n459), .ZN(n460) );
  NAND2_X1 U525 ( .A1(n460), .A2(n479), .ZN(n461) );
  OR2_X1 U526 ( .A1(n584), .A2(n461), .ZN(n462) );
  XNOR2_X1 U527 ( .A(n463), .B(n462), .ZN(n464) );
  NAND2_X1 U528 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U529 ( .A1(n545), .A2(n519), .ZN(n470) );
  XNOR2_X1 U530 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n468) );
  XNOR2_X1 U531 ( .A(n468), .B(KEYINPUT54), .ZN(n469) );
  XNOR2_X1 U532 ( .A(n470), .B(n469), .ZN(n471) );
  NAND2_X1 U533 ( .A1(n471), .A2(n548), .ZN(n573) );
  NOR2_X1 U534 ( .A1(n472), .A2(n573), .ZN(n473) );
  XNOR2_X1 U535 ( .A(n473), .B(KEYINPUT55), .ZN(n474) );
  INV_X1 U536 ( .A(n479), .ZN(n556) );
  NAND2_X1 U537 ( .A1(n569), .A2(n556), .ZN(n478) );
  XOR2_X1 U538 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n476) );
  XNOR2_X1 U539 ( .A(G190GAT), .B(KEYINPUT122), .ZN(n475) );
  XOR2_X1 U540 ( .A(KEYINPUT16), .B(KEYINPUT80), .Z(n481) );
  NAND2_X1 U541 ( .A1(n584), .A2(n479), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n481), .B(n480), .ZN(n484) );
  INV_X1 U543 ( .A(n482), .ZN(n483) );
  NAND2_X1 U544 ( .A1(n484), .A2(n483), .ZN(n507) );
  NOR2_X1 U545 ( .A1(n485), .A2(n507), .ZN(n486) );
  XNOR2_X1 U546 ( .A(KEYINPUT95), .B(n486), .ZN(n495) );
  NOR2_X1 U547 ( .A1(n548), .A2(n495), .ZN(n488) );
  XNOR2_X1 U548 ( .A(KEYINPUT96), .B(KEYINPUT34), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(n489) );
  XOR2_X1 U550 ( .A(G1GAT), .B(n489), .Z(G1324GAT) );
  NOR2_X1 U551 ( .A1(n500), .A2(n495), .ZN(n491) );
  XNOR2_X1 U552 ( .A(G8GAT), .B(KEYINPUT97), .ZN(n490) );
  XNOR2_X1 U553 ( .A(n491), .B(n490), .ZN(G1325GAT) );
  NOR2_X1 U554 ( .A1(n530), .A2(n495), .ZN(n493) );
  XNOR2_X1 U555 ( .A(KEYINPUT98), .B(KEYINPUT35), .ZN(n492) );
  XNOR2_X1 U556 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U557 ( .A(G15GAT), .B(n494), .ZN(G1326GAT) );
  NOR2_X1 U558 ( .A1(n504), .A2(n495), .ZN(n497) );
  XNOR2_X1 U559 ( .A(G22GAT), .B(KEYINPUT99), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n497), .B(n496), .ZN(G1327GAT) );
  NOR2_X1 U561 ( .A1(n503), .A2(n548), .ZN(n499) );
  XNOR2_X1 U562 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n499), .B(n498), .ZN(G1328GAT) );
  XNOR2_X1 U564 ( .A(G36GAT), .B(KEYINPUT101), .ZN(n502) );
  NOR2_X1 U565 ( .A1(n500), .A2(n503), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n502), .B(n501), .ZN(G1329GAT) );
  NOR2_X1 U567 ( .A1(n504), .A2(n503), .ZN(n505) );
  XOR2_X1 U568 ( .A(G50GAT), .B(n505), .Z(G1331GAT) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n509) );
  XOR2_X1 U570 ( .A(KEYINPUT103), .B(n550), .Z(n566) );
  NAND2_X1 U571 ( .A1(n506), .A2(n566), .ZN(n515) );
  NAND2_X1 U572 ( .A1(n517), .A2(n512), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(G1332GAT) );
  NAND2_X1 U574 ( .A1(n519), .A2(n512), .ZN(n510) );
  XNOR2_X1 U575 ( .A(n510), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U576 ( .A1(n512), .A2(n522), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n511), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U579 ( .A1(n512), .A2(n524), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  NOR2_X1 U581 ( .A1(n516), .A2(n515), .ZN(n525) );
  NAND2_X1 U582 ( .A1(n517), .A2(n525), .ZN(n518) );
  XNOR2_X1 U583 ( .A(G85GAT), .B(n518), .ZN(G1336GAT) );
  NAND2_X1 U584 ( .A1(n519), .A2(n525), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n520), .B(KEYINPUT104), .ZN(n521) );
  XNOR2_X1 U586 ( .A(G92GAT), .B(n521), .ZN(G1337GAT) );
  NAND2_X1 U587 ( .A1(n525), .A2(n522), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n523), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT44), .B(KEYINPUT105), .Z(n527) );
  NAND2_X1 U590 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U591 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  NOR2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n531) );
  NAND2_X1 U594 ( .A1(n545), .A2(n531), .ZN(n532) );
  XNOR2_X1 U595 ( .A(n532), .B(KEYINPUT109), .ZN(n541) );
  NAND2_X1 U596 ( .A1(n541), .A2(n575), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n533), .B(KEYINPUT110), .ZN(n534) );
  XNOR2_X1 U598 ( .A(G113GAT), .B(n534), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT111), .B(KEYINPUT49), .Z(n536) );
  NAND2_X1 U600 ( .A1(n541), .A2(n566), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U602 ( .A(G120GAT), .B(n537), .Z(G1341GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT112), .B(KEYINPUT50), .Z(n539) );
  NAND2_X1 U604 ( .A1(n541), .A2(n584), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U606 ( .A(G127GAT), .B(n540), .Z(G1342GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U608 ( .A1(n541), .A2(n556), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U610 ( .A(G134GAT), .B(n544), .Z(G1343GAT) );
  NAND2_X1 U611 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U612 ( .A1(n548), .A2(n547), .ZN(n557) );
  NAND2_X1 U613 ( .A1(n557), .A2(n575), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n549), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n552) );
  NAND2_X1 U616 ( .A1(n557), .A2(n550), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(n553), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n557), .A2(n584), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n554), .B(KEYINPUT114), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(n555), .ZN(G1346GAT) );
  XOR2_X1 U622 ( .A(G162GAT), .B(KEYINPUT115), .Z(n559) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(G1347GAT) );
  NAND2_X1 U625 ( .A1(n569), .A2(n575), .ZN(n562) );
  XOR2_X1 U626 ( .A(G169GAT), .B(KEYINPUT118), .Z(n560) );
  XNOR2_X1 U627 ( .A(KEYINPUT119), .B(n560), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1348GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT57), .B(KEYINPUT121), .Z(n564) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U632 ( .A(KEYINPUT56), .B(n565), .Z(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n566), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1349GAT) );
  NAND2_X1 U635 ( .A1(n569), .A2(n584), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(KEYINPUT60), .ZN(n572) );
  XOR2_X1 U639 ( .A(KEYINPUT124), .B(n572), .Z(n577) );
  NOR2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n587) );
  NAND2_X1 U641 ( .A1(n587), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  INV_X1 U643 ( .A(n587), .ZN(n579) );
  NOR2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n583) );
  XOR2_X1 U645 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n581) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NAND2_X1 U649 ( .A1(n587), .A2(n584), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n585), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U651 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n589) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U654 ( .A(G218GAT), .B(n590), .ZN(G1355GAT) );
endmodule

