

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U550 ( .A1(n676), .A2(n780), .ZN(n720) );
  NOR2_X2 U551 ( .A1(n690), .A2(n689), .ZN(n695) );
  OR2_X1 U552 ( .A1(n673), .A2(n714), .ZN(n674) );
  INV_X1 U553 ( .A(KEYINPUT101), .ZN(n715) );
  XOR2_X1 U554 ( .A(n711), .B(KEYINPUT29), .Z(n516) );
  XOR2_X1 U555 ( .A(n760), .B(KEYINPUT94), .Z(n517) );
  INV_X1 U556 ( .A(KEYINPUT100), .ZN(n696) );
  INV_X1 U557 ( .A(G8), .ZN(n672) );
  OR2_X1 U558 ( .A1(n717), .A2(n672), .ZN(n673) );
  AND2_X1 U559 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U560 ( .A1(n731), .A2(G8), .ZN(n732) );
  NAND2_X1 U561 ( .A1(G8), .A2(n720), .ZN(n759) );
  AND2_X1 U562 ( .A1(n761), .A2(n517), .ZN(n762) );
  NOR2_X1 U563 ( .A1(G651), .A2(n629), .ZN(n638) );
  NOR2_X2 U564 ( .A1(n580), .A2(n579), .ZN(n962) );
  XOR2_X1 U565 ( .A(KEYINPUT66), .B(KEYINPUT23), .Z(n519) );
  INV_X1 U566 ( .A(G2105), .ZN(n524) );
  AND2_X4 U567 ( .A1(n524), .A2(G2104), .ZN(n862) );
  NAND2_X1 U568 ( .A1(G101), .A2(n862), .ZN(n518) );
  XNOR2_X1 U569 ( .A(n519), .B(n518), .ZN(n521) );
  AND2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n864) );
  NAND2_X1 U571 ( .A1(n864), .A2(G113), .ZN(n520) );
  NAND2_X1 U572 ( .A1(n521), .A2(n520), .ZN(n528) );
  XNOR2_X1 U573 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n523) );
  NOR2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  XNOR2_X2 U575 ( .A(n523), .B(n522), .ZN(n861) );
  NAND2_X1 U576 ( .A1(G137), .A2(n861), .ZN(n526) );
  NOR2_X2 U577 ( .A1(G2104), .A2(n524), .ZN(n865) );
  NAND2_X1 U578 ( .A1(G125), .A2(n865), .ZN(n525) );
  NAND2_X1 U579 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U580 ( .A1(n528), .A2(n527), .ZN(G160) );
  NAND2_X1 U581 ( .A1(G102), .A2(n862), .ZN(n530) );
  NAND2_X1 U582 ( .A1(G138), .A2(n861), .ZN(n529) );
  NAND2_X1 U583 ( .A1(n530), .A2(n529), .ZN(n534) );
  NAND2_X1 U584 ( .A1(G114), .A2(n864), .ZN(n532) );
  NAND2_X1 U585 ( .A1(G126), .A2(n865), .ZN(n531) );
  NAND2_X1 U586 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U587 ( .A1(n534), .A2(n533), .ZN(G164) );
  XOR2_X1 U588 ( .A(G543), .B(KEYINPUT0), .Z(n629) );
  NAND2_X1 U589 ( .A1(G52), .A2(n638), .ZN(n537) );
  INV_X1 U590 ( .A(G651), .ZN(n538) );
  NOR2_X1 U591 ( .A1(G543), .A2(n538), .ZN(n535) );
  XOR2_X2 U592 ( .A(KEYINPUT1), .B(n535), .Z(n633) );
  NAND2_X1 U593 ( .A1(G64), .A2(n633), .ZN(n536) );
  NAND2_X1 U594 ( .A1(n537), .A2(n536), .ZN(n543) );
  NOR2_X2 U595 ( .A1(n629), .A2(n538), .ZN(n634) );
  NAND2_X1 U596 ( .A1(G77), .A2(n634), .ZN(n540) );
  NOR2_X1 U597 ( .A1(G543), .A2(G651), .ZN(n635) );
  NAND2_X1 U598 ( .A1(G90), .A2(n635), .ZN(n539) );
  NAND2_X1 U599 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U600 ( .A(KEYINPUT9), .B(n541), .Z(n542) );
  NOR2_X1 U601 ( .A1(n543), .A2(n542), .ZN(G171) );
  AND2_X1 U602 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U603 ( .A1(G111), .A2(n864), .ZN(n545) );
  NAND2_X1 U604 ( .A1(G135), .A2(n861), .ZN(n544) );
  NAND2_X1 U605 ( .A1(n545), .A2(n544), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n865), .A2(G123), .ZN(n546) );
  XOR2_X1 U607 ( .A(KEYINPUT18), .B(n546), .Z(n547) );
  NOR2_X1 U608 ( .A1(n548), .A2(n547), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n862), .A2(G99), .ZN(n549) );
  NAND2_X1 U610 ( .A1(n550), .A2(n549), .ZN(n915) );
  XNOR2_X1 U611 ( .A(G2096), .B(n915), .ZN(n551) );
  OR2_X1 U612 ( .A1(G2100), .A2(n551), .ZN(G156) );
  INV_X1 U613 ( .A(G57), .ZN(G237) );
  INV_X1 U614 ( .A(G69), .ZN(G235) );
  INV_X1 U615 ( .A(G108), .ZN(G238) );
  INV_X1 U616 ( .A(G120), .ZN(G236) );
  INV_X1 U617 ( .A(G132), .ZN(G219) );
  INV_X1 U618 ( .A(G82), .ZN(G220) );
  NAND2_X1 U619 ( .A1(G88), .A2(n635), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n552), .B(KEYINPUT82), .ZN(n554) );
  NAND2_X1 U621 ( .A1(n634), .A2(G75), .ZN(n553) );
  NAND2_X1 U622 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U623 ( .A1(G50), .A2(n638), .ZN(n556) );
  NAND2_X1 U624 ( .A1(G62), .A2(n633), .ZN(n555) );
  NAND2_X1 U625 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U626 ( .A1(n558), .A2(n557), .ZN(G166) );
  NAND2_X1 U627 ( .A1(n635), .A2(G89), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n559), .B(KEYINPUT4), .ZN(n561) );
  NAND2_X1 U629 ( .A1(G76), .A2(n634), .ZN(n560) );
  NAND2_X1 U630 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n562), .B(KEYINPUT5), .ZN(n567) );
  NAND2_X1 U632 ( .A1(G51), .A2(n638), .ZN(n564) );
  NAND2_X1 U633 ( .A1(G63), .A2(n633), .ZN(n563) );
  NAND2_X1 U634 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U635 ( .A(KEYINPUT6), .B(n565), .Z(n566) );
  NAND2_X1 U636 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U637 ( .A(n568), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U638 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U639 ( .A1(G7), .A2(G661), .ZN(n569) );
  XNOR2_X1 U640 ( .A(n569), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U641 ( .A(G223), .ZN(n818) );
  AND2_X1 U642 ( .A1(n818), .A2(G567), .ZN(n571) );
  XNOR2_X1 U643 ( .A(KEYINPUT11), .B(KEYINPUT72), .ZN(n570) );
  XNOR2_X1 U644 ( .A(n571), .B(n570), .ZN(G234) );
  NAND2_X1 U645 ( .A1(G68), .A2(n634), .ZN(n574) );
  NAND2_X1 U646 ( .A1(n635), .A2(G81), .ZN(n572) );
  XNOR2_X1 U647 ( .A(n572), .B(KEYINPUT12), .ZN(n573) );
  NAND2_X1 U648 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U649 ( .A(n575), .B(KEYINPUT13), .ZN(n577) );
  NAND2_X1 U650 ( .A1(G43), .A2(n638), .ZN(n576) );
  NAND2_X1 U651 ( .A1(n577), .A2(n576), .ZN(n580) );
  NAND2_X1 U652 ( .A1(n633), .A2(G56), .ZN(n578) );
  XOR2_X1 U653 ( .A(KEYINPUT14), .B(n578), .Z(n579) );
  NAND2_X1 U654 ( .A1(n962), .A2(G860), .ZN(G153) );
  INV_X1 U655 ( .A(G171), .ZN(G301) );
  NAND2_X1 U656 ( .A1(G868), .A2(G301), .ZN(n589) );
  NAND2_X1 U657 ( .A1(G79), .A2(n634), .ZN(n582) );
  NAND2_X1 U658 ( .A1(G92), .A2(n635), .ZN(n581) );
  NAND2_X1 U659 ( .A1(n582), .A2(n581), .ZN(n586) );
  NAND2_X1 U660 ( .A1(G54), .A2(n638), .ZN(n584) );
  NAND2_X1 U661 ( .A1(G66), .A2(n633), .ZN(n583) );
  NAND2_X1 U662 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U663 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U664 ( .A(KEYINPUT15), .B(n587), .Z(n967) );
  OR2_X1 U665 ( .A1(n967), .A2(G868), .ZN(n588) );
  NAND2_X1 U666 ( .A1(n589), .A2(n588), .ZN(G284) );
  NAND2_X1 U667 ( .A1(G78), .A2(n634), .ZN(n591) );
  NAND2_X1 U668 ( .A1(G91), .A2(n635), .ZN(n590) );
  NAND2_X1 U669 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U670 ( .A1(G65), .A2(n633), .ZN(n592) );
  XNOR2_X1 U671 ( .A(KEYINPUT71), .B(n592), .ZN(n593) );
  NOR2_X1 U672 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U673 ( .A1(n638), .A2(G53), .ZN(n595) );
  NAND2_X1 U674 ( .A1(n596), .A2(n595), .ZN(G299) );
  XNOR2_X1 U675 ( .A(KEYINPUT73), .B(G868), .ZN(n597) );
  NOR2_X1 U676 ( .A1(G286), .A2(n597), .ZN(n600) );
  NOR2_X1 U677 ( .A1(G868), .A2(G299), .ZN(n598) );
  XNOR2_X1 U678 ( .A(n598), .B(KEYINPUT74), .ZN(n599) );
  NOR2_X1 U679 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U680 ( .A(KEYINPUT75), .B(n601), .Z(G297) );
  INV_X1 U681 ( .A(G860), .ZN(n602) );
  NAND2_X1 U682 ( .A1(n602), .A2(G559), .ZN(n603) );
  NAND2_X1 U683 ( .A1(n603), .A2(n967), .ZN(n604) );
  XNOR2_X1 U684 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  INV_X1 U685 ( .A(G868), .ZN(n653) );
  NAND2_X1 U686 ( .A1(n962), .A2(n653), .ZN(n605) );
  XOR2_X1 U687 ( .A(KEYINPUT76), .B(n605), .Z(n608) );
  NAND2_X1 U688 ( .A1(G868), .A2(n967), .ZN(n606) );
  NOR2_X1 U689 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U690 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U691 ( .A1(G72), .A2(n634), .ZN(n610) );
  NAND2_X1 U692 ( .A1(G85), .A2(n635), .ZN(n609) );
  NAND2_X1 U693 ( .A1(n610), .A2(n609), .ZN(n611) );
  XOR2_X1 U694 ( .A(KEYINPUT68), .B(n611), .Z(n617) );
  NAND2_X1 U695 ( .A1(n638), .A2(G47), .ZN(n612) );
  XOR2_X1 U696 ( .A(KEYINPUT69), .B(n612), .Z(n614) );
  NAND2_X1 U697 ( .A1(n633), .A2(G60), .ZN(n613) );
  NAND2_X1 U698 ( .A1(n614), .A2(n613), .ZN(n615) );
  XOR2_X1 U699 ( .A(KEYINPUT70), .B(n615), .Z(n616) );
  NAND2_X1 U700 ( .A1(n617), .A2(n616), .ZN(G290) );
  NAND2_X1 U701 ( .A1(n634), .A2(G73), .ZN(n618) );
  XNOR2_X1 U702 ( .A(n618), .B(KEYINPUT2), .ZN(n620) );
  NAND2_X1 U703 ( .A1(G86), .A2(n635), .ZN(n619) );
  NAND2_X1 U704 ( .A1(n620), .A2(n619), .ZN(n623) );
  NAND2_X1 U705 ( .A1(G48), .A2(n638), .ZN(n621) );
  XNOR2_X1 U706 ( .A(KEYINPUT81), .B(n621), .ZN(n622) );
  NOR2_X1 U707 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n633), .A2(G61), .ZN(n624) );
  NAND2_X1 U709 ( .A1(n625), .A2(n624), .ZN(G305) );
  NAND2_X1 U710 ( .A1(G49), .A2(n638), .ZN(n627) );
  NAND2_X1 U711 ( .A1(G74), .A2(G651), .ZN(n626) );
  NAND2_X1 U712 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U713 ( .A1(n633), .A2(n628), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n629), .A2(G87), .ZN(n630) );
  NAND2_X1 U715 ( .A1(n631), .A2(n630), .ZN(G288) );
  NAND2_X1 U716 ( .A1(G559), .A2(n967), .ZN(n632) );
  XOR2_X1 U717 ( .A(n962), .B(n632), .Z(n907) );
  NAND2_X1 U718 ( .A1(n633), .A2(G67), .ZN(n643) );
  NAND2_X1 U719 ( .A1(G80), .A2(n634), .ZN(n637) );
  NAND2_X1 U720 ( .A1(G93), .A2(n635), .ZN(n636) );
  NAND2_X1 U721 ( .A1(n637), .A2(n636), .ZN(n641) );
  NAND2_X1 U722 ( .A1(G55), .A2(n638), .ZN(n639) );
  XNOR2_X1 U723 ( .A(KEYINPUT79), .B(n639), .ZN(n640) );
  NOR2_X1 U724 ( .A1(n641), .A2(n640), .ZN(n642) );
  NAND2_X1 U725 ( .A1(n643), .A2(n642), .ZN(n644) );
  XOR2_X1 U726 ( .A(KEYINPUT80), .B(n644), .Z(n911) );
  INV_X1 U727 ( .A(G299), .ZN(n971) );
  XNOR2_X1 U728 ( .A(KEYINPUT83), .B(KEYINPUT84), .ZN(n646) );
  XNOR2_X1 U729 ( .A(G305), .B(KEYINPUT19), .ZN(n645) );
  XNOR2_X1 U730 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U731 ( .A(n971), .B(n647), .ZN(n649) );
  XNOR2_X1 U732 ( .A(G288), .B(G166), .ZN(n648) );
  XNOR2_X1 U733 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U734 ( .A(n911), .B(n650), .ZN(n651) );
  XNOR2_X1 U735 ( .A(G290), .B(n651), .ZN(n884) );
  XNOR2_X1 U736 ( .A(n907), .B(n884), .ZN(n652) );
  NAND2_X1 U737 ( .A1(n652), .A2(G868), .ZN(n655) );
  NAND2_X1 U738 ( .A1(n653), .A2(n911), .ZN(n654) );
  NAND2_X1 U739 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U740 ( .A(KEYINPUT85), .B(n656), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2084), .A2(G2078), .ZN(n657) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n657), .Z(n658) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n658), .ZN(n659) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(n659), .ZN(n660) );
  NAND2_X1 U745 ( .A1(n660), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U746 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U747 ( .A1(G220), .A2(G219), .ZN(n661) );
  XOR2_X1 U748 ( .A(KEYINPUT22), .B(n661), .Z(n662) );
  NOR2_X1 U749 ( .A1(G218), .A2(n662), .ZN(n663) );
  NAND2_X1 U750 ( .A1(G96), .A2(n663), .ZN(n905) );
  NAND2_X1 U751 ( .A1(G2106), .A2(n905), .ZN(n664) );
  XOR2_X1 U752 ( .A(KEYINPUT86), .B(n664), .Z(n669) );
  NOR2_X1 U753 ( .A1(G236), .A2(G238), .ZN(n666) );
  NOR2_X1 U754 ( .A1(G235), .A2(G237), .ZN(n665) );
  NAND2_X1 U755 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U756 ( .A(KEYINPUT87), .B(n667), .Z(n906) );
  AND2_X1 U757 ( .A1(n906), .A2(G567), .ZN(n668) );
  NOR2_X1 U758 ( .A1(n669), .A2(n668), .ZN(G319) );
  INV_X1 U759 ( .A(G319), .ZN(n671) );
  NAND2_X1 U760 ( .A1(G661), .A2(G483), .ZN(n670) );
  NOR2_X1 U761 ( .A1(n671), .A2(n670), .ZN(n822) );
  NAND2_X1 U762 ( .A1(n822), .A2(G36), .ZN(G176) );
  INV_X1 U763 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U764 ( .A(G1981), .B(G305), .ZN(n965) );
  NAND2_X1 U765 ( .A1(G160), .A2(G40), .ZN(n781) );
  INV_X1 U766 ( .A(n781), .ZN(n676) );
  NOR2_X1 U767 ( .A1(G164), .A2(G1384), .ZN(n780) );
  NOR2_X1 U768 ( .A1(G1966), .A2(n759), .ZN(n714) );
  NOR2_X1 U769 ( .A1(G2084), .A2(n720), .ZN(n717) );
  XNOR2_X1 U770 ( .A(KEYINPUT30), .B(n674), .ZN(n675) );
  NOR2_X1 U771 ( .A1(G168), .A2(n675), .ZN(n681) );
  INV_X1 U772 ( .A(G1961), .ZN(n991) );
  NAND2_X1 U773 ( .A1(n720), .A2(n991), .ZN(n679) );
  AND2_X2 U774 ( .A1(n676), .A2(n780), .ZN(n701) );
  XOR2_X1 U775 ( .A(G2078), .B(KEYINPUT95), .Z(n677) );
  XNOR2_X1 U776 ( .A(KEYINPUT25), .B(n677), .ZN(n948) );
  NAND2_X1 U777 ( .A1(n701), .A2(n948), .ZN(n678) );
  NAND2_X1 U778 ( .A1(n679), .A2(n678), .ZN(n683) );
  NOR2_X1 U779 ( .A1(G171), .A2(n683), .ZN(n680) );
  NOR2_X1 U780 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U781 ( .A(KEYINPUT31), .B(n682), .Z(n724) );
  NAND2_X1 U782 ( .A1(n683), .A2(G171), .ZN(n712) );
  NAND2_X1 U783 ( .A1(G1996), .A2(n701), .ZN(n686) );
  XOR2_X1 U784 ( .A(KEYINPUT26), .B(KEYINPUT98), .Z(n684) );
  XNOR2_X1 U785 ( .A(KEYINPUT65), .B(n684), .ZN(n685) );
  XNOR2_X1 U786 ( .A(n686), .B(n685), .ZN(n687) );
  NAND2_X1 U787 ( .A1(n687), .A2(n962), .ZN(n690) );
  NAND2_X1 U788 ( .A1(G1341), .A2(n720), .ZN(n688) );
  XNOR2_X1 U789 ( .A(n688), .B(KEYINPUT99), .ZN(n689) );
  NAND2_X1 U790 ( .A1(n695), .A2(n967), .ZN(n694) );
  NOR2_X1 U791 ( .A1(G2067), .A2(n720), .ZN(n692) );
  NOR2_X1 U792 ( .A1(n701), .A2(G1348), .ZN(n691) );
  NOR2_X1 U793 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U794 ( .A1(n694), .A2(n693), .ZN(n699) );
  NOR2_X1 U795 ( .A1(n695), .A2(n967), .ZN(n697) );
  XNOR2_X1 U796 ( .A(n697), .B(n696), .ZN(n698) );
  NAND2_X1 U797 ( .A1(n699), .A2(n698), .ZN(n705) );
  NAND2_X1 U798 ( .A1(n701), .A2(G2072), .ZN(n700) );
  XNOR2_X1 U799 ( .A(n700), .B(KEYINPUT27), .ZN(n703) );
  XOR2_X1 U800 ( .A(G1956), .B(KEYINPUT96), .Z(n997) );
  NOR2_X1 U801 ( .A1(n701), .A2(n997), .ZN(n702) );
  NOR2_X1 U802 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U803 ( .A1(n971), .A2(n706), .ZN(n704) );
  NAND2_X1 U804 ( .A1(n705), .A2(n704), .ZN(n710) );
  NOR2_X1 U805 ( .A1(n971), .A2(n706), .ZN(n708) );
  XNOR2_X1 U806 ( .A(KEYINPUT97), .B(KEYINPUT28), .ZN(n707) );
  XNOR2_X1 U807 ( .A(n708), .B(n707), .ZN(n709) );
  NAND2_X1 U808 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U809 ( .A1(n712), .A2(n516), .ZN(n726) );
  AND2_X1 U810 ( .A1(n724), .A2(n726), .ZN(n713) );
  NOR2_X1 U811 ( .A1(n714), .A2(n713), .ZN(n716) );
  XNOR2_X1 U812 ( .A(n716), .B(n715), .ZN(n719) );
  NAND2_X1 U813 ( .A1(G8), .A2(n717), .ZN(n718) );
  NAND2_X1 U814 ( .A1(n719), .A2(n718), .ZN(n753) );
  NOR2_X1 U815 ( .A1(G1971), .A2(n759), .ZN(n722) );
  NOR2_X1 U816 ( .A1(G2090), .A2(n720), .ZN(n721) );
  NOR2_X1 U817 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U818 ( .A1(n723), .A2(G303), .ZN(n727) );
  AND2_X1 U819 ( .A1(n724), .A2(n727), .ZN(n725) );
  NAND2_X1 U820 ( .A1(n726), .A2(n725), .ZN(n730) );
  INV_X1 U821 ( .A(n727), .ZN(n728) );
  OR2_X1 U822 ( .A1(n728), .A2(G286), .ZN(n729) );
  XNOR2_X1 U823 ( .A(n732), .B(KEYINPUT32), .ZN(n752) );
  INV_X1 U824 ( .A(n759), .ZN(n733) );
  NAND2_X1 U825 ( .A1(G1976), .A2(G288), .ZN(n969) );
  AND2_X1 U826 ( .A1(n733), .A2(n969), .ZN(n735) );
  AND2_X1 U827 ( .A1(n752), .A2(n735), .ZN(n734) );
  NAND2_X1 U828 ( .A1(n753), .A2(n734), .ZN(n740) );
  INV_X1 U829 ( .A(n735), .ZN(n738) );
  NOR2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n972) );
  NOR2_X1 U831 ( .A1(G1971), .A2(G303), .ZN(n736) );
  NOR2_X1 U832 ( .A1(n972), .A2(n736), .ZN(n737) );
  OR2_X1 U833 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U834 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U835 ( .A(n741), .B(KEYINPUT64), .ZN(n742) );
  NOR2_X1 U836 ( .A1(KEYINPUT33), .A2(n742), .ZN(n746) );
  NAND2_X1 U837 ( .A1(KEYINPUT33), .A2(n972), .ZN(n743) );
  NOR2_X1 U838 ( .A1(n759), .A2(n743), .ZN(n744) );
  XNOR2_X1 U839 ( .A(n744), .B(KEYINPUT102), .ZN(n745) );
  NOR2_X1 U840 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U841 ( .A(n747), .B(KEYINPUT103), .ZN(n748) );
  NOR2_X1 U842 ( .A1(n965), .A2(n748), .ZN(n749) );
  INV_X1 U843 ( .A(n749), .ZN(n763) );
  NOR2_X1 U844 ( .A1(G2090), .A2(G303), .ZN(n750) );
  NAND2_X1 U845 ( .A1(G8), .A2(n750), .ZN(n751) );
  XNOR2_X1 U846 ( .A(n751), .B(KEYINPUT104), .ZN(n755) );
  NAND2_X1 U847 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U848 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U849 ( .A1(n756), .A2(n759), .ZN(n761) );
  NOR2_X1 U850 ( .A1(G1981), .A2(G305), .ZN(n757) );
  XOR2_X1 U851 ( .A(n757), .B(KEYINPUT24), .Z(n758) );
  NOR2_X1 U852 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U853 ( .A1(n763), .A2(n762), .ZN(n785) );
  NAND2_X1 U854 ( .A1(G107), .A2(n864), .ZN(n765) );
  NAND2_X1 U855 ( .A1(G119), .A2(n865), .ZN(n764) );
  NAND2_X1 U856 ( .A1(n765), .A2(n764), .ZN(n768) );
  NAND2_X1 U857 ( .A1(G131), .A2(n861), .ZN(n766) );
  XNOR2_X1 U858 ( .A(KEYINPUT91), .B(n766), .ZN(n767) );
  NOR2_X1 U859 ( .A1(n768), .A2(n767), .ZN(n770) );
  NAND2_X1 U860 ( .A1(n862), .A2(G95), .ZN(n769) );
  NAND2_X1 U861 ( .A1(n770), .A2(n769), .ZN(n848) );
  XNOR2_X1 U862 ( .A(KEYINPUT92), .B(G1991), .ZN(n943) );
  NAND2_X1 U863 ( .A1(n848), .A2(n943), .ZN(n779) );
  NAND2_X1 U864 ( .A1(G117), .A2(n864), .ZN(n772) );
  NAND2_X1 U865 ( .A1(G141), .A2(n861), .ZN(n771) );
  NAND2_X1 U866 ( .A1(n772), .A2(n771), .ZN(n775) );
  NAND2_X1 U867 ( .A1(n862), .A2(G105), .ZN(n773) );
  XOR2_X1 U868 ( .A(KEYINPUT38), .B(n773), .Z(n774) );
  NOR2_X1 U869 ( .A1(n775), .A2(n774), .ZN(n777) );
  NAND2_X1 U870 ( .A1(n865), .A2(G129), .ZN(n776) );
  NAND2_X1 U871 ( .A1(n777), .A2(n776), .ZN(n878) );
  NAND2_X1 U872 ( .A1(G1996), .A2(n878), .ZN(n778) );
  NAND2_X1 U873 ( .A1(n779), .A2(n778), .ZN(n931) );
  NOR2_X1 U874 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U875 ( .A(n782), .B(KEYINPUT88), .ZN(n812) );
  NAND2_X1 U876 ( .A1(n931), .A2(n812), .ZN(n783) );
  XNOR2_X1 U877 ( .A(n783), .B(KEYINPUT93), .ZN(n804) );
  INV_X1 U878 ( .A(n804), .ZN(n784) );
  NAND2_X1 U879 ( .A1(n785), .A2(n784), .ZN(n788) );
  INV_X1 U880 ( .A(n812), .ZN(n786) );
  XOR2_X1 U881 ( .A(G1986), .B(G290), .Z(n980) );
  NOR2_X1 U882 ( .A1(n786), .A2(n980), .ZN(n787) );
  NOR2_X1 U883 ( .A1(n788), .A2(n787), .ZN(n800) );
  NAND2_X1 U884 ( .A1(G104), .A2(n862), .ZN(n790) );
  NAND2_X1 U885 ( .A1(G140), .A2(n861), .ZN(n789) );
  NAND2_X1 U886 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U887 ( .A(KEYINPUT34), .B(n791), .ZN(n797) );
  NAND2_X1 U888 ( .A1(G116), .A2(n864), .ZN(n793) );
  NAND2_X1 U889 ( .A1(G128), .A2(n865), .ZN(n792) );
  NAND2_X1 U890 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U891 ( .A(KEYINPUT90), .B(n794), .Z(n795) );
  XNOR2_X1 U892 ( .A(KEYINPUT35), .B(n795), .ZN(n796) );
  NOR2_X1 U893 ( .A1(n797), .A2(n796), .ZN(n798) );
  XOR2_X1 U894 ( .A(KEYINPUT36), .B(n798), .Z(n875) );
  XNOR2_X1 U895 ( .A(G2067), .B(KEYINPUT37), .ZN(n799) );
  XNOR2_X1 U896 ( .A(n799), .B(KEYINPUT89), .ZN(n801) );
  AND2_X1 U897 ( .A1(n875), .A2(n801), .ZN(n914) );
  NAND2_X1 U898 ( .A1(n812), .A2(n914), .ZN(n807) );
  NAND2_X1 U899 ( .A1(n800), .A2(n807), .ZN(n816) );
  NOR2_X1 U900 ( .A1(n875), .A2(n801), .ZN(n913) );
  NOR2_X1 U901 ( .A1(G1996), .A2(n878), .ZN(n928) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n802) );
  NOR2_X1 U903 ( .A1(n943), .A2(n848), .ZN(n917) );
  NOR2_X1 U904 ( .A1(n802), .A2(n917), .ZN(n803) );
  NOR2_X1 U905 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U906 ( .A1(n928), .A2(n805), .ZN(n806) );
  XOR2_X1 U907 ( .A(KEYINPUT39), .B(n806), .Z(n809) );
  INV_X1 U908 ( .A(n807), .ZN(n808) );
  NOR2_X1 U909 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U910 ( .A1(n913), .A2(n810), .ZN(n811) );
  XNOR2_X1 U911 ( .A(n811), .B(KEYINPUT105), .ZN(n813) );
  NAND2_X1 U912 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U913 ( .A(n814), .B(KEYINPUT106), .ZN(n815) );
  NAND2_X1 U914 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U915 ( .A(KEYINPUT40), .B(n817), .ZN(G329) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n818), .ZN(G217) );
  NAND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n819) );
  XNOR2_X1 U918 ( .A(KEYINPUT109), .B(n819), .ZN(n820) );
  NAND2_X1 U919 ( .A1(n820), .A2(G661), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n821) );
  NAND2_X1 U921 ( .A1(n822), .A2(n821), .ZN(G188) );
  XOR2_X1 U922 ( .A(G2100), .B(G2096), .Z(n824) );
  XNOR2_X1 U923 ( .A(KEYINPUT42), .B(G2678), .ZN(n823) );
  XNOR2_X1 U924 ( .A(n824), .B(n823), .ZN(n828) );
  XOR2_X1 U925 ( .A(KEYINPUT43), .B(G2090), .Z(n826) );
  XNOR2_X1 U926 ( .A(G2072), .B(G2067), .ZN(n825) );
  XNOR2_X1 U927 ( .A(n826), .B(n825), .ZN(n827) );
  XOR2_X1 U928 ( .A(n828), .B(n827), .Z(n830) );
  XNOR2_X1 U929 ( .A(G2084), .B(G2078), .ZN(n829) );
  XNOR2_X1 U930 ( .A(n830), .B(n829), .ZN(G227) );
  XOR2_X1 U931 ( .A(G1956), .B(G1966), .Z(n832) );
  XNOR2_X1 U932 ( .A(G1976), .B(G1971), .ZN(n831) );
  XNOR2_X1 U933 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U934 ( .A(n833), .B(G2474), .Z(n835) );
  XNOR2_X1 U935 ( .A(G1961), .B(G1986), .ZN(n834) );
  XNOR2_X1 U936 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U937 ( .A(KEYINPUT41), .B(G1991), .Z(n837) );
  XNOR2_X1 U938 ( .A(G1981), .B(G1996), .ZN(n836) );
  XNOR2_X1 U939 ( .A(n837), .B(n836), .ZN(n838) );
  XNOR2_X1 U940 ( .A(n839), .B(n838), .ZN(G229) );
  NAND2_X1 U941 ( .A1(G124), .A2(n865), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n840), .B(KEYINPUT44), .ZN(n842) );
  NAND2_X1 U943 ( .A1(n864), .A2(G112), .ZN(n841) );
  NAND2_X1 U944 ( .A1(n842), .A2(n841), .ZN(n846) );
  NAND2_X1 U945 ( .A1(G100), .A2(n862), .ZN(n844) );
  NAND2_X1 U946 ( .A1(G136), .A2(n861), .ZN(n843) );
  NAND2_X1 U947 ( .A1(n844), .A2(n843), .ZN(n845) );
  NOR2_X1 U948 ( .A1(n846), .A2(n845), .ZN(G162) );
  XOR2_X1 U949 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n847) );
  XNOR2_X1 U950 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U951 ( .A(n849), .B(KEYINPUT110), .Z(n851) );
  XNOR2_X1 U952 ( .A(G164), .B(KEYINPUT46), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n860) );
  NAND2_X1 U954 ( .A1(G118), .A2(n864), .ZN(n853) );
  NAND2_X1 U955 ( .A1(G130), .A2(n865), .ZN(n852) );
  NAND2_X1 U956 ( .A1(n853), .A2(n852), .ZN(n858) );
  NAND2_X1 U957 ( .A1(G106), .A2(n862), .ZN(n855) );
  NAND2_X1 U958 ( .A1(G142), .A2(n861), .ZN(n854) );
  NAND2_X1 U959 ( .A1(n855), .A2(n854), .ZN(n856) );
  XOR2_X1 U960 ( .A(KEYINPUT45), .B(n856), .Z(n857) );
  NOR2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n859) );
  XOR2_X1 U962 ( .A(n860), .B(n859), .Z(n877) );
  NAND2_X1 U963 ( .A1(G139), .A2(n861), .ZN(n873) );
  NAND2_X1 U964 ( .A1(n862), .A2(G103), .ZN(n863) );
  XNOR2_X1 U965 ( .A(KEYINPUT111), .B(n863), .ZN(n871) );
  NAND2_X1 U966 ( .A1(G115), .A2(n864), .ZN(n867) );
  NAND2_X1 U967 ( .A1(G127), .A2(n865), .ZN(n866) );
  NAND2_X1 U968 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U969 ( .A(KEYINPUT112), .B(n868), .Z(n869) );
  XNOR2_X1 U970 ( .A(KEYINPUT47), .B(n869), .ZN(n870) );
  NOR2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n872) );
  NAND2_X1 U972 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U973 ( .A(n874), .B(KEYINPUT113), .ZN(n922) );
  XNOR2_X1 U974 ( .A(n875), .B(n922), .ZN(n876) );
  XNOR2_X1 U975 ( .A(n877), .B(n876), .ZN(n882) );
  XNOR2_X1 U976 ( .A(G162), .B(n878), .ZN(n879) );
  XNOR2_X1 U977 ( .A(n879), .B(n915), .ZN(n880) );
  XOR2_X1 U978 ( .A(G160), .B(n880), .Z(n881) );
  XNOR2_X1 U979 ( .A(n882), .B(n881), .ZN(n883) );
  NOR2_X1 U980 ( .A1(G37), .A2(n883), .ZN(G395) );
  XOR2_X1 U981 ( .A(n884), .B(G286), .Z(n886) );
  XNOR2_X1 U982 ( .A(G171), .B(n967), .ZN(n885) );
  XNOR2_X1 U983 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n962), .B(n887), .ZN(n888) );
  NOR2_X1 U985 ( .A1(G37), .A2(n888), .ZN(G397) );
  XNOR2_X1 U986 ( .A(G1341), .B(G2454), .ZN(n889) );
  XNOR2_X1 U987 ( .A(n889), .B(G2430), .ZN(n890) );
  XNOR2_X1 U988 ( .A(n890), .B(G1348), .ZN(n896) );
  XOR2_X1 U989 ( .A(G2443), .B(G2427), .Z(n892) );
  XNOR2_X1 U990 ( .A(G2438), .B(G2446), .ZN(n891) );
  XNOR2_X1 U991 ( .A(n892), .B(n891), .ZN(n894) );
  XOR2_X1 U992 ( .A(G2451), .B(G2435), .Z(n893) );
  XNOR2_X1 U993 ( .A(n894), .B(n893), .ZN(n895) );
  XNOR2_X1 U994 ( .A(n896), .B(n895), .ZN(n897) );
  NAND2_X1 U995 ( .A1(n897), .A2(G14), .ZN(n898) );
  XNOR2_X1 U996 ( .A(KEYINPUT107), .B(n898), .ZN(n912) );
  NOR2_X1 U997 ( .A1(G227), .A2(G229), .ZN(n899) );
  XNOR2_X1 U998 ( .A(n899), .B(KEYINPUT49), .ZN(n900) );
  NOR2_X1 U999 ( .A1(n912), .A2(n900), .ZN(n901) );
  NAND2_X1 U1000 ( .A1(G319), .A2(n901), .ZN(n902) );
  XNOR2_X1 U1001 ( .A(KEYINPUT115), .B(n902), .ZN(n904) );
  NOR2_X1 U1002 ( .A1(G395), .A2(G397), .ZN(n903) );
  NAND2_X1 U1003 ( .A1(n904), .A2(n903), .ZN(G225) );
  XOR2_X1 U1004 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  INV_X1 U1006 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1007 ( .A1(n906), .A2(n905), .ZN(G325) );
  INV_X1 U1008 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1009 ( .A(n907), .B(KEYINPUT77), .Z(n908) );
  NOR2_X1 U1010 ( .A1(G860), .A2(n908), .ZN(n909) );
  XOR2_X1 U1011 ( .A(KEYINPUT78), .B(n909), .Z(n910) );
  XOR2_X1 U1012 ( .A(n911), .B(n910), .Z(G145) );
  XNOR2_X1 U1013 ( .A(n912), .B(KEYINPUT108), .ZN(G401) );
  NOR2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n921) );
  XNOR2_X1 U1015 ( .A(G160), .B(G2084), .ZN(n916) );
  NAND2_X1 U1016 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1018 ( .A(KEYINPUT117), .B(n919), .Z(n920) );
  NAND2_X1 U1019 ( .A1(n921), .A2(n920), .ZN(n935) );
  XOR2_X1 U1020 ( .A(G2072), .B(n922), .Z(n924) );
  XOR2_X1 U1021 ( .A(G164), .B(G2078), .Z(n923) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(KEYINPUT118), .B(n925), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(n926), .B(KEYINPUT50), .ZN(n933) );
  XOR2_X1 U1025 ( .A(G2090), .B(G162), .Z(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1027 ( .A(n929), .B(KEYINPUT51), .ZN(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1031 ( .A(KEYINPUT52), .B(n936), .ZN(n937) );
  XNOR2_X1 U1032 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n939) );
  NAND2_X1 U1033 ( .A1(n937), .A2(n939), .ZN(n938) );
  NAND2_X1 U1034 ( .A1(n938), .A2(G29), .ZN(n1021) );
  XNOR2_X1 U1035 ( .A(n939), .B(KEYINPUT121), .ZN(n959) );
  XNOR2_X1 U1036 ( .A(G2090), .B(G35), .ZN(n953) );
  XNOR2_X1 U1037 ( .A(G2072), .B(G33), .ZN(n941) );
  XNOR2_X1 U1038 ( .A(G1996), .B(G32), .ZN(n940) );
  NOR2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n947) );
  XOR2_X1 U1040 ( .A(G2067), .B(G26), .Z(n942) );
  NAND2_X1 U1041 ( .A1(n942), .A2(G28), .ZN(n945) );
  XNOR2_X1 U1042 ( .A(G25), .B(n943), .ZN(n944) );
  NOR2_X1 U1043 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n950) );
  XOR2_X1 U1045 ( .A(G27), .B(n948), .Z(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(KEYINPUT53), .B(n951), .ZN(n952) );
  NOR2_X1 U1048 ( .A1(n953), .A2(n952), .ZN(n957) );
  XOR2_X1 U1049 ( .A(KEYINPUT120), .B(G34), .Z(n955) );
  XNOR2_X1 U1050 ( .A(G2084), .B(KEYINPUT54), .ZN(n954) );
  XNOR2_X1 U1051 ( .A(n955), .B(n954), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(n959), .B(n958), .ZN(n960) );
  OR2_X1 U1054 ( .A1(G29), .A2(n960), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(G11), .A2(n961), .ZN(n1019) );
  XNOR2_X1 U1056 ( .A(G16), .B(KEYINPUT56), .ZN(n990) );
  XNOR2_X1 U1057 ( .A(G1341), .B(n962), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(n963), .B(KEYINPUT126), .ZN(n988) );
  XOR2_X1 U1059 ( .A(G1966), .B(G168), .Z(n964) );
  NOR2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(KEYINPUT57), .B(n966), .ZN(n986) );
  XNOR2_X1 U1062 ( .A(G1348), .B(n967), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(n968), .B(KEYINPUT122), .ZN(n979) );
  XNOR2_X1 U1064 ( .A(G1971), .B(G166), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n976) );
  XNOR2_X1 U1066 ( .A(G1956), .B(n971), .ZN(n974) );
  XNOR2_X1 U1067 ( .A(n972), .B(KEYINPUT123), .ZN(n973) );
  NAND2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n975) );
  NOR2_X1 U1069 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1070 ( .A(n977), .B(KEYINPUT124), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(G171), .B(G1961), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(KEYINPUT125), .B(n984), .ZN(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n1017) );
  INV_X1 U1079 ( .A(G16), .ZN(n1015) );
  XNOR2_X1 U1080 ( .A(G5), .B(n991), .ZN(n1005) );
  XNOR2_X1 U1081 ( .A(G1348), .B(KEYINPUT59), .ZN(n992) );
  XNOR2_X1 U1082 ( .A(n992), .B(G4), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(G1981), .B(G6), .ZN(n994) );
  XNOR2_X1 U1084 ( .A(G1341), .B(G19), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(G20), .B(n997), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(KEYINPUT127), .B(n998), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1090 ( .A(KEYINPUT60), .B(n1001), .Z(n1003) );
  XNOR2_X1 U1091 ( .A(G1966), .B(G21), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1012) );
  XNOR2_X1 U1094 ( .A(G1971), .B(G22), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(G24), .B(G1986), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  XOR2_X1 U1097 ( .A(G1976), .B(G23), .Z(n1008) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(KEYINPUT58), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(KEYINPUT61), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1105 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1022), .Z(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

