//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n555, new_n557, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n611, new_n612, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  INV_X1    g030(.A(new_n452), .ZN(new_n456));
  AOI22_X1  g031(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT65), .Z(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n462), .B1(new_n459), .B2(KEYINPUT66), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n461), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n471), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(new_n467), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n470), .A2(new_n473), .ZN(G160));
  AOI21_X1  g049(.A(new_n467), .B1(new_n463), .B2(new_n465), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n467), .A2(G112), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n468), .A2(KEYINPUT67), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n463), .B2(new_n465), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n479), .B1(new_n484), .B2(G136), .ZN(G162));
  NAND2_X1  g060(.A1(new_n475), .A2(G126), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT68), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT69), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n488), .B1(new_n467), .B2(G114), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n490), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n489), .A2(new_n491), .A3(new_n492), .A4(G2104), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT70), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n471), .A2(G138), .A3(new_n467), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  AND2_X1   g071(.A1(KEYINPUT4), .A2(G138), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n495), .A2(new_n496), .B1(new_n481), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n487), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  AND2_X1   g075(.A1(KEYINPUT6), .A2(G651), .ZN(new_n501));
  NOR2_X1   g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  OAI211_X1 g077(.A(G50), .B(G543), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n506), .A2(KEYINPUT71), .A3(G50), .A4(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g087(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g089(.A1(G75), .A2(G543), .ZN(new_n515));
  OAI21_X1  g090(.A(G651), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n512), .A2(new_n513), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n517), .A2(G88), .A3(new_n506), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n508), .A2(new_n516), .A3(new_n518), .ZN(G303));
  INV_X1    g094(.A(G303), .ZN(G166));
  OAI21_X1  g095(.A(G543), .B1(new_n501), .B2(new_n502), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT73), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n523));
  OAI211_X1 g098(.A(new_n523), .B(G543), .C1(new_n501), .C2(new_n502), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n525), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  AND3_X1   g105(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n531));
  AOI21_X1  g106(.A(G543), .B1(KEYINPUT72), .B2(KEYINPUT5), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n531), .A2(new_n532), .B1(new_n501), .B2(new_n502), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n527), .B(new_n529), .C1(new_n530), .C2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n526), .A2(new_n534), .ZN(G168));
  AOI22_X1  g110(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G651), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n525), .A2(G52), .ZN(new_n539));
  INV_X1    g114(.A(new_n533), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G90), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(G68), .A2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n531), .A2(new_n532), .ZN(new_n545));
  INV_X1    g120(.A(G56), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n537), .B1(new_n547), .B2(KEYINPUT74), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n548), .B1(KEYINPUT74), .B2(new_n547), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n525), .A2(G43), .B1(G81), .B2(new_n540), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G860), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT75), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  XOR2_X1   g131(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n557));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n555), .A2(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n545), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n563), .A2(G651), .B1(new_n540), .B2(G91), .ZN(new_n564));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  OR3_X1    g140(.A1(new_n521), .A2(KEYINPUT9), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT9), .B1(new_n521), .B2(new_n565), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n564), .A2(new_n568), .ZN(G299));
  INV_X1    g144(.A(KEYINPUT77), .ZN(new_n570));
  NOR3_X1   g145(.A1(new_n526), .A2(new_n570), .A3(new_n534), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n534), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n525), .A2(G51), .ZN(new_n574));
  AOI21_X1  g149(.A(KEYINPUT77), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G286));
  INV_X1    g153(.A(new_n521), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G49), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n517), .A2(G87), .A3(new_n506), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(G288));
  AOI22_X1  g158(.A1(new_n540), .A2(G86), .B1(new_n579), .B2(G48), .ZN(new_n584));
  OAI21_X1  g159(.A(G61), .B1(new_n531), .B2(new_n532), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g162(.A(KEYINPUT78), .B1(new_n587), .B2(G651), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n589));
  AOI211_X1 g164(.A(new_n589), .B(new_n537), .C1(new_n585), .C2(new_n586), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n584), .B1(new_n588), .B2(new_n590), .ZN(G305));
  NAND2_X1  g166(.A1(G72), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G60), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n545), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(new_n540), .B2(G85), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n525), .A2(G47), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n533), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n525), .A2(G54), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(new_n537), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n601), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n598), .B1(new_n606), .B2(G868), .ZN(G284));
  OAI21_X1  g182(.A(new_n598), .B1(new_n606), .B2(G868), .ZN(G321));
  AND2_X1   g183(.A1(new_n564), .A2(new_n568), .ZN(new_n609));
  OAI21_X1  g184(.A(KEYINPUT79), .B1(new_n609), .B2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n577), .A2(new_n611), .ZN(new_n612));
  MUX2_X1   g187(.A(new_n610), .B(KEYINPUT79), .S(new_n612), .Z(G297));
  MUX2_X1   g188(.A(new_n610), .B(KEYINPUT79), .S(new_n612), .Z(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n606), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n551), .A2(new_n611), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n605), .A2(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n611), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n484), .A2(G135), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n475), .A2(G123), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n467), .A2(G111), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n621), .B(new_n622), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT80), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(G2096), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(G2096), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT12), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT13), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2100), .ZN(new_n633));
  NAND3_X1  g208(.A1(new_n628), .A2(new_n629), .A3(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(new_n639), .A3(KEYINPUT14), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n640), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2451), .B(G2454), .Z(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(G14), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n644), .A2(new_n647), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n649), .A2(new_n650), .ZN(G401));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT82), .ZN(new_n653));
  XOR2_X1   g228(.A(G2072), .B(G2078), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n653), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT18), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n656), .B(KEYINPUT83), .ZN(new_n659));
  OAI21_X1  g234(.A(KEYINPUT17), .B1(new_n653), .B2(new_n659), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n660), .A2(new_n654), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n653), .A2(new_n659), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n660), .B2(new_n654), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n658), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2100), .ZN(new_n665));
  XNOR2_X1  g240(.A(KEYINPUT84), .B(G2096), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1991), .B(G1996), .Z(new_n668));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT85), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT86), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n671), .A2(KEYINPUT86), .A3(new_n672), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT19), .Z(new_n678));
  NAND3_X1  g253(.A1(new_n675), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT20), .ZN(new_n680));
  OR2_X1    g255(.A1(new_n671), .A2(new_n672), .ZN(new_n681));
  INV_X1    g256(.A(new_n678), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n681), .A2(new_n673), .A3(new_n682), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n680), .B(new_n683), .C1(new_n682), .C2(new_n681), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n684), .A2(new_n686), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n668), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n689), .ZN(new_n691));
  INV_X1    g266(.A(new_n668), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n691), .A2(new_n692), .A3(new_n687), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  AND3_X1   g269(.A1(new_n690), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n694), .B1(new_n690), .B2(new_n693), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(G229));
  MUX2_X1   g272(.A(G24), .B(G290), .S(G16), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1986), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n484), .A2(G131), .ZN(new_n700));
  OAI21_X1  g275(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n701));
  INV_X1    g276(.A(G107), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(G2105), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT87), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n704), .ZN(new_n706));
  AOI22_X1  g281(.A1(new_n705), .A2(new_n706), .B1(G119), .B2(new_n475), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n700), .A2(new_n707), .ZN(new_n708));
  MUX2_X1   g283(.A(G25), .B(new_n708), .S(G29), .Z(new_n709));
  XOR2_X1   g284(.A(KEYINPUT35), .B(G1991), .Z(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n709), .B(new_n711), .ZN(new_n712));
  AOI211_X1 g287(.A(new_n699), .B(new_n712), .C1(KEYINPUT89), .C2(KEYINPUT36), .ZN(new_n713));
  NOR2_X1   g288(.A1(G16), .A2(G23), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT88), .Z(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(G288), .B2(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT33), .ZN(new_n718));
  INV_X1    g293(.A(G1976), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n716), .A2(G6), .ZN(new_n721));
  INV_X1    g296(.A(G305), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(new_n716), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT32), .B(G1981), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n716), .A2(G22), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G166), .B2(new_n716), .ZN(new_n727));
  INV_X1    g302(.A(G1971), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n720), .A2(new_n725), .A3(new_n729), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(KEYINPUT34), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n713), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(KEYINPUT34), .B2(new_n730), .ZN(new_n733));
  OR3_X1    g308(.A1(new_n733), .A2(KEYINPUT89), .A3(KEYINPUT36), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(KEYINPUT89), .B2(KEYINPUT36), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n716), .A2(G21), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G168), .B2(new_n716), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G1966), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT31), .B(G11), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT93), .B(G28), .Z(new_n740));
  AOI21_X1  g315(.A(G29), .B1(new_n740), .B2(KEYINPUT30), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(KEYINPUT30), .B2(new_n740), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n738), .A2(new_n739), .A3(new_n742), .ZN(new_n743));
  NOR2_X1   g318(.A1(G171), .A2(new_n716), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G5), .B2(new_n716), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n743), .B1(new_n746), .B2(G1961), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n737), .A2(G1966), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT94), .ZN(new_n749));
  INV_X1    g324(.A(G29), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n747), .B(new_n749), .C1(new_n750), .C2(new_n627), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT95), .Z(new_n752));
  NOR2_X1   g327(.A1(new_n606), .A2(new_n716), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G4), .B2(new_n716), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT90), .B(G1348), .Z(new_n755));
  NOR2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(G1961), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(new_n745), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n750), .A2(G33), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n760), .A2(new_n467), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT25), .ZN(new_n763));
  AOI211_X1 g338(.A(new_n761), .B(new_n763), .C1(new_n484), .C2(G139), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n759), .B1(new_n764), .B2(new_n750), .ZN(new_n765));
  INV_X1    g340(.A(G2078), .ZN(new_n766));
  NAND2_X1  g341(.A1(G164), .A2(G29), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G27), .B2(G29), .ZN(new_n768));
  OAI221_X1 g343(.A(new_n758), .B1(G2072), .B2(new_n765), .C1(new_n766), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n754), .A2(new_n755), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n766), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n765), .A2(G2072), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n484), .A2(G141), .ZN(new_n774));
  NAND3_X1  g349(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT26), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  AOI22_X1  g353(.A1(new_n777), .A2(new_n778), .B1(G105), .B2(new_n460), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n475), .A2(G129), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n774), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT92), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  MUX2_X1   g359(.A(G32), .B(new_n784), .S(G29), .Z(new_n785));
  XOR2_X1   g360(.A(KEYINPUT27), .B(G1996), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  AND2_X1   g362(.A1(new_n549), .A2(new_n550), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n788), .A2(new_n716), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n716), .B2(G19), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(G1341), .ZN(new_n792));
  INV_X1    g367(.A(G2084), .ZN(new_n793));
  AND2_X1   g368(.A1(KEYINPUT24), .A2(G34), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n750), .B1(KEYINPUT24), .B2(G34), .ZN(new_n795));
  OAI22_X1  g370(.A1(G160), .A2(new_n750), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT91), .Z(new_n797));
  AOI22_X1  g372(.A1(new_n791), .A2(G1341), .B1(new_n793), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n750), .A2(G26), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT28), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n484), .A2(G140), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n802));
  INV_X1    g377(.A(G116), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(G2105), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n475), .B2(G128), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n800), .B1(new_n806), .B2(G29), .ZN(new_n807));
  INV_X1    g382(.A(G2067), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n750), .A2(G35), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G162), .B2(new_n750), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT29), .B(G2090), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n716), .A2(G20), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT23), .Z(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G299), .B2(G16), .ZN(new_n817));
  INV_X1    g392(.A(G1956), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n797), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(G2084), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n792), .A2(new_n798), .A3(new_n814), .A4(new_n821), .ZN(new_n822));
  NOR4_X1   g397(.A1(new_n769), .A2(new_n773), .A3(new_n787), .A4(new_n822), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n734), .A2(new_n735), .A3(new_n752), .A4(new_n823), .ZN(G150));
  INV_X1    g399(.A(G150), .ZN(G311));
  INV_X1    g400(.A(G67), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(new_n512), .B2(new_n513), .ZN(new_n827));
  NAND2_X1  g402(.A1(G80), .A2(G543), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  OAI21_X1  g404(.A(KEYINPUT96), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT96), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n831), .B(new_n828), .C1(new_n545), .C2(new_n826), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n830), .A2(new_n832), .A3(G651), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT98), .ZN(new_n834));
  XNOR2_X1  g409(.A(KEYINPUT97), .B(G55), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n523), .B1(new_n506), .B2(G543), .ZN(new_n836));
  INV_X1    g411(.A(new_n524), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(G93), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n533), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n834), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n835), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n843), .B1(new_n522), .B2(new_n524), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n844), .A2(KEYINPUT98), .A3(new_n840), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n833), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT99), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n848), .B(new_n833), .C1(new_n842), .C2(new_n845), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n847), .A2(new_n788), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n846), .A2(KEYINPUT99), .A3(new_n551), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT38), .Z(new_n853));
  NOR2_X1   g428(.A1(new_n605), .A2(new_n615), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n856));
  AOI21_X1  g431(.A(G860), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n856), .B2(new_n855), .ZN(new_n858));
  INV_X1    g433(.A(new_n833), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n838), .A2(new_n834), .A3(new_n841), .ZN(new_n860));
  OAI21_X1  g435(.A(KEYINPUT98), .B1(new_n844), .B2(new_n840), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n859), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n862), .A2(new_n552), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT37), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n858), .A2(new_n864), .ZN(G145));
  XOR2_X1   g440(.A(G162), .B(G160), .Z(new_n866));
  NAND2_X1  g441(.A1(new_n784), .A2(new_n764), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n764), .A2(new_n782), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n806), .B(new_n499), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n871), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n867), .A2(new_n873), .A3(new_n869), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n708), .B(new_n631), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n475), .A2(G130), .ZN(new_n877));
  OR2_X1    g452(.A1(G106), .A2(G2105), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n878), .B(G2104), .C1(G118), .C2(new_n467), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n880), .B1(new_n484), .B2(G142), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n876), .B(new_n881), .Z(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(KEYINPUT100), .B1(new_n875), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n872), .A3(new_n874), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(new_n627), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n627), .B1(new_n884), .B2(new_n885), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n866), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n888), .ZN(new_n890));
  INV_X1    g465(.A(new_n866), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(new_n886), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(G37), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n889), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g470(.A1(new_n846), .A2(new_n611), .ZN(new_n896));
  AOI21_X1  g471(.A(G288), .B1(new_n595), .B2(new_n596), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n595), .A2(G288), .A3(new_n596), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n901));
  NAND2_X1  g476(.A1(G303), .A2(new_n901), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n508), .A2(KEYINPUT102), .A3(new_n516), .A4(new_n518), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n902), .A2(G305), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(G305), .B1(new_n902), .B2(new_n903), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n900), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n902), .A2(new_n903), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n722), .ZN(new_n908));
  INV_X1    g483(.A(new_n899), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n909), .A2(new_n897), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n902), .A2(G305), .A3(new_n903), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n908), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n906), .A2(new_n912), .A3(KEYINPUT103), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT103), .B1(new_n906), .B2(new_n912), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n915), .A2(KEYINPUT42), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n906), .A2(new_n912), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n917), .A2(KEYINPUT42), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n916), .B1(KEYINPUT104), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(KEYINPUT104), .B2(new_n916), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n852), .B(new_n618), .ZN(new_n921));
  XOR2_X1   g496(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n922));
  NOR2_X1   g497(.A1(new_n605), .A2(G299), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n604), .A2(new_n602), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n609), .B1(new_n601), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n922), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n605), .A2(G299), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(new_n609), .A3(new_n601), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n926), .B1(new_n929), .B2(KEYINPUT41), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n921), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n929), .B2(new_n921), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n920), .B(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n896), .B1(new_n933), .B2(new_n611), .ZN(G295));
  OAI21_X1  g509(.A(new_n896), .B1(new_n933), .B2(new_n611), .ZN(G331));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT106), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n923), .A2(new_n925), .ZN(new_n938));
  OAI21_X1  g513(.A(G171), .B1(new_n571), .B2(new_n575), .ZN(new_n939));
  INV_X1    g514(.A(G168), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(G301), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n850), .A2(new_n942), .A3(new_n851), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n942), .B1(new_n850), .B2(new_n851), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n938), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n939), .A2(new_n941), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n849), .A2(new_n788), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n862), .A2(new_n848), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n851), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n946), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n850), .A2(new_n942), .A3(new_n851), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT41), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n929), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n927), .A2(new_n928), .A3(new_n922), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n951), .A2(new_n952), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n945), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n915), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n937), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AOI211_X1 g534(.A(KEYINPUT106), .B(new_n915), .C1(new_n945), .C2(new_n956), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n951), .A2(new_n930), .A3(new_n952), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT105), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n951), .A2(new_n930), .A3(new_n964), .A4(new_n952), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n963), .A2(new_n915), .A3(new_n965), .A4(new_n945), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n966), .A2(new_n893), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n961), .A2(new_n967), .A3(KEYINPUT43), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n966), .A2(new_n893), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n945), .A2(new_n965), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n915), .B1(new_n971), .B2(new_n963), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n969), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n936), .B1(new_n968), .B2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n961), .A2(new_n967), .A3(new_n969), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT43), .B1(new_n970), .B2(new_n972), .ZN(new_n976));
  AOI21_X1  g551(.A(KEYINPUT44), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT107), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n954), .A2(new_n955), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n943), .A2(new_n944), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n929), .B1(new_n951), .B2(new_n952), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n958), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT106), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n957), .A2(new_n937), .A3(new_n958), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n985), .A2(new_n969), .A3(new_n970), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n971), .A2(new_n963), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n958), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT43), .B1(new_n967), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT44), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n985), .A2(KEYINPUT43), .A3(new_n970), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n969), .B1(new_n967), .B2(new_n988), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n936), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT107), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n990), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n978), .A2(new_n995), .ZN(G397));
  XNOR2_X1  g571(.A(new_n806), .B(new_n808), .ZN(new_n997));
  INV_X1    g572(.A(G1384), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT45), .B1(new_n499), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT108), .B(G40), .ZN(new_n1000));
  NOR3_X1   g575(.A1(new_n470), .A2(new_n473), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n997), .A2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1003), .A2(KEYINPUT109), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n1003), .A2(KEYINPUT109), .ZN(new_n1005));
  INV_X1    g580(.A(G1996), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n784), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n782), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1002), .B1(G1996), .B2(new_n1008), .ZN(new_n1009));
  AOI211_X1 g584(.A(new_n1004), .B(new_n1005), .C1(new_n1007), .C2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n708), .B(new_n710), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1010), .B1(new_n1002), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1002), .ZN(new_n1013));
  XNOR2_X1  g588(.A(G290), .B(G1986), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OR2_X1    g590(.A1(G305), .A2(G1981), .ZN(new_n1016));
  INV_X1    g591(.A(new_n584), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n537), .B1(new_n585), .B2(new_n586), .ZN(new_n1018));
  OAI21_X1  g593(.A(G1981), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT49), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1016), .A2(KEYINPUT49), .A3(new_n1019), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n499), .A2(new_n998), .A3(new_n1001), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1022), .A2(G8), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G288), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(G1976), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n1027), .B(KEYINPUT112), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1028), .A2(new_n1024), .A3(G8), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT52), .ZN(new_n1030));
  AOI21_X1  g605(.A(KEYINPUT52), .B1(G288), .B2(new_n719), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1028), .A2(new_n1024), .A3(G8), .A4(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1025), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT113), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT113), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1025), .A2(new_n1030), .A3(new_n1035), .A4(new_n1032), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n499), .A2(new_n998), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT50), .ZN(new_n1039));
  AND2_X1   g614(.A1(new_n494), .A2(new_n498), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1384), .B1(new_n1040), .B2(new_n487), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1039), .A2(new_n1043), .A3(new_n1001), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT110), .B1(new_n1044), .B2(G2090), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1001), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n999), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n998), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n728), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1046), .B1(new_n1038), .B2(KEYINPUT50), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT110), .ZN(new_n1052));
  INV_X1    g627(.A(G2090), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1043), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1045), .A2(new_n1050), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G8), .ZN(new_n1056));
  NOR2_X1   g631(.A1(G166), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1058), .A2(KEYINPUT111), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1058), .A2(KEYINPUT111), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1057), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1055), .A2(G8), .A3(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1037), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1024), .A2(G8), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1025), .A2(new_n719), .A3(new_n1026), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1065), .B1(new_n1066), .B2(new_n1016), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT123), .B(KEYINPUT54), .Z(new_n1069));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1070), .B1(new_n1049), .B2(G2078), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT114), .B1(new_n999), .B2(new_n1046), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT114), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1074), .B(new_n1001), .C1(new_n1041), .C2(KEYINPUT45), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1070), .A2(G2078), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1073), .A2(new_n1048), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1044), .A2(new_n757), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT124), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1077), .A2(KEYINPUT124), .A3(new_n1078), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1072), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(G301), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT45), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1038), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1076), .A2(G40), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n472), .A2(KEYINPUT125), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1088), .A2(new_n467), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n472), .A2(KEYINPUT125), .ZN(new_n1090));
  AOI211_X1 g665(.A(new_n470), .B(new_n1087), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1086), .A2(new_n1048), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1071), .A2(new_n1078), .A3(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(G171), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1069), .B1(new_n1084), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT61), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n1097), .B(G2072), .ZN(new_n1098));
  AND4_X1   g673(.A1(new_n1086), .A2(new_n1001), .A3(new_n1048), .A4(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(G1956), .B1(new_n1051), .B2(new_n1043), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n609), .B(KEYINPUT57), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1099), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1044), .A2(new_n818), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1047), .A2(new_n1048), .A3(new_n1098), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1101), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1096), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1102), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1104), .A2(new_n1105), .A3(new_n1101), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(new_n1109), .A3(KEYINPUT61), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1086), .A2(new_n1006), .A3(new_n1001), .A4(new_n1048), .ZN(new_n1111));
  XOR2_X1   g686(.A(KEYINPUT58), .B(G1341), .Z(new_n1112));
  NAND2_X1  g687(.A1(new_n1024), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n788), .A2(KEYINPUT119), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT59), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n1118));
  AOI211_X1 g693(.A(new_n1118), .B(new_n1115), .C1(new_n1111), .C2(new_n1113), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1107), .A2(new_n1110), .A3(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1024), .A2(G2067), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1122), .B1(new_n1044), .B2(new_n755), .ZN(new_n1123));
  OR2_X1    g698(.A1(new_n1123), .A2(KEYINPUT60), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT120), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(KEYINPUT60), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1125), .B1(new_n1126), .B2(new_n606), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT60), .ZN(new_n1128));
  AOI211_X1 g703(.A(new_n1128), .B(new_n1122), .C1(new_n1044), .C2(new_n755), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT121), .B1(new_n1129), .B2(new_n605), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1126), .A2(new_n1131), .A3(new_n606), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1129), .A2(KEYINPUT120), .A3(new_n605), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1127), .A2(new_n1130), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1121), .B1(new_n1124), .B2(new_n1134), .ZN(new_n1135));
  OR2_X1    g710(.A1(new_n1123), .A2(new_n605), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1103), .B1(new_n1136), .B2(new_n1108), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1095), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1044), .A2(G2090), .ZN(new_n1139));
  AOI21_X1  g714(.A(G1971), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1140));
  OAI21_X1  g715(.A(G8), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1062), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1033), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(new_n1063), .ZN(new_n1144));
  AOI211_X1 g719(.A(KEYINPUT50), .B(G1384), .C1(new_n1040), .C2(new_n487), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1042), .B1(new_n499), .B2(new_n998), .ZN(new_n1146));
  XOR2_X1   g721(.A(KEYINPUT115), .B(G2084), .Z(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  NOR4_X1   g723(.A1(new_n1145), .A2(new_n1146), .A3(new_n1046), .A4(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1073), .A2(new_n1048), .A3(new_n1075), .ZN(new_n1150));
  INV_X1    g725(.A(G1966), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1149), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1152), .A2(new_n1056), .A3(G168), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT51), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1056), .B1(KEYINPUT122), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1149), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1155), .B1(new_n1158), .B2(new_n940), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1154), .A2(KEYINPUT122), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1153), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1155), .ZN(new_n1162));
  AOI211_X1 g737(.A(new_n1162), .B(new_n1160), .C1(new_n1152), .C2(G168), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1144), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1083), .A2(G301), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1093), .A2(G171), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1166), .A2(KEYINPUT54), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1165), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1068), .B1(new_n1138), .B2(new_n1169), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1144), .A2(new_n1083), .A3(G301), .ZN(new_n1171));
  AOI21_X1  g746(.A(KEYINPUT62), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1158), .A2(G8), .A3(new_n940), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1162), .B1(new_n1152), .B2(G168), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1160), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1173), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT62), .ZN(new_n1177));
  NOR3_X1   g752(.A1(new_n1176), .A2(new_n1177), .A3(new_n1163), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1171), .B1(new_n1172), .B2(new_n1178), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1152), .A2(new_n1056), .A3(G286), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1180), .A2(new_n1143), .A3(new_n1063), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(KEYINPUT116), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT63), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT116), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1180), .A2(new_n1143), .A3(new_n1063), .A4(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1182), .A2(new_n1183), .A3(new_n1185), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1062), .B1(new_n1055), .B2(G8), .ZN(new_n1187));
  OAI21_X1  g762(.A(KEYINPUT117), .B1(new_n1037), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT117), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1034), .A2(new_n1036), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1055), .A2(G8), .ZN(new_n1191));
  OAI211_X1 g766(.A(new_n1189), .B(new_n1190), .C1(new_n1191), .C2(new_n1062), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1180), .A2(new_n1063), .A3(KEYINPUT63), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1188), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1186), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1179), .A2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1015), .B1(new_n1170), .B2(new_n1196), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1010), .A2(new_n710), .A3(new_n700), .A4(new_n707), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n801), .A2(new_n808), .A3(new_n805), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1002), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n1201));
  AND2_X1   g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1002), .B1(new_n997), .B2(new_n1008), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT46), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1013), .A2(new_n1006), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1204), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1207), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1208), .B(KEYINPUT47), .ZN(new_n1209));
  NOR3_X1   g784(.A1(new_n1002), .A2(G1986), .A3(G290), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n1210), .B(KEYINPUT48), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1209), .B1(new_n1012), .B2(new_n1211), .ZN(new_n1212));
  NOR3_X1   g787(.A1(new_n1202), .A2(new_n1203), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1197), .A2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g789(.A(new_n457), .B1(new_n649), .B2(new_n650), .ZN(new_n1216));
  NOR2_X1   g790(.A1(G227), .A2(new_n1216), .ZN(new_n1217));
  OAI21_X1  g791(.A(new_n1217), .B1(new_n695), .B2(new_n696), .ZN(new_n1218));
  NAND2_X1  g792(.A1(new_n1218), .A2(KEYINPUT127), .ZN(new_n1219));
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n1220));
  OAI211_X1 g794(.A(new_n1217), .B(new_n1220), .C1(new_n695), .C2(new_n696), .ZN(new_n1221));
  NAND2_X1  g795(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  OAI211_X1 g796(.A(new_n894), .B(new_n1222), .C1(new_n992), .C2(new_n991), .ZN(G225));
  INV_X1    g797(.A(G225), .ZN(G308));
endmodule


