

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U556 ( .A(KEYINPUT23), .B(n528), .Z(n531) );
  NOR2_X1 U557 ( .A1(n813), .A2(n800), .ZN(n522) );
  XOR2_X1 U558 ( .A(n740), .B(n739), .Z(n523) );
  INV_X1 U559 ( .A(n774), .ZN(n757) );
  NOR2_X2 U560 ( .A1(G2105), .A2(G2104), .ZN(n524) );
  OR2_X1 U561 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U562 ( .A(n534), .B(KEYINPUT65), .ZN(G160) );
  XOR2_X2 U563 ( .A(KEYINPUT17), .B(n524), .Z(n879) );
  NAND2_X1 U564 ( .A1(G137), .A2(n879), .ZN(n526) );
  INV_X1 U565 ( .A(G2105), .ZN(n527) );
  NOR2_X1 U566 ( .A1(G2104), .A2(n527), .ZN(n876) );
  NAND2_X1 U567 ( .A1(G125), .A2(n876), .ZN(n525) );
  NAND2_X1 U568 ( .A1(n526), .A2(n525), .ZN(n533) );
  AND2_X2 U569 ( .A1(n527), .A2(G2104), .ZN(n880) );
  NAND2_X1 U570 ( .A1(G101), .A2(n880), .ZN(n528) );
  AND2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n875) );
  NAND2_X1 U572 ( .A1(G113), .A2(n875), .ZN(n529) );
  XNOR2_X1 U573 ( .A(n529), .B(KEYINPUT66), .ZN(n530) );
  NAND2_X1 U574 ( .A1(n531), .A2(n530), .ZN(n532) );
  INV_X1 U575 ( .A(G651), .ZN(n538) );
  NOR2_X1 U576 ( .A1(G543), .A2(n538), .ZN(n535) );
  XOR2_X1 U577 ( .A(KEYINPUT1), .B(n535), .Z(n644) );
  NAND2_X1 U578 ( .A1(G60), .A2(n644), .ZN(n537) );
  NOR2_X1 U579 ( .A1(G651), .A2(G543), .ZN(n645) );
  NAND2_X1 U580 ( .A1(G85), .A2(n645), .ZN(n536) );
  NAND2_X1 U581 ( .A1(n537), .A2(n536), .ZN(n543) );
  XOR2_X1 U582 ( .A(KEYINPUT0), .B(G543), .Z(n634) );
  NOR2_X1 U583 ( .A1(n634), .A2(n538), .ZN(n648) );
  NAND2_X1 U584 ( .A1(n648), .A2(G72), .ZN(n541) );
  NOR2_X1 U585 ( .A1(G651), .A2(n634), .ZN(n539) );
  XNOR2_X1 U586 ( .A(KEYINPUT64), .B(n539), .ZN(n652) );
  NAND2_X1 U587 ( .A1(G47), .A2(n652), .ZN(n540) );
  NAND2_X1 U588 ( .A1(n541), .A2(n540), .ZN(n542) );
  OR2_X1 U589 ( .A1(n543), .A2(n542), .ZN(G290) );
  NAND2_X1 U590 ( .A1(G52), .A2(n652), .ZN(n544) );
  XNOR2_X1 U591 ( .A(KEYINPUT67), .B(n544), .ZN(n552) );
  NAND2_X1 U592 ( .A1(G90), .A2(n645), .ZN(n546) );
  NAND2_X1 U593 ( .A1(G77), .A2(n648), .ZN(n545) );
  NAND2_X1 U594 ( .A1(n546), .A2(n545), .ZN(n548) );
  XNOR2_X1 U595 ( .A(KEYINPUT68), .B(KEYINPUT9), .ZN(n547) );
  XNOR2_X1 U596 ( .A(n548), .B(n547), .ZN(n550) );
  NAND2_X1 U597 ( .A1(G64), .A2(n644), .ZN(n549) );
  NAND2_X1 U598 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U599 ( .A1(n552), .A2(n551), .ZN(G171) );
  AND2_X1 U600 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U601 ( .A(G57), .ZN(G237) );
  INV_X1 U602 ( .A(G132), .ZN(G219) );
  INV_X1 U603 ( .A(G82), .ZN(G220) );
  NAND2_X1 U604 ( .A1(n875), .A2(G114), .ZN(n555) );
  NAND2_X1 U605 ( .A1(n879), .A2(G138), .ZN(n553) );
  XOR2_X1 U606 ( .A(KEYINPUT81), .B(n553), .Z(n554) );
  NAND2_X1 U607 ( .A1(n555), .A2(n554), .ZN(n559) );
  NAND2_X1 U608 ( .A1(G102), .A2(n880), .ZN(n557) );
  NAND2_X1 U609 ( .A1(G126), .A2(n876), .ZN(n556) );
  NAND2_X1 U610 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U611 ( .A1(n559), .A2(n558), .ZN(n679) );
  BUF_X1 U612 ( .A(n679), .Z(G164) );
  NAND2_X1 U613 ( .A1(n644), .A2(G63), .ZN(n561) );
  NAND2_X1 U614 ( .A1(G51), .A2(n652), .ZN(n560) );
  NAND2_X1 U615 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U616 ( .A(KEYINPUT6), .B(n562), .ZN(n569) );
  NAND2_X1 U617 ( .A1(G89), .A2(n645), .ZN(n563) );
  XNOR2_X1 U618 ( .A(n563), .B(KEYINPUT4), .ZN(n564) );
  XNOR2_X1 U619 ( .A(n564), .B(KEYINPUT72), .ZN(n566) );
  NAND2_X1 U620 ( .A1(G76), .A2(n648), .ZN(n565) );
  NAND2_X1 U621 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U622 ( .A(n567), .B(KEYINPUT5), .Z(n568) );
  NOR2_X1 U623 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U624 ( .A(KEYINPUT7), .B(n570), .Z(n571) );
  XOR2_X1 U625 ( .A(KEYINPUT73), .B(n571), .Z(G168) );
  XOR2_X1 U626 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U627 ( .A1(G7), .A2(G661), .ZN(n572) );
  XNOR2_X1 U628 ( .A(n572), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U629 ( .A(G223), .ZN(n823) );
  NAND2_X1 U630 ( .A1(n823), .A2(G567), .ZN(n573) );
  XOR2_X1 U631 ( .A(KEYINPUT11), .B(n573), .Z(G234) );
  NAND2_X1 U632 ( .A1(G56), .A2(n644), .ZN(n574) );
  XOR2_X1 U633 ( .A(KEYINPUT14), .B(n574), .Z(n580) );
  NAND2_X1 U634 ( .A1(n645), .A2(G81), .ZN(n575) );
  XNOR2_X1 U635 ( .A(n575), .B(KEYINPUT12), .ZN(n577) );
  NAND2_X1 U636 ( .A1(G68), .A2(n648), .ZN(n576) );
  NAND2_X1 U637 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U638 ( .A(KEYINPUT13), .B(n578), .Z(n579) );
  NOR2_X1 U639 ( .A1(n580), .A2(n579), .ZN(n582) );
  NAND2_X1 U640 ( .A1(G43), .A2(n652), .ZN(n581) );
  NAND2_X1 U641 ( .A1(n582), .A2(n581), .ZN(n950) );
  INV_X1 U642 ( .A(G860), .ZN(n604) );
  OR2_X1 U643 ( .A1(n950), .A2(n604), .ZN(G153) );
  INV_X1 U644 ( .A(G171), .ZN(G301) );
  NAND2_X1 U645 ( .A1(G66), .A2(n644), .ZN(n584) );
  NAND2_X1 U646 ( .A1(G92), .A2(n645), .ZN(n583) );
  NAND2_X1 U647 ( .A1(n584), .A2(n583), .ZN(n588) );
  NAND2_X1 U648 ( .A1(n648), .A2(G79), .ZN(n586) );
  NAND2_X1 U649 ( .A1(G54), .A2(n652), .ZN(n585) );
  NAND2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U651 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U652 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n589) );
  XNOR2_X1 U653 ( .A(n590), .B(n589), .ZN(n591) );
  XOR2_X1 U654 ( .A(KEYINPUT15), .B(n591), .Z(n954) );
  NOR2_X1 U655 ( .A1(n954), .A2(G868), .ZN(n593) );
  INV_X1 U656 ( .A(G868), .ZN(n663) );
  NOR2_X1 U657 ( .A1(n663), .A2(G301), .ZN(n592) );
  NOR2_X1 U658 ( .A1(n593), .A2(n592), .ZN(G284) );
  NAND2_X1 U659 ( .A1(G91), .A2(n645), .ZN(n595) );
  NAND2_X1 U660 ( .A1(G78), .A2(n648), .ZN(n594) );
  NAND2_X1 U661 ( .A1(n595), .A2(n594), .ZN(n598) );
  NAND2_X1 U662 ( .A1(G65), .A2(n644), .ZN(n596) );
  XNOR2_X1 U663 ( .A(KEYINPUT69), .B(n596), .ZN(n597) );
  NOR2_X1 U664 ( .A1(n598), .A2(n597), .ZN(n600) );
  NAND2_X1 U665 ( .A1(G53), .A2(n652), .ZN(n599) );
  NAND2_X1 U666 ( .A1(n600), .A2(n599), .ZN(G299) );
  NOR2_X1 U667 ( .A1(G286), .A2(n663), .ZN(n601) );
  XNOR2_X1 U668 ( .A(n601), .B(KEYINPUT74), .ZN(n603) );
  NOR2_X1 U669 ( .A1(G299), .A2(G868), .ZN(n602) );
  NOR2_X1 U670 ( .A1(n603), .A2(n602), .ZN(G297) );
  NAND2_X1 U671 ( .A1(n604), .A2(G559), .ZN(n605) );
  INV_X1 U672 ( .A(n954), .ZN(n899) );
  NAND2_X1 U673 ( .A1(n605), .A2(n899), .ZN(n606) );
  XNOR2_X1 U674 ( .A(n606), .B(KEYINPUT75), .ZN(n607) );
  XOR2_X1 U675 ( .A(KEYINPUT16), .B(n607), .Z(G148) );
  NOR2_X1 U676 ( .A1(G868), .A2(n950), .ZN(n610) );
  NAND2_X1 U677 ( .A1(n899), .A2(G868), .ZN(n608) );
  NOR2_X1 U678 ( .A1(G559), .A2(n608), .ZN(n609) );
  NOR2_X1 U679 ( .A1(n610), .A2(n609), .ZN(G282) );
  NAND2_X1 U680 ( .A1(G123), .A2(n876), .ZN(n611) );
  XNOR2_X1 U681 ( .A(n611), .B(KEYINPUT18), .ZN(n613) );
  NAND2_X1 U682 ( .A1(n875), .A2(G111), .ZN(n612) );
  NAND2_X1 U683 ( .A1(n613), .A2(n612), .ZN(n617) );
  NAND2_X1 U684 ( .A1(G135), .A2(n879), .ZN(n615) );
  NAND2_X1 U685 ( .A1(G99), .A2(n880), .ZN(n614) );
  NAND2_X1 U686 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U687 ( .A1(n617), .A2(n616), .ZN(n975) );
  XNOR2_X1 U688 ( .A(G2096), .B(n975), .ZN(n619) );
  INV_X1 U689 ( .A(G2100), .ZN(n618) );
  NAND2_X1 U690 ( .A1(n619), .A2(n618), .ZN(G156) );
  NAND2_X1 U691 ( .A1(G67), .A2(n644), .ZN(n621) );
  NAND2_X1 U692 ( .A1(G93), .A2(n645), .ZN(n620) );
  NAND2_X1 U693 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U694 ( .A1(G80), .A2(n648), .ZN(n622) );
  XNOR2_X1 U695 ( .A(KEYINPUT77), .B(n622), .ZN(n623) );
  NOR2_X1 U696 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U697 ( .A1(G55), .A2(n652), .ZN(n625) );
  NAND2_X1 U698 ( .A1(n626), .A2(n625), .ZN(n664) );
  XNOR2_X1 U699 ( .A(n950), .B(KEYINPUT76), .ZN(n628) );
  NAND2_X1 U700 ( .A1(n899), .A2(G559), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n628), .B(n627), .ZN(n661) );
  NOR2_X1 U702 ( .A1(n661), .A2(G860), .ZN(n629) );
  XOR2_X1 U703 ( .A(n664), .B(n629), .Z(G145) );
  NAND2_X1 U704 ( .A1(G651), .A2(G74), .ZN(n631) );
  NAND2_X1 U705 ( .A1(G49), .A2(n652), .ZN(n630) );
  NAND2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U707 ( .A1(n644), .A2(n632), .ZN(n633) );
  XNOR2_X1 U708 ( .A(n633), .B(KEYINPUT78), .ZN(n636) );
  NAND2_X1 U709 ( .A1(G87), .A2(n634), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n636), .A2(n635), .ZN(G288) );
  NAND2_X1 U711 ( .A1(G62), .A2(n644), .ZN(n638) );
  NAND2_X1 U712 ( .A1(G88), .A2(n645), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n641) );
  NAND2_X1 U714 ( .A1(G75), .A2(n648), .ZN(n639) );
  XNOR2_X1 U715 ( .A(KEYINPUT79), .B(n639), .ZN(n640) );
  NOR2_X1 U716 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U717 ( .A1(G50), .A2(n652), .ZN(n642) );
  NAND2_X1 U718 ( .A1(n643), .A2(n642), .ZN(G303) );
  NAND2_X1 U719 ( .A1(G61), .A2(n644), .ZN(n647) );
  NAND2_X1 U720 ( .A1(G86), .A2(n645), .ZN(n646) );
  NAND2_X1 U721 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U722 ( .A1(n648), .A2(G73), .ZN(n649) );
  XOR2_X1 U723 ( .A(KEYINPUT2), .B(n649), .Z(n650) );
  NOR2_X1 U724 ( .A1(n651), .A2(n650), .ZN(n654) );
  NAND2_X1 U725 ( .A1(G48), .A2(n652), .ZN(n653) );
  NAND2_X1 U726 ( .A1(n654), .A2(n653), .ZN(G305) );
  INV_X1 U727 ( .A(G299), .ZN(n951) );
  XNOR2_X1 U728 ( .A(n951), .B(G288), .ZN(n655) );
  XNOR2_X1 U729 ( .A(n655), .B(n664), .ZN(n656) );
  XNOR2_X1 U730 ( .A(KEYINPUT80), .B(n656), .ZN(n658) );
  XNOR2_X1 U731 ( .A(G290), .B(KEYINPUT19), .ZN(n657) );
  XNOR2_X1 U732 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U733 ( .A(n659), .B(G303), .ZN(n660) );
  XNOR2_X1 U734 ( .A(n660), .B(G305), .ZN(n896) );
  XNOR2_X1 U735 ( .A(n661), .B(n896), .ZN(n662) );
  NAND2_X1 U736 ( .A1(n662), .A2(G868), .ZN(n666) );
  NAND2_X1 U737 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U738 ( .A1(n666), .A2(n665), .ZN(G295) );
  NAND2_X1 U739 ( .A1(G2078), .A2(G2084), .ZN(n667) );
  XOR2_X1 U740 ( .A(KEYINPUT20), .B(n667), .Z(n668) );
  NAND2_X1 U741 ( .A1(G2090), .A2(n668), .ZN(n669) );
  XNOR2_X1 U742 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U743 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U744 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U745 ( .A1(G220), .A2(G219), .ZN(n671) );
  XOR2_X1 U746 ( .A(KEYINPUT22), .B(n671), .Z(n672) );
  NOR2_X1 U747 ( .A1(G218), .A2(n672), .ZN(n673) );
  NAND2_X1 U748 ( .A1(G96), .A2(n673), .ZN(n829) );
  NAND2_X1 U749 ( .A1(n829), .A2(G2106), .ZN(n677) );
  NAND2_X1 U750 ( .A1(G120), .A2(G108), .ZN(n674) );
  NOR2_X1 U751 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U752 ( .A1(G69), .A2(n675), .ZN(n830) );
  NAND2_X1 U753 ( .A1(n830), .A2(G567), .ZN(n676) );
  NAND2_X1 U754 ( .A1(n677), .A2(n676), .ZN(n831) );
  NAND2_X1 U755 ( .A1(G483), .A2(G661), .ZN(n678) );
  NOR2_X1 U756 ( .A1(n831), .A2(n678), .ZN(n828) );
  NAND2_X1 U757 ( .A1(n828), .A2(G36), .ZN(G176) );
  INV_X1 U758 ( .A(G303), .ZN(G166) );
  NOR2_X1 U759 ( .A1(n679), .A2(G1384), .ZN(n731) );
  NAND2_X1 U760 ( .A1(G160), .A2(G40), .ZN(n730) );
  NOR2_X1 U761 ( .A1(n731), .A2(n730), .ZN(n726) );
  NAND2_X1 U762 ( .A1(G140), .A2(n879), .ZN(n681) );
  NAND2_X1 U763 ( .A1(G104), .A2(n880), .ZN(n680) );
  NAND2_X1 U764 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U765 ( .A(KEYINPUT34), .B(n682), .ZN(n688) );
  NAND2_X1 U766 ( .A1(G116), .A2(n875), .ZN(n684) );
  NAND2_X1 U767 ( .A1(G128), .A2(n876), .ZN(n683) );
  NAND2_X1 U768 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U769 ( .A(KEYINPUT35), .B(n685), .Z(n686) );
  XNOR2_X1 U770 ( .A(KEYINPUT82), .B(n686), .ZN(n687) );
  NOR2_X1 U771 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U772 ( .A(KEYINPUT36), .B(n689), .ZN(n889) );
  XNOR2_X1 U773 ( .A(G2067), .B(KEYINPUT37), .ZN(n719) );
  NOR2_X1 U774 ( .A1(n889), .A2(n719), .ZN(n974) );
  NAND2_X1 U775 ( .A1(n974), .A2(n726), .ZN(n690) );
  XOR2_X1 U776 ( .A(KEYINPUT83), .B(n690), .Z(n723) );
  NAND2_X1 U777 ( .A1(n875), .A2(G117), .ZN(n697) );
  NAND2_X1 U778 ( .A1(G141), .A2(n879), .ZN(n692) );
  NAND2_X1 U779 ( .A1(G129), .A2(n876), .ZN(n691) );
  NAND2_X1 U780 ( .A1(n692), .A2(n691), .ZN(n695) );
  NAND2_X1 U781 ( .A1(n880), .A2(G105), .ZN(n693) );
  XOR2_X1 U782 ( .A(KEYINPUT38), .B(n693), .Z(n694) );
  NOR2_X1 U783 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U784 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U785 ( .A(KEYINPUT85), .B(n698), .Z(n892) );
  NOR2_X1 U786 ( .A1(G1996), .A2(n892), .ZN(n985) );
  NAND2_X1 U787 ( .A1(G1996), .A2(n892), .ZN(n699) );
  XNOR2_X1 U788 ( .A(n699), .B(KEYINPUT86), .ZN(n708) );
  NAND2_X1 U789 ( .A1(G131), .A2(n879), .ZN(n701) );
  NAND2_X1 U790 ( .A1(G119), .A2(n876), .ZN(n700) );
  NAND2_X1 U791 ( .A1(n701), .A2(n700), .ZN(n705) );
  NAND2_X1 U792 ( .A1(G107), .A2(n875), .ZN(n703) );
  NAND2_X1 U793 ( .A1(G95), .A2(n880), .ZN(n702) );
  NAND2_X1 U794 ( .A1(n703), .A2(n702), .ZN(n704) );
  OR2_X1 U795 ( .A1(n705), .A2(n704), .ZN(n865) );
  NAND2_X1 U796 ( .A1(G1991), .A2(n865), .ZN(n706) );
  XNOR2_X1 U797 ( .A(KEYINPUT84), .B(n706), .ZN(n707) );
  NAND2_X1 U798 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U799 ( .A(n709), .B(KEYINPUT87), .ZN(n971) );
  INV_X1 U800 ( .A(n971), .ZN(n710) );
  NAND2_X1 U801 ( .A1(n710), .A2(n726), .ZN(n724) );
  INV_X1 U802 ( .A(n724), .ZN(n713) );
  NOR2_X1 U803 ( .A1(G1986), .A2(G290), .ZN(n711) );
  NOR2_X1 U804 ( .A1(G1991), .A2(n865), .ZN(n976) );
  NOR2_X1 U805 ( .A1(n711), .A2(n976), .ZN(n712) );
  NOR2_X1 U806 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U807 ( .A1(n985), .A2(n714), .ZN(n715) );
  XOR2_X1 U808 ( .A(n715), .B(KEYINPUT99), .Z(n716) );
  XNOR2_X1 U809 ( .A(KEYINPUT39), .B(n716), .ZN(n717) );
  NAND2_X1 U810 ( .A1(n723), .A2(n717), .ZN(n718) );
  XNOR2_X1 U811 ( .A(n718), .B(KEYINPUT100), .ZN(n720) );
  NAND2_X1 U812 ( .A1(n889), .A2(n719), .ZN(n989) );
  NAND2_X1 U813 ( .A1(n720), .A2(n989), .ZN(n721) );
  NAND2_X1 U814 ( .A1(n726), .A2(n721), .ZN(n722) );
  XNOR2_X1 U815 ( .A(n722), .B(KEYINPUT101), .ZN(n821) );
  NAND2_X1 U816 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U817 ( .A(KEYINPUT88), .B(n725), .Z(n728) );
  XNOR2_X1 U818 ( .A(G1986), .B(G290), .ZN(n949) );
  NAND2_X1 U819 ( .A1(n726), .A2(n949), .ZN(n727) );
  NAND2_X1 U820 ( .A1(n728), .A2(n727), .ZN(n819) );
  XNOR2_X1 U821 ( .A(G1981), .B(KEYINPUT97), .ZN(n729) );
  XNOR2_X1 U822 ( .A(n729), .B(G305), .ZN(n959) );
  INV_X1 U823 ( .A(n730), .ZN(n732) );
  NAND2_X1 U824 ( .A1(n732), .A2(n731), .ZN(n774) );
  NAND2_X1 U825 ( .A1(n774), .A2(G8), .ZN(n733) );
  XOR2_X2 U826 ( .A(KEYINPUT89), .B(n733), .Z(n813) );
  INV_X1 U827 ( .A(n813), .ZN(n807) );
  NOR2_X1 U828 ( .A1(G288), .A2(G1976), .ZN(n734) );
  XOR2_X1 U829 ( .A(n734), .B(KEYINPUT95), .Z(n798) );
  AND2_X1 U830 ( .A1(n807), .A2(n798), .ZN(n735) );
  NAND2_X1 U831 ( .A1(KEYINPUT33), .A2(n735), .ZN(n736) );
  NAND2_X1 U832 ( .A1(n959), .A2(n736), .ZN(n804) );
  NOR2_X1 U833 ( .A1(G1966), .A2(n813), .ZN(n792) );
  NOR2_X1 U834 ( .A1(G2084), .A2(n774), .ZN(n788) );
  NOR2_X1 U835 ( .A1(n792), .A2(n788), .ZN(n737) );
  NAND2_X1 U836 ( .A1(n737), .A2(G8), .ZN(n740) );
  XNOR2_X1 U837 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n738) );
  XNOR2_X1 U838 ( .A(n738), .B(KEYINPUT30), .ZN(n739) );
  NOR2_X1 U839 ( .A1(G168), .A2(n523), .ZN(n744) );
  OR2_X1 U840 ( .A1(n757), .A2(G1961), .ZN(n742) );
  XNOR2_X1 U841 ( .A(G2078), .B(KEYINPUT25), .ZN(n930) );
  NAND2_X1 U842 ( .A1(n757), .A2(n930), .ZN(n741) );
  NAND2_X1 U843 ( .A1(n742), .A2(n741), .ZN(n746) );
  NOR2_X1 U844 ( .A1(G171), .A2(n746), .ZN(n743) );
  NOR2_X1 U845 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U846 ( .A(KEYINPUT31), .B(n745), .Z(n789) );
  NAND2_X1 U847 ( .A1(n746), .A2(G171), .ZN(n772) );
  INV_X1 U848 ( .A(KEYINPUT29), .ZN(n770) );
  NAND2_X1 U849 ( .A1(G2072), .A2(n757), .ZN(n747) );
  XNOR2_X1 U850 ( .A(n747), .B(KEYINPUT90), .ZN(n748) );
  XNOR2_X1 U851 ( .A(KEYINPUT27), .B(n748), .ZN(n750) );
  AND2_X1 U852 ( .A1(n774), .A2(G1956), .ZN(n749) );
  NOR2_X1 U853 ( .A1(n750), .A2(n749), .ZN(n752) );
  OR2_X1 U854 ( .A1(n752), .A2(n951), .ZN(n751) );
  XNOR2_X1 U855 ( .A(n751), .B(KEYINPUT28), .ZN(n768) );
  NAND2_X1 U856 ( .A1(n752), .A2(n951), .ZN(n766) );
  INV_X1 U857 ( .A(G1996), .ZN(n924) );
  NOR2_X1 U858 ( .A1(n774), .A2(n924), .ZN(n753) );
  XOR2_X1 U859 ( .A(n753), .B(KEYINPUT26), .Z(n755) );
  NAND2_X1 U860 ( .A1(n774), .A2(G1341), .ZN(n754) );
  NAND2_X1 U861 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U862 ( .A1(n950), .A2(n756), .ZN(n762) );
  NAND2_X1 U863 ( .A1(n899), .A2(n762), .ZN(n761) );
  NAND2_X1 U864 ( .A1(G1348), .A2(n774), .ZN(n759) );
  NAND2_X1 U865 ( .A1(n757), .A2(G2067), .ZN(n758) );
  NAND2_X1 U866 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U867 ( .A1(n761), .A2(n760), .ZN(n764) );
  OR2_X1 U868 ( .A1(n762), .A2(n899), .ZN(n763) );
  NAND2_X1 U869 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U870 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U871 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U872 ( .A(n770), .B(n769), .ZN(n771) );
  NAND2_X1 U873 ( .A1(n772), .A2(n771), .ZN(n790) );
  INV_X1 U874 ( .A(G8), .ZN(n780) );
  NOR2_X1 U875 ( .A1(G1971), .A2(n813), .ZN(n773) );
  XNOR2_X1 U876 ( .A(KEYINPUT93), .B(n773), .ZN(n778) );
  NOR2_X1 U877 ( .A1(G2090), .A2(n774), .ZN(n775) );
  XNOR2_X1 U878 ( .A(KEYINPUT94), .B(n775), .ZN(n776) );
  NOR2_X1 U879 ( .A1(G166), .A2(n776), .ZN(n777) );
  NAND2_X1 U880 ( .A1(n778), .A2(n777), .ZN(n779) );
  OR2_X1 U881 ( .A1(n780), .A2(n779), .ZN(n782) );
  AND2_X1 U882 ( .A1(n790), .A2(n782), .ZN(n781) );
  NAND2_X1 U883 ( .A1(n789), .A2(n781), .ZN(n786) );
  INV_X1 U884 ( .A(n782), .ZN(n784) );
  AND2_X1 U885 ( .A1(G286), .A2(G8), .ZN(n783) );
  OR2_X1 U886 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U887 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U888 ( .A(n787), .B(KEYINPUT32), .ZN(n796) );
  NAND2_X1 U889 ( .A1(G8), .A2(n788), .ZN(n794) );
  AND2_X1 U890 ( .A1(n790), .A2(n789), .ZN(n791) );
  NOR2_X1 U891 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U892 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U893 ( .A1(n796), .A2(n795), .ZN(n811) );
  NOR2_X1 U894 ( .A1(G1971), .A2(G303), .ZN(n797) );
  NOR2_X1 U895 ( .A1(n798), .A2(n797), .ZN(n965) );
  XNOR2_X1 U896 ( .A(KEYINPUT96), .B(n965), .ZN(n799) );
  NAND2_X1 U897 ( .A1(n811), .A2(n799), .ZN(n801) );
  NAND2_X1 U898 ( .A1(G1976), .A2(G288), .ZN(n946) );
  INV_X1 U899 ( .A(n946), .ZN(n800) );
  AND2_X1 U900 ( .A1(n801), .A2(n522), .ZN(n802) );
  NOR2_X1 U901 ( .A1(KEYINPUT33), .A2(n802), .ZN(n803) );
  NOR2_X1 U902 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U903 ( .A(n805), .B(KEYINPUT98), .ZN(n817) );
  NOR2_X1 U904 ( .A1(G1981), .A2(G305), .ZN(n806) );
  XNOR2_X1 U905 ( .A(KEYINPUT24), .B(n806), .ZN(n808) );
  NAND2_X1 U906 ( .A1(n808), .A2(n807), .ZN(n815) );
  NOR2_X1 U907 ( .A1(G2090), .A2(G303), .ZN(n809) );
  NAND2_X1 U908 ( .A1(G8), .A2(n809), .ZN(n810) );
  NAND2_X1 U909 ( .A1(n811), .A2(n810), .ZN(n812) );
  NAND2_X1 U910 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U911 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U912 ( .A1(n817), .A2(n816), .ZN(n818) );
  NOR2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n822) );
  XOR2_X1 U915 ( .A(KEYINPUT40), .B(n822), .Z(G329) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n823), .ZN(G217) );
  NAND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n825) );
  INV_X1 U918 ( .A(G661), .ZN(n824) );
  NOR2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U920 ( .A(n826), .B(KEYINPUT105), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n828), .A2(n827), .ZN(G188) );
  XNOR2_X1 U923 ( .A(G108), .B(KEYINPUT115), .ZN(G238) );
  INV_X1 U925 ( .A(G120), .ZN(G236) );
  INV_X1 U926 ( .A(G96), .ZN(G221) );
  NOR2_X1 U927 ( .A1(n830), .A2(n829), .ZN(G325) );
  INV_X1 U928 ( .A(G325), .ZN(G261) );
  INV_X1 U929 ( .A(n831), .ZN(G319) );
  XOR2_X1 U930 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n833) );
  XNOR2_X1 U931 ( .A(G2678), .B(G2096), .ZN(n832) );
  XNOR2_X1 U932 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U933 ( .A(n834), .B(KEYINPUT43), .Z(n836) );
  XNOR2_X1 U934 ( .A(G2072), .B(G2090), .ZN(n835) );
  XNOR2_X1 U935 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U936 ( .A(G2100), .B(G2084), .Z(n838) );
  XNOR2_X1 U937 ( .A(G2078), .B(G2067), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U939 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U940 ( .A(KEYINPUT107), .B(KEYINPUT106), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(G227) );
  XOR2_X1 U942 ( .A(G1981), .B(G1971), .Z(n844) );
  XNOR2_X1 U943 ( .A(G1966), .B(G1961), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U945 ( .A(G1991), .B(G1986), .Z(n846) );
  XNOR2_X1 U946 ( .A(G1996), .B(G1976), .ZN(n845) );
  XNOR2_X1 U947 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U948 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U949 ( .A(G2474), .B(KEYINPUT109), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(n851) );
  XNOR2_X1 U951 ( .A(KEYINPUT41), .B(n851), .ZN(n852) );
  XOR2_X1 U952 ( .A(n852), .B(G1956), .Z(G229) );
  NAND2_X1 U953 ( .A1(n880), .A2(G100), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n853), .B(KEYINPUT110), .ZN(n855) );
  NAND2_X1 U955 ( .A1(G112), .A2(n875), .ZN(n854) );
  NAND2_X1 U956 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n856), .B(KEYINPUT111), .ZN(n858) );
  NAND2_X1 U958 ( .A1(G136), .A2(n879), .ZN(n857) );
  NAND2_X1 U959 ( .A1(n858), .A2(n857), .ZN(n861) );
  NAND2_X1 U960 ( .A1(n876), .A2(G124), .ZN(n859) );
  XOR2_X1 U961 ( .A(KEYINPUT44), .B(n859), .Z(n860) );
  NOR2_X1 U962 ( .A1(n861), .A2(n860), .ZN(G162) );
  XOR2_X1 U963 ( .A(KEYINPUT48), .B(KEYINPUT113), .Z(n863) );
  XNOR2_X1 U964 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n862) );
  XNOR2_X1 U965 ( .A(n863), .B(n862), .ZN(n867) );
  XOR2_X1 U966 ( .A(G164), .B(G162), .Z(n864) );
  XNOR2_X1 U967 ( .A(n865), .B(n864), .ZN(n866) );
  XNOR2_X1 U968 ( .A(n867), .B(n866), .ZN(n891) );
  NAND2_X1 U969 ( .A1(G139), .A2(n879), .ZN(n869) );
  NAND2_X1 U970 ( .A1(G103), .A2(n880), .ZN(n868) );
  NAND2_X1 U971 ( .A1(n869), .A2(n868), .ZN(n874) );
  NAND2_X1 U972 ( .A1(G115), .A2(n875), .ZN(n871) );
  NAND2_X1 U973 ( .A1(G127), .A2(n876), .ZN(n870) );
  NAND2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U975 ( .A(KEYINPUT47), .B(n872), .Z(n873) );
  NOR2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n980) );
  XNOR2_X1 U977 ( .A(n980), .B(n975), .ZN(n887) );
  NAND2_X1 U978 ( .A1(G118), .A2(n875), .ZN(n878) );
  NAND2_X1 U979 ( .A1(G130), .A2(n876), .ZN(n877) );
  NAND2_X1 U980 ( .A1(n878), .A2(n877), .ZN(n885) );
  NAND2_X1 U981 ( .A1(G142), .A2(n879), .ZN(n882) );
  NAND2_X1 U982 ( .A1(G106), .A2(n880), .ZN(n881) );
  NAND2_X1 U983 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U984 ( .A(KEYINPUT45), .B(n883), .Z(n884) );
  NOR2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U986 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U987 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U988 ( .A(n891), .B(n890), .ZN(n894) );
  XOR2_X1 U989 ( .A(n892), .B(G160), .Z(n893) );
  XNOR2_X1 U990 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U991 ( .A1(G37), .A2(n895), .ZN(G395) );
  XNOR2_X1 U992 ( .A(n896), .B(KEYINPUT114), .ZN(n898) );
  XNOR2_X1 U993 ( .A(n950), .B(G286), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n898), .B(n897), .ZN(n901) );
  XOR2_X1 U995 ( .A(n899), .B(G171), .Z(n900) );
  XNOR2_X1 U996 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U997 ( .A1(G37), .A2(n902), .ZN(G397) );
  XOR2_X1 U998 ( .A(KEYINPUT102), .B(G2446), .Z(n904) );
  XNOR2_X1 U999 ( .A(G2454), .B(G2451), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n904), .B(n903), .ZN(n908) );
  XOR2_X1 U1001 ( .A(KEYINPUT104), .B(KEYINPUT103), .Z(n906) );
  XNOR2_X1 U1002 ( .A(G2438), .B(G2435), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1004 ( .A(n908), .B(n907), .Z(n910) );
  XNOR2_X1 U1005 ( .A(G2443), .B(G2427), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n910), .B(n909), .ZN(n913) );
  XOR2_X1 U1007 ( .A(G1348), .B(G1341), .Z(n911) );
  XNOR2_X1 U1008 ( .A(G2430), .B(n911), .ZN(n912) );
  XOR2_X1 U1009 ( .A(n913), .B(n912), .Z(n914) );
  NAND2_X1 U1010 ( .A1(G14), .A2(n914), .ZN(n920) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n920), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(G227), .A2(G229), .ZN(n915) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(n915), .ZN(n916) );
  NOR2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(n919) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(G69), .ZN(G235) );
  INV_X1 U1019 ( .A(n920), .ZN(G401) );
  XNOR2_X1 U1020 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n994) );
  XNOR2_X1 U1021 ( .A(G2072), .B(G33), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(G1991), .B(G25), .ZN(n921) );
  NOR2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n929) );
  XOR2_X1 U1024 ( .A(G2067), .B(G26), .Z(n923) );
  NAND2_X1 U1025 ( .A1(n923), .A2(G28), .ZN(n927) );
  XOR2_X1 U1026 ( .A(G32), .B(n924), .Z(n925) );
  XNOR2_X1 U1027 ( .A(KEYINPUT120), .B(n925), .ZN(n926) );
  NOR2_X1 U1028 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n932) );
  XOR2_X1 U1030 ( .A(G27), .B(n930), .Z(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1032 ( .A(KEYINPUT121), .B(n933), .ZN(n934) );
  XNOR2_X1 U1033 ( .A(n934), .B(KEYINPUT53), .ZN(n940) );
  XNOR2_X1 U1034 ( .A(KEYINPUT54), .B(G34), .ZN(n935) );
  XNOR2_X1 U1035 ( .A(n935), .B(KEYINPUT122), .ZN(n936) );
  XNOR2_X1 U1036 ( .A(G2084), .B(n936), .ZN(n938) );
  XNOR2_X1 U1037 ( .A(G2090), .B(G35), .ZN(n937) );
  NOR2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1040 ( .A(n994), .B(n941), .ZN(n943) );
  INV_X1 U1041 ( .A(G29), .ZN(n942) );
  NAND2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1043 ( .A1(n944), .A2(G11), .ZN(n945) );
  XNOR2_X1 U1044 ( .A(KEYINPUT123), .B(n945), .ZN(n1002) );
  XOR2_X1 U1045 ( .A(G16), .B(KEYINPUT56), .Z(n970) );
  XNOR2_X1 U1046 ( .A(G171), .B(G1961), .ZN(n947) );
  NAND2_X1 U1047 ( .A1(n947), .A2(n946), .ZN(n967) );
  AND2_X1 U1048 ( .A1(G303), .A2(G1971), .ZN(n948) );
  NOR2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n958) );
  XOR2_X1 U1050 ( .A(n950), .B(G1341), .Z(n953) );
  XNOR2_X1 U1051 ( .A(n951), .B(G1956), .ZN(n952) );
  NAND2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n956) );
  XNOR2_X1 U1053 ( .A(n954), .B(G1348), .ZN(n955) );
  NOR2_X1 U1054 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(G1966), .B(G168), .ZN(n960) );
  NAND2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1058 ( .A(KEYINPUT57), .B(n961), .Z(n962) );
  NOR2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1062 ( .A(n968), .B(KEYINPUT124), .ZN(n969) );
  NOR2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n1000) );
  XNOR2_X1 U1064 ( .A(G160), .B(G2084), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  NOR2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n978) );
  NOR2_X1 U1067 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1069 ( .A(KEYINPUT116), .B(n979), .ZN(n992) );
  XOR2_X1 U1070 ( .A(G2072), .B(n980), .Z(n982) );
  XOR2_X1 U1071 ( .A(G164), .B(G2078), .Z(n981) );
  NOR2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n983) );
  XOR2_X1 U1073 ( .A(KEYINPUT50), .B(n983), .Z(n988) );
  XOR2_X1 U1074 ( .A(G2090), .B(G162), .Z(n984) );
  NOR2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1076 ( .A(KEYINPUT51), .B(n986), .ZN(n987) );
  NOR2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n990) );
  NAND2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1079 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1080 ( .A(n993), .B(KEYINPUT52), .ZN(n995) );
  NAND2_X1 U1081 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1082 ( .A(KEYINPUT118), .B(n996), .ZN(n997) );
  NAND2_X1 U1083 ( .A1(n997), .A2(G29), .ZN(n998) );
  XNOR2_X1 U1084 ( .A(KEYINPUT119), .B(n998), .ZN(n999) );
  NOR2_X1 U1085 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1086 ( .A1(n1002), .A2(n1001), .ZN(n1028) );
  XNOR2_X1 U1087 ( .A(G1966), .B(G21), .ZN(n1003) );
  XNOR2_X1 U1088 ( .A(n1003), .B(KEYINPUT126), .ZN(n1011) );
  XNOR2_X1 U1089 ( .A(G1971), .B(G22), .ZN(n1005) );
  XNOR2_X1 U1090 ( .A(G1986), .B(G24), .ZN(n1004) );
  NOR2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1008) );
  XNOR2_X1 U1092 ( .A(G1976), .B(KEYINPUT127), .ZN(n1006) );
  XNOR2_X1 U1093 ( .A(n1006), .B(G23), .ZN(n1007) );
  NAND2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(KEYINPUT58), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1096 ( .A1(n1011), .A2(n1010), .ZN(n1022) );
  XOR2_X1 U1097 ( .A(G1341), .B(G19), .Z(n1013) );
  XOR2_X1 U1098 ( .A(G1956), .B(G20), .Z(n1012) );
  NAND2_X1 U1099 ( .A1(n1013), .A2(n1012), .ZN(n1019) );
  XOR2_X1 U1100 ( .A(G1981), .B(G6), .Z(n1017) );
  XOR2_X1 U1101 ( .A(G1348), .B(KEYINPUT125), .Z(n1014) );
  XNOR2_X1 U1102 ( .A(G4), .B(n1014), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(n1015), .B(KEYINPUT59), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1106 ( .A(n1020), .B(KEYINPUT60), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  XNOR2_X1 U1108 ( .A(G5), .B(G1961), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1110 ( .A(KEYINPUT61), .B(n1025), .Z(n1026) );
  NOR2_X1 U1111 ( .A1(G16), .A2(n1026), .ZN(n1027) );
  NOR2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1113 ( .A(n1029), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1114 ( .A(G311), .ZN(G150) );
endmodule

