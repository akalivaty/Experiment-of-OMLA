

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592;

  XOR2_X1 U324 ( .A(n398), .B(n397), .Z(n400) );
  XOR2_X1 U325 ( .A(KEYINPUT36), .B(n486), .Z(n590) );
  INV_X1 U326 ( .A(n585), .ZN(n554) );
  AND2_X1 U327 ( .A1(n574), .A2(n292), .ZN(n480) );
  NOR2_X1 U328 ( .A1(n531), .A2(n523), .ZN(n477) );
  XNOR2_X1 U329 ( .A(n476), .B(n475), .ZN(n531) );
  XOR2_X2 U330 ( .A(n462), .B(n582), .Z(n565) );
  XNOR2_X1 U331 ( .A(n455), .B(n454), .ZN(n582) );
  XOR2_X2 U332 ( .A(n327), .B(n324), .Z(n336) );
  INV_X1 U333 ( .A(KEYINPUT85), .ZN(n320) );
  NOR2_X1 U334 ( .A1(n576), .A2(n335), .ZN(n547) );
  XNOR2_X1 U335 ( .A(n326), .B(n306), .ZN(n307) );
  XNOR2_X1 U336 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U337 ( .A(n563), .B(n562), .ZN(n564) );
  NOR2_X1 U338 ( .A1(n479), .A2(n478), .ZN(n292) );
  AND2_X1 U339 ( .A1(G227GAT), .A2(G233GAT), .ZN(n293) );
  AND2_X1 U340 ( .A1(n565), .A2(n577), .ZN(n463) );
  XNOR2_X1 U341 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n433) );
  AND2_X1 U342 ( .A1(n466), .A2(n559), .ZN(n467) );
  XNOR2_X1 U343 ( .A(n402), .B(n293), .ZN(n315) );
  INV_X1 U344 ( .A(KEYINPUT23), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n315), .B(n449), .ZN(n316) );
  XNOR2_X1 U346 ( .A(n341), .B(KEYINPUT100), .ZN(n367) );
  XNOR2_X1 U347 ( .A(n474), .B(KEYINPUT64), .ZN(n475) );
  XNOR2_X1 U348 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U350 ( .A(n451), .B(n450), .ZN(n452) );
  NOR2_X1 U351 ( .A1(n413), .A2(n590), .ZN(n414) );
  XNOR2_X1 U352 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U353 ( .A(n453), .B(n452), .ZN(n455) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n479) );
  XNOR2_X1 U355 ( .A(KEYINPUT120), .B(n482), .ZN(n570) );
  INV_X1 U356 ( .A(G43GAT), .ZN(n459) );
  XNOR2_X1 U357 ( .A(n483), .B(G190GAT), .ZN(n484) );
  XNOR2_X1 U358 ( .A(n459), .B(KEYINPUT40), .ZN(n460) );
  XNOR2_X1 U359 ( .A(n485), .B(n484), .ZN(G1351GAT) );
  XNOR2_X1 U360 ( .A(n461), .B(n460), .ZN(G1330GAT) );
  XNOR2_X1 U361 ( .A(G106GAT), .B(G78GAT), .ZN(n294) );
  XNOR2_X1 U362 ( .A(n294), .B(G148GAT), .ZN(n451) );
  XOR2_X1 U363 ( .A(G50GAT), .B(G162GAT), .Z(n397) );
  XOR2_X1 U364 ( .A(n451), .B(n397), .Z(n296) );
  NAND2_X1 U365 ( .A1(G228GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U366 ( .A(n296), .B(n295), .ZN(n301) );
  XNOR2_X1 U367 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n297) );
  XNOR2_X1 U368 ( .A(n297), .B(KEYINPUT2), .ZN(n352) );
  XNOR2_X1 U369 ( .A(n352), .B(KEYINPUT24), .ZN(n299) );
  XOR2_X1 U370 ( .A(n302), .B(G204GAT), .Z(n308) );
  XOR2_X1 U371 ( .A(KEYINPUT21), .B(G218GAT), .Z(n304) );
  XNOR2_X1 U372 ( .A(KEYINPUT89), .B(G211GAT), .ZN(n303) );
  XNOR2_X1 U373 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U374 ( .A(G197GAT), .B(n305), .Z(n326) );
  XOR2_X1 U375 ( .A(G22GAT), .B(G155GAT), .Z(n379) );
  XNOR2_X1 U376 ( .A(KEYINPUT22), .B(n379), .ZN(n306) );
  XOR2_X1 U377 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n310) );
  XNOR2_X1 U378 ( .A(G190GAT), .B(KEYINPUT19), .ZN(n309) );
  XNOR2_X1 U379 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U380 ( .A(n311), .B(G183GAT), .Z(n313) );
  XNOR2_X1 U381 ( .A(G169GAT), .B(G176GAT), .ZN(n312) );
  XNOR2_X1 U382 ( .A(n313), .B(n312), .ZN(n327) );
  XOR2_X1 U383 ( .A(G43GAT), .B(G134GAT), .Z(n402) );
  XNOR2_X1 U384 ( .A(G99GAT), .B(G71GAT), .ZN(n314) );
  XNOR2_X1 U385 ( .A(n314), .B(G120GAT), .ZN(n449) );
  XOR2_X1 U386 ( .A(n316), .B(KEYINPUT87), .Z(n319) );
  XNOR2_X1 U387 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n317) );
  XNOR2_X1 U388 ( .A(n317), .B(KEYINPUT84), .ZN(n342) );
  XNOR2_X1 U389 ( .A(KEYINPUT20), .B(n342), .ZN(n318) );
  XNOR2_X1 U390 ( .A(n319), .B(n318), .ZN(n323) );
  XOR2_X1 U391 ( .A(G15GAT), .B(G127GAT), .Z(n380) );
  XNOR2_X1 U392 ( .A(n380), .B(KEYINPUT86), .ZN(n321) );
  NAND2_X1 U393 ( .A1(n479), .A2(n336), .ZN(n325) );
  XNOR2_X1 U394 ( .A(n325), .B(KEYINPUT26), .ZN(n576) );
  XNOR2_X1 U395 ( .A(n327), .B(n326), .ZN(n334) );
  XOR2_X1 U396 ( .A(G92GAT), .B(KEYINPUT97), .Z(n329) );
  NAND2_X1 U397 ( .A1(G226GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U398 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U399 ( .A(G36GAT), .B(KEYINPUT81), .Z(n398) );
  XOR2_X1 U400 ( .A(n330), .B(n398), .Z(n332) );
  XOR2_X1 U401 ( .A(G204GAT), .B(G64GAT), .Z(n437) );
  XNOR2_X1 U402 ( .A(G8GAT), .B(n437), .ZN(n331) );
  XNOR2_X1 U403 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U404 ( .A(n334), .B(n333), .ZN(n523) );
  XOR2_X1 U405 ( .A(n523), .B(KEYINPUT27), .Z(n369) );
  INV_X1 U406 ( .A(n369), .ZN(n335) );
  XNOR2_X1 U407 ( .A(n547), .B(KEYINPUT99), .ZN(n340) );
  NOR2_X1 U408 ( .A1(n336), .A2(n523), .ZN(n337) );
  NOR2_X1 U409 ( .A1(n479), .A2(n337), .ZN(n338) );
  XNOR2_X1 U410 ( .A(KEYINPUT25), .B(n338), .ZN(n339) );
  NAND2_X1 U411 ( .A1(n340), .A2(n339), .ZN(n341) );
  XOR2_X1 U412 ( .A(G85GAT), .B(G162GAT), .Z(n344) );
  XNOR2_X1 U413 ( .A(n342), .B(G134GAT), .ZN(n343) );
  XNOR2_X1 U414 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U415 ( .A(G29GAT), .B(n345), .ZN(n366) );
  XOR2_X1 U416 ( .A(KEYINPUT4), .B(KEYINPUT93), .Z(n347) );
  XNOR2_X1 U417 ( .A(G1GAT), .B(G57GAT), .ZN(n346) );
  XNOR2_X1 U418 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U419 ( .A(G148GAT), .B(G155GAT), .Z(n349) );
  XNOR2_X1 U420 ( .A(G127GAT), .B(G120GAT), .ZN(n348) );
  XNOR2_X1 U421 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U422 ( .A(n351), .B(n350), .ZN(n364) );
  XOR2_X1 U423 ( .A(n352), .B(KEYINPUT1), .Z(n354) );
  NAND2_X1 U424 ( .A1(G225GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U425 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U426 ( .A(KEYINPUT6), .B(KEYINPUT91), .Z(n356) );
  XNOR2_X1 U427 ( .A(KEYINPUT94), .B(KEYINPUT92), .ZN(n355) );
  XNOR2_X1 U428 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U429 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U430 ( .A(KEYINPUT5), .B(KEYINPUT90), .Z(n360) );
  XNOR2_X1 U431 ( .A(KEYINPUT96), .B(KEYINPUT95), .ZN(n359) );
  XNOR2_X1 U432 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U433 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U434 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U435 ( .A(n366), .B(n365), .ZN(n573) );
  NAND2_X1 U436 ( .A1(n367), .A2(n573), .ZN(n374) );
  XNOR2_X1 U437 ( .A(n336), .B(KEYINPUT88), .ZN(n371) );
  XNOR2_X1 U438 ( .A(KEYINPUT28), .B(KEYINPUT67), .ZN(n368) );
  XNOR2_X1 U439 ( .A(n368), .B(n479), .ZN(n528) );
  NAND2_X1 U440 ( .A1(n369), .A2(n528), .ZN(n370) );
  NOR2_X1 U441 ( .A1(n573), .A2(n370), .ZN(n533) );
  NAND2_X1 U442 ( .A1(n371), .A2(n533), .ZN(n372) );
  XNOR2_X1 U443 ( .A(n372), .B(KEYINPUT98), .ZN(n373) );
  NAND2_X1 U444 ( .A1(n374), .A2(n373), .ZN(n489) );
  XOR2_X1 U445 ( .A(KEYINPUT82), .B(G64GAT), .Z(n376) );
  XNOR2_X1 U446 ( .A(G183GAT), .B(G71GAT), .ZN(n375) );
  XNOR2_X1 U447 ( .A(n376), .B(n375), .ZN(n378) );
  XNOR2_X1 U448 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n377) );
  XNOR2_X1 U449 ( .A(n377), .B(KEYINPUT13), .ZN(n448) );
  XOR2_X1 U450 ( .A(n378), .B(n448), .Z(n382) );
  XNOR2_X1 U451 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U452 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U453 ( .A(n383), .B(G78GAT), .Z(n385) );
  XOR2_X1 U454 ( .A(G8GAT), .B(G1GAT), .Z(n418) );
  XNOR2_X1 U455 ( .A(n418), .B(G211GAT), .ZN(n384) );
  XNOR2_X1 U456 ( .A(n385), .B(n384), .ZN(n390) );
  XOR2_X1 U457 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n387) );
  NAND2_X1 U458 ( .A1(G231GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U459 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U460 ( .A(KEYINPUT15), .B(n388), .Z(n389) );
  XNOR2_X1 U461 ( .A(n390), .B(n389), .ZN(n585) );
  NAND2_X1 U462 ( .A1(n489), .A2(n554), .ZN(n413) );
  XOR2_X1 U463 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n392) );
  XNOR2_X1 U464 ( .A(G218GAT), .B(KEYINPUT77), .ZN(n391) );
  XNOR2_X1 U465 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U466 ( .A(KEYINPUT66), .B(G106GAT), .Z(n394) );
  XNOR2_X1 U467 ( .A(G190GAT), .B(G99GAT), .ZN(n393) );
  XNOR2_X1 U468 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U469 ( .A(n396), .B(n395), .Z(n404) );
  NAND2_X1 U470 ( .A1(G232GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U471 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U472 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U473 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U474 ( .A(KEYINPUT9), .B(KEYINPUT80), .Z(n406) );
  XNOR2_X1 U475 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n405) );
  XNOR2_X1 U476 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U477 ( .A(n408), .B(n407), .Z(n412) );
  XNOR2_X1 U478 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n409) );
  XNOR2_X1 U479 ( .A(n409), .B(KEYINPUT7), .ZN(n422) );
  XNOR2_X1 U480 ( .A(G85GAT), .B(KEYINPUT74), .ZN(n410) );
  XOR2_X1 U481 ( .A(n410), .B(G92GAT), .Z(n454) );
  XOR2_X1 U482 ( .A(n422), .B(n454), .Z(n411) );
  XNOR2_X1 U483 ( .A(n412), .B(n411), .ZN(n486) );
  XNOR2_X1 U484 ( .A(n414), .B(KEYINPUT37), .ZN(n521) );
  XOR2_X1 U485 ( .A(G141GAT), .B(G36GAT), .Z(n416) );
  XNOR2_X1 U486 ( .A(G43GAT), .B(G50GAT), .ZN(n415) );
  XNOR2_X1 U487 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U488 ( .A(n418), .B(n417), .Z(n420) );
  NAND2_X1 U489 ( .A1(G229GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U490 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U491 ( .A(n421), .B(KEYINPUT29), .Z(n424) );
  XNOR2_X1 U492 ( .A(n422), .B(KEYINPUT68), .ZN(n423) );
  XNOR2_X1 U493 ( .A(n424), .B(n423), .ZN(n432) );
  XOR2_X1 U494 ( .A(G113GAT), .B(G15GAT), .Z(n426) );
  XNOR2_X1 U495 ( .A(G22GAT), .B(G197GAT), .ZN(n425) );
  XNOR2_X1 U496 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U497 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n428) );
  XNOR2_X1 U498 ( .A(G169GAT), .B(KEYINPUT70), .ZN(n427) );
  XNOR2_X1 U499 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U500 ( .A(n430), .B(n429), .Z(n431) );
  XNOR2_X1 U501 ( .A(n432), .B(n431), .ZN(n548) );
  INV_X1 U502 ( .A(n548), .ZN(n577) );
  INV_X1 U503 ( .A(n433), .ZN(n435) );
  XNOR2_X1 U504 ( .A(G176GAT), .B(KEYINPUT32), .ZN(n434) );
  XNOR2_X1 U505 ( .A(n435), .B(n434), .ZN(n438) );
  INV_X1 U506 ( .A(n438), .ZN(n436) );
  NAND2_X1 U507 ( .A1(n436), .A2(n437), .ZN(n441) );
  INV_X1 U508 ( .A(n437), .ZN(n439) );
  NAND2_X1 U509 ( .A1(n439), .A2(n438), .ZN(n440) );
  NAND2_X1 U510 ( .A1(n441), .A2(n440), .ZN(n443) );
  NAND2_X1 U511 ( .A1(G230GAT), .A2(G233GAT), .ZN(n442) );
  XNOR2_X1 U512 ( .A(n443), .B(n442), .ZN(n447) );
  XOR2_X1 U513 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n445) );
  XNOR2_X1 U514 ( .A(KEYINPUT73), .B(KEYINPUT72), .ZN(n444) );
  XOR2_X1 U515 ( .A(n445), .B(n444), .Z(n446) );
  XNOR2_X1 U516 ( .A(n447), .B(n446), .ZN(n453) );
  XNOR2_X1 U517 ( .A(n449), .B(n448), .ZN(n450) );
  NAND2_X1 U518 ( .A1(n577), .A2(n582), .ZN(n491) );
  NOR2_X1 U519 ( .A1(n521), .A2(n491), .ZN(n457) );
  XNOR2_X1 U520 ( .A(KEYINPUT106), .B(KEYINPUT38), .ZN(n456) );
  XNOR2_X1 U521 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U522 ( .A(KEYINPUT105), .B(n458), .ZN(n506) );
  NOR2_X1 U523 ( .A1(n506), .A2(n336), .ZN(n461) );
  XNOR2_X1 U524 ( .A(KEYINPUT41), .B(KEYINPUT65), .ZN(n462) );
  XNOR2_X1 U525 ( .A(n463), .B(KEYINPUT46), .ZN(n464) );
  NOR2_X1 U526 ( .A1(n585), .A2(n464), .ZN(n465) );
  XNOR2_X1 U527 ( .A(KEYINPUT112), .B(n465), .ZN(n466) );
  INV_X1 U528 ( .A(n486), .ZN(n559) );
  XNOR2_X1 U529 ( .A(n467), .B(KEYINPUT47), .ZN(n473) );
  NOR2_X1 U530 ( .A1(n590), .A2(n554), .ZN(n468) );
  XNOR2_X1 U531 ( .A(n468), .B(KEYINPUT45), .ZN(n469) );
  NAND2_X1 U532 ( .A1(n469), .A2(n582), .ZN(n470) );
  XNOR2_X1 U533 ( .A(n470), .B(KEYINPUT113), .ZN(n471) );
  NAND2_X1 U534 ( .A1(n471), .A2(n548), .ZN(n472) );
  NAND2_X1 U535 ( .A1(n473), .A2(n472), .ZN(n476) );
  INV_X1 U536 ( .A(KEYINPUT48), .ZN(n474) );
  XNOR2_X1 U537 ( .A(KEYINPUT54), .B(n477), .ZN(n574) );
  INV_X1 U538 ( .A(n573), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n480), .B(KEYINPUT55), .ZN(n481) );
  NOR2_X1 U540 ( .A1(n336), .A2(n481), .ZN(n482) );
  NAND2_X1 U541 ( .A1(n486), .A2(n570), .ZN(n485) );
  XOR2_X1 U542 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n483) );
  NOR2_X1 U543 ( .A1(n486), .A2(n554), .ZN(n487) );
  XOR2_X1 U544 ( .A(KEYINPUT16), .B(n487), .Z(n488) );
  XNOR2_X1 U545 ( .A(n488), .B(KEYINPUT83), .ZN(n490) );
  NAND2_X1 U546 ( .A1(n490), .A2(n489), .ZN(n508) );
  NOR2_X1 U547 ( .A1(n508), .A2(n491), .ZN(n492) );
  XNOR2_X1 U548 ( .A(n492), .B(KEYINPUT101), .ZN(n500) );
  NOR2_X1 U549 ( .A1(n573), .A2(n500), .ZN(n494) );
  XNOR2_X1 U550 ( .A(KEYINPUT34), .B(KEYINPUT102), .ZN(n493) );
  XNOR2_X1 U551 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U552 ( .A(G1GAT), .B(n495), .Z(G1324GAT) );
  NOR2_X1 U553 ( .A1(n523), .A2(n500), .ZN(n496) );
  XOR2_X1 U554 ( .A(G8GAT), .B(n496), .Z(G1325GAT) );
  NOR2_X1 U555 ( .A1(n336), .A2(n500), .ZN(n498) );
  XNOR2_X1 U556 ( .A(KEYINPUT35), .B(KEYINPUT103), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U558 ( .A(G15GAT), .B(n499), .Z(G1326GAT) );
  NOR2_X1 U559 ( .A1(n528), .A2(n500), .ZN(n501) );
  XOR2_X1 U560 ( .A(KEYINPUT104), .B(n501), .Z(n502) );
  XNOR2_X1 U561 ( .A(G22GAT), .B(n502), .ZN(G1327GAT) );
  NOR2_X1 U562 ( .A1(n573), .A2(n506), .ZN(n504) );
  XNOR2_X1 U563 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n504), .B(n503), .ZN(G1328GAT) );
  NOR2_X1 U565 ( .A1(n523), .A2(n506), .ZN(n505) );
  XOR2_X1 U566 ( .A(n505), .B(G36GAT), .Z(G1329GAT) );
  NOR2_X1 U567 ( .A1(n528), .A2(n506), .ZN(n507) );
  XOR2_X1 U568 ( .A(G50GAT), .B(n507), .Z(G1331GAT) );
  NAND2_X1 U569 ( .A1(n565), .A2(n548), .ZN(n520) );
  NOR2_X1 U570 ( .A1(n520), .A2(n508), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n509), .B(KEYINPUT107), .ZN(n516) );
  NOR2_X1 U572 ( .A1(n573), .A2(n516), .ZN(n511) );
  XNOR2_X1 U573 ( .A(KEYINPUT42), .B(KEYINPUT108), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U575 ( .A(G57GAT), .B(n512), .Z(G1332GAT) );
  NOR2_X1 U576 ( .A1(n523), .A2(n516), .ZN(n513) );
  XOR2_X1 U577 ( .A(G64GAT), .B(n513), .Z(G1333GAT) );
  NOR2_X1 U578 ( .A1(n336), .A2(n516), .ZN(n515) );
  XNOR2_X1 U579 ( .A(G71GAT), .B(KEYINPUT109), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n515), .B(n514), .ZN(G1334GAT) );
  NOR2_X1 U581 ( .A1(n528), .A2(n516), .ZN(n518) );
  XNOR2_X1 U582 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U584 ( .A(G78GAT), .B(n519), .ZN(G1335GAT) );
  OR2_X1 U585 ( .A1(n521), .A2(n520), .ZN(n527) );
  NOR2_X1 U586 ( .A1(n573), .A2(n527), .ZN(n522) );
  XOR2_X1 U587 ( .A(G85GAT), .B(n522), .Z(G1336GAT) );
  NOR2_X1 U588 ( .A1(n523), .A2(n527), .ZN(n525) );
  XNOR2_X1 U589 ( .A(G92GAT), .B(KEYINPUT111), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(G1337GAT) );
  NOR2_X1 U591 ( .A1(n336), .A2(n527), .ZN(n526) );
  XOR2_X1 U592 ( .A(G99GAT), .B(n526), .Z(G1338GAT) );
  NOR2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U594 ( .A(KEYINPUT44), .B(n529), .Z(n530) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  BUF_X1 U596 ( .A(n531), .Z(n545) );
  NOR2_X1 U597 ( .A1(n336), .A2(n545), .ZN(n532) );
  NAND2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n541) );
  NOR2_X1 U599 ( .A1(n548), .A2(n541), .ZN(n534) );
  XOR2_X1 U600 ( .A(KEYINPUT114), .B(n534), .Z(n535) );
  XNOR2_X1 U601 ( .A(G113GAT), .B(n535), .ZN(G1340GAT) );
  INV_X1 U602 ( .A(n565), .ZN(n550) );
  NOR2_X1 U603 ( .A1(n550), .A2(n541), .ZN(n537) );
  XNOR2_X1 U604 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U606 ( .A(G120GAT), .B(n538), .Z(G1341GAT) );
  NOR2_X1 U607 ( .A1(n554), .A2(n541), .ZN(n539) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(n539), .Z(n540) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  NOR2_X1 U610 ( .A1(n559), .A2(n541), .ZN(n543) );
  XNOR2_X1 U611 ( .A(KEYINPUT116), .B(KEYINPUT51), .ZN(n542) );
  XNOR2_X1 U612 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U613 ( .A(G134GAT), .B(n544), .ZN(G1343GAT) );
  NOR2_X1 U614 ( .A1(n573), .A2(n545), .ZN(n546) );
  NAND2_X1 U615 ( .A1(n547), .A2(n546), .ZN(n558) );
  NOR2_X1 U616 ( .A1(n548), .A2(n558), .ZN(n549) );
  XOR2_X1 U617 ( .A(G141GAT), .B(n549), .Z(G1344GAT) );
  NOR2_X1 U618 ( .A1(n550), .A2(n558), .ZN(n552) );
  XNOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(n553), .ZN(G1345GAT) );
  NOR2_X1 U622 ( .A1(n554), .A2(n558), .ZN(n556) );
  XNOR2_X1 U623 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(G155GAT), .B(n557), .ZN(G1346GAT) );
  NOR2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G162GAT), .B(KEYINPUT119), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n577), .A2(n570), .ZN(n563) );
  XOR2_X1 U630 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n562) );
  XNOR2_X1 U631 ( .A(G169GAT), .B(n564), .ZN(G1348GAT) );
  XOR2_X1 U632 ( .A(G176GAT), .B(KEYINPUT123), .Z(n567) );
  NAND2_X1 U633 ( .A1(n565), .A2(n570), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n569) );
  XOR2_X1 U635 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  NAND2_X1 U637 ( .A1(n570), .A2(n585), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(KEYINPUT124), .ZN(n572) );
  XNOR2_X1 U639 ( .A(G183GAT), .B(n572), .ZN(G1350GAT) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n586) );
  NAND2_X1 U642 ( .A1(n586), .A2(n577), .ZN(n581) );
  XOR2_X1 U643 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n579) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  INV_X1 U648 ( .A(n586), .ZN(n589) );
  OR2_X1 U649 ( .A1(n589), .A2(n582), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  XOR2_X1 U651 ( .A(G211GAT), .B(KEYINPUT127), .Z(n588) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U655 ( .A(KEYINPUT62), .B(n591), .Z(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

