//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n570, new_n571,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n585, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n628, new_n629, new_n632,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1220;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT66), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  NAND2_X1  g033(.A1(G113), .A2(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n466), .A2(G2105), .B1(G101), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n461), .B1(new_n471), .B2(KEYINPUT67), .ZN(new_n472));
  OR3_X1    g047(.A1(new_n462), .A2(KEYINPUT67), .A3(G2104), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n472), .A2(G137), .A3(new_n467), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G112), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G2105), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n472), .A2(G2105), .A3(new_n473), .ZN(new_n480));
  INV_X1    g055(.A(G124), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT69), .Z(new_n483));
  NAND3_X1  g058(.A1(new_n472), .A2(new_n467), .A3(new_n473), .ZN(new_n484));
  OR2_X1    g059(.A1(new_n484), .A2(KEYINPUT68), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n484), .A2(KEYINPUT68), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI211_X1 g062(.A(new_n479), .B(new_n483), .C1(G136), .C2(new_n487), .ZN(G162));
  NAND2_X1  g063(.A1(new_n467), .A2(G138), .ZN(new_n489));
  NOR3_X1   g064(.A1(new_n464), .A2(KEYINPUT4), .A3(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n472), .A2(G138), .A3(new_n467), .A4(new_n473), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(G126), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n467), .A2(G114), .ZN(new_n495));
  OAI22_X1  g070(.A1(new_n480), .A2(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n492), .A2(new_n496), .ZN(G164));
  INV_X1    g072(.A(G651), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT6), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G651), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT71), .ZN(new_n503));
  OAI21_X1  g078(.A(G543), .B1(new_n503), .B2(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n503), .A2(KEYINPUT70), .A3(KEYINPUT5), .A4(G543), .ZN(new_n507));
  AOI211_X1 g082(.A(KEYINPUT72), .B(new_n502), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n510), .B1(KEYINPUT71), .B2(new_n511), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n507), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n499), .A2(new_n501), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n509), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n508), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n502), .A2(new_n510), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n517), .A2(G88), .B1(G50), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT73), .ZN(new_n520));
  INV_X1    g095(.A(new_n514), .ZN(new_n521));
  INV_X1    g096(.A(G62), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n514), .A2(KEYINPUT73), .A3(G62), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n519), .A2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  INV_X1    g104(.A(G89), .ZN(new_n530));
  NOR3_X1   g105(.A1(new_n508), .A2(new_n516), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n498), .B1(new_n506), .B2(new_n507), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G63), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n499), .A2(new_n501), .A3(G51), .A4(G543), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n533), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n531), .A2(new_n537), .ZN(G168));
  NAND2_X1  g113(.A1(new_n518), .A2(G52), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n540), .B2(new_n498), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n541), .B1(G90), .B2(new_n517), .ZN(G171));
  INV_X1    g117(.A(KEYINPUT76), .ZN(new_n543));
  INV_X1    g118(.A(new_n518), .ZN(new_n544));
  XOR2_X1   g119(.A(KEYINPUT75), .B(G43), .Z(new_n545));
  NOR2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n546), .B1(new_n517), .B2(G81), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n548), .B1(new_n506), .B2(new_n507), .ZN(new_n549));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  OAI21_X1  g126(.A(KEYINPUT74), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n511), .A2(KEYINPUT71), .ZN(new_n553));
  AOI21_X1  g128(.A(new_n513), .B1(new_n553), .B2(G543), .ZN(new_n554));
  INV_X1    g129(.A(new_n507), .ZN(new_n555));
  OAI21_X1  g130(.A(G56), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT74), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n556), .A2(new_n557), .A3(new_n550), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n552), .A2(new_n558), .A3(G651), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n543), .B1(new_n547), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n515), .B1(new_n554), .B2(new_n555), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT72), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n514), .A2(new_n509), .A3(new_n515), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n562), .A2(G81), .A3(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n546), .ZN(new_n565));
  AND4_X1   g140(.A1(new_n543), .A2(new_n559), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n560), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G860), .ZN(G153));
  AND3_X1   g144(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G36), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT77), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n570), .A2(new_n574), .ZN(G188));
  AOI22_X1  g150(.A1(new_n514), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n576), .A2(new_n498), .ZN(new_n577));
  INV_X1    g152(.A(G53), .ZN(new_n578));
  OAI21_X1  g153(.A(KEYINPUT9), .B1(new_n544), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT9), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n518), .A2(new_n580), .A3(G53), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n562), .A2(G91), .A3(new_n563), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n577), .A2(new_n582), .A3(new_n583), .ZN(G299));
  NAND3_X1  g159(.A1(new_n562), .A2(G90), .A3(new_n563), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n585), .B(new_n539), .C1(new_n498), .C2(new_n540), .ZN(G301));
  INV_X1    g161(.A(G168), .ZN(G286));
  NAND2_X1  g162(.A1(new_n517), .A2(G87), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n518), .A2(G49), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G288));
  AOI22_X1  g166(.A1(new_n514), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n592), .A2(new_n498), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n518), .A2(G48), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n562), .A2(new_n563), .ZN(new_n596));
  INV_X1    g171(.A(G86), .ZN(new_n597));
  OAI21_X1  g172(.A(KEYINPUT78), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n517), .A2(new_n599), .A3(G86), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n595), .B1(new_n598), .B2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G305));
  NAND2_X1  g177(.A1(new_n518), .A2(G47), .ZN(new_n603));
  INV_X1    g178(.A(G85), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n596), .B2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT79), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n605), .A2(new_n606), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n609));
  OAI22_X1  g184(.A1(new_n607), .A2(new_n608), .B1(new_n498), .B2(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n562), .A2(G92), .A3(new_n563), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(KEYINPUT10), .ZN(new_n613));
  NAND2_X1  g188(.A1(G79), .A2(G543), .ZN(new_n614));
  INV_X1    g189(.A(G66), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n521), .B2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n616), .A2(G651), .B1(G54), .B2(new_n518), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT10), .ZN(new_n618));
  NAND4_X1  g193(.A1(new_n562), .A2(new_n618), .A3(G92), .A4(new_n563), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n613), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n621));
  OR2_X1    g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n611), .B1(new_n625), .B2(G868), .ZN(G321));
  XOR2_X1   g201(.A(G321), .B(KEYINPUT81), .Z(G284));
  NAND2_X1  g202(.A1(G286), .A2(G868), .ZN(new_n628));
  AND3_X1   g203(.A1(new_n577), .A2(new_n582), .A3(new_n583), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n628), .B1(G868), .B2(new_n629), .ZN(G297));
  OAI21_X1  g205(.A(new_n628), .B1(G868), .B2(new_n629), .ZN(G280));
  INV_X1    g206(.A(G559), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n625), .B1(new_n632), .B2(G860), .ZN(G148));
  NAND2_X1  g208(.A1(new_n625), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G868), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(G868), .B2(new_n568), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g212(.A(G123), .ZN(new_n638));
  NOR2_X1   g213(.A1(new_n480), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT82), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n487), .A2(G135), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n467), .A2(G111), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n640), .B(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  NAND3_X1  g220(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT12), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT13), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2100), .Z(new_n649));
  NAND2_X1  g224(.A1(new_n645), .A2(new_n649), .ZN(G156));
  XOR2_X1   g225(.A(KEYINPUT83), .B(G2438), .Z(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT15), .B(G2435), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2427), .B(G2430), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT84), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT14), .ZN(new_n657));
  AND2_X1   g232(.A1(new_n657), .A2(KEYINPUT85), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(KEYINPUT85), .ZN(new_n659));
  OAI22_X1  g234(.A1(new_n658), .A2(new_n659), .B1(new_n655), .B2(new_n653), .ZN(new_n660));
  XOR2_X1   g235(.A(G2451), .B(G2454), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT16), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n660), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G1341), .B(G1348), .Z(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT86), .ZN(new_n668));
  INV_X1    g243(.A(G14), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n665), .B2(new_n666), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G401));
  XOR2_X1   g247(.A(G2072), .B(G2078), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  XOR2_X1   g250(.A(G2084), .B(G2090), .Z(new_n676));
  NAND3_X1  g251(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT18), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(KEYINPUT87), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(new_n673), .ZN(new_n680));
  INV_X1    g255(.A(new_n676), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n673), .B(KEYINPUT17), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n680), .B(new_n681), .C1(new_n679), .C2(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n682), .A2(new_n679), .A3(new_n676), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n678), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G2096), .B(G2100), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(G227));
  XOR2_X1   g263(.A(G1956), .B(G2474), .Z(new_n689));
  XOR2_X1   g264(.A(G1961), .B(G1966), .Z(new_n690));
  AND2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g266(.A1(new_n691), .A2(KEYINPUT88), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1971), .B(G1976), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT19), .ZN(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n691), .A2(KEYINPUT88), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n692), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT20), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n689), .A2(new_n690), .ZN(new_n699));
  AOI22_X1  g274(.A1(new_n697), .A2(new_n698), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  OR3_X1    g275(.A1(new_n695), .A2(new_n691), .A3(new_n699), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n700), .B(new_n701), .C1(new_n698), .C2(new_n697), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1991), .B(G1996), .ZN(new_n705));
  INV_X1    g280(.A(G1981), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G1986), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n704), .B(new_n708), .ZN(G229));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G4), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n625), .B2(new_n710), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT97), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1348), .ZN(new_n714));
  INV_X1    g289(.A(G11), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n715), .A2(KEYINPUT31), .ZN(new_n716));
  NOR2_X1   g291(.A1(G29), .A2(G32), .ZN(new_n717));
  NAND3_X1  g292(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT26), .Z(new_n719));
  INV_X1    g294(.A(G105), .ZN(new_n720));
  INV_X1    g295(.A(G129), .ZN(new_n721));
  OAI221_X1 g296(.A(new_n719), .B1(new_n720), .B2(new_n468), .C1(new_n480), .C2(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(new_n487), .B2(G141), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n717), .B1(new_n723), .B2(G29), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT27), .B(G1996), .Z(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G1966), .ZN(new_n727));
  NAND2_X1  g302(.A1(G168), .A2(G16), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G16), .B2(G21), .ZN(new_n729));
  AOI211_X1 g304(.A(new_n716), .B(new_n726), .C1(new_n727), .C2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G27), .ZN(new_n731));
  OAI21_X1  g306(.A(KEYINPUT99), .B1(new_n731), .B2(G29), .ZN(new_n732));
  OR3_X1    g307(.A1(new_n731), .A2(KEYINPUT99), .A3(G29), .ZN(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n732), .B(new_n733), .C1(G164), .C2(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT100), .B(G2078), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  AND2_X1   g312(.A1(KEYINPUT24), .A2(G34), .ZN(new_n738));
  NOR2_X1   g313(.A1(KEYINPUT24), .A2(G34), .ZN(new_n739));
  NOR3_X1   g314(.A1(new_n738), .A2(new_n739), .A3(G29), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n475), .B2(G29), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G2084), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT30), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(G28), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(G28), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n744), .A2(new_n745), .A3(new_n734), .ZN(new_n746));
  AND3_X1   g321(.A1(new_n737), .A2(new_n742), .A3(new_n746), .ZN(new_n747));
  OAI211_X1 g322(.A(new_n730), .B(new_n747), .C1(new_n734), .C2(new_n644), .ZN(new_n748));
  NOR2_X1   g323(.A1(G29), .A2(G33), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n487), .A2(G139), .ZN(new_n751));
  NAND2_X1  g326(.A1(G115), .A2(G2104), .ZN(new_n752));
  INV_X1    g327(.A(G127), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n752), .B1(new_n464), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G2105), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n469), .A2(G103), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT25), .Z(new_n757));
  NAND3_X1  g332(.A1(new_n751), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT98), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n750), .B1(new_n760), .B2(new_n734), .ZN(new_n761));
  INV_X1    g336(.A(G2072), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI211_X1 g338(.A(G2072), .B(new_n750), .C1(new_n760), .C2(new_n734), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n724), .A2(new_n725), .ZN(new_n765));
  NAND2_X1  g340(.A1(G171), .A2(G16), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G5), .B2(G16), .ZN(new_n767));
  INV_X1    g342(.A(G1961), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n763), .A2(new_n764), .A3(new_n765), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n748), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n715), .A2(KEYINPUT31), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n767), .A2(new_n768), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n729), .A2(new_n727), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n771), .A2(new_n772), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT101), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n748), .A2(new_n770), .A3(new_n774), .ZN(new_n779));
  NAND4_X1  g354(.A1(new_n779), .A2(KEYINPUT101), .A3(new_n772), .A4(new_n773), .ZN(new_n780));
  AND2_X1   g355(.A1(KEYINPUT91), .A2(G16), .ZN(new_n781));
  NOR2_X1   g356(.A1(KEYINPUT91), .A2(G16), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n784), .A2(KEYINPUT23), .A3(G20), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT23), .ZN(new_n786));
  INV_X1    g361(.A(G20), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n783), .B2(new_n787), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n785), .B(new_n788), .C1(new_n629), .C2(new_n710), .ZN(new_n789));
  INV_X1    g364(.A(G1956), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n783), .A2(G19), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n568), .B2(new_n783), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(G1341), .Z(new_n794));
  NAND4_X1  g369(.A1(new_n778), .A2(new_n780), .A3(new_n791), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n710), .A2(G6), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n601), .B2(new_n710), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT32), .B(G1981), .Z(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n796), .B(new_n798), .C1(new_n601), .C2(new_n710), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT92), .B(KEYINPUT33), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(G1976), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(G288), .A2(G16), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n710), .A2(G23), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n807), .ZN(new_n809));
  AOI211_X1 g384(.A(new_n804), .B(new_n809), .C1(G288), .C2(G16), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT34), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n784), .A2(G22), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT93), .B(G1971), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n813), .B(new_n814), .C1(G166), .C2(new_n784), .ZN(new_n815));
  INV_X1    g390(.A(new_n814), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n784), .B1(new_n519), .B2(new_n527), .ZN(new_n817));
  INV_X1    g392(.A(new_n813), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n816), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n802), .A2(new_n811), .A3(new_n812), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(G290), .A2(new_n783), .ZN(new_n822));
  INV_X1    g397(.A(G1986), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n784), .A2(G24), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n823), .B1(new_n822), .B2(new_n824), .ZN(new_n826));
  INV_X1    g401(.A(new_n826), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n487), .A2(G131), .ZN(new_n828));
  INV_X1    g403(.A(G119), .ZN(new_n829));
  OAI21_X1  g404(.A(G2104), .B1(new_n467), .B2(G107), .ZN(new_n830));
  NOR2_X1   g405(.A1(G95), .A2(G2105), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT89), .ZN(new_n832));
  OAI22_X1  g407(.A1(new_n480), .A2(new_n829), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n828), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(G29), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n734), .A2(G25), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT35), .B(G1991), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT90), .Z(new_n839));
  AND3_X1   g414(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n839), .B1(new_n836), .B2(new_n837), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n821), .A2(new_n825), .A3(new_n827), .A4(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT94), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n815), .B(new_n819), .C1(new_n808), .C2(new_n810), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n800), .A2(new_n801), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n826), .B1(new_n848), .B2(new_n812), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n849), .A2(KEYINPUT94), .A3(new_n825), .A4(new_n842), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n845), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(KEYINPUT34), .B1(new_n846), .B2(new_n847), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT95), .B(KEYINPUT36), .Z(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT36), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(new_n851), .B2(new_n852), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT96), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n854), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n851), .A2(KEYINPUT96), .A3(new_n852), .A4(new_n853), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n795), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n734), .A2(G35), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n861), .B1(G162), .B2(new_n734), .ZN(new_n862));
  XOR2_X1   g437(.A(KEYINPUT29), .B(G2090), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n734), .A2(G26), .ZN(new_n865));
  INV_X1    g440(.A(G128), .ZN(new_n866));
  OAI21_X1  g441(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n467), .A2(G116), .ZN(new_n868));
  OAI22_X1  g443(.A1(new_n480), .A2(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(new_n487), .B2(G140), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n865), .B1(new_n870), .B2(new_n734), .ZN(new_n871));
  MUX2_X1   g446(.A(new_n865), .B(new_n871), .S(KEYINPUT28), .Z(new_n872));
  INV_X1    g447(.A(G2067), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  AND4_X1   g449(.A1(new_n714), .A2(new_n860), .A3(new_n864), .A4(new_n874), .ZN(G311));
  NAND4_X1  g450(.A1(new_n860), .A2(new_n714), .A3(new_n864), .A4(new_n874), .ZN(G150));
  NAND2_X1  g451(.A1(new_n518), .A2(G55), .ZN(new_n877));
  AOI22_X1  g452(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n877), .B1(new_n878), .B2(new_n498), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n879), .B1(G93), .B2(new_n517), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(G860), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n882), .B(KEYINPUT37), .Z(new_n883));
  NAND2_X1  g458(.A1(new_n625), .A2(G559), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n881), .B1(new_n560), .B2(new_n566), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n559), .A2(new_n564), .A3(new_n565), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n884), .B(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n883), .B1(new_n891), .B2(G860), .ZN(G145));
  XNOR2_X1  g467(.A(new_n758), .B(KEYINPUT98), .ZN(new_n893));
  INV_X1    g468(.A(new_n723), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n760), .A2(new_n723), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n870), .B(G164), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(KEYINPUT103), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT102), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n487), .A2(G142), .ZN(new_n905));
  OR2_X1    g480(.A1(G106), .A2(G2105), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n906), .B(G2104), .C1(G118), .C2(new_n467), .ZN(new_n907));
  INV_X1    g482(.A(G130), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n905), .B(new_n907), .C1(new_n908), .C2(new_n480), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n834), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n834), .A2(new_n909), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n904), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n910), .A2(new_n904), .A3(new_n911), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n913), .A2(new_n647), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n647), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n900), .A2(new_n918), .A3(new_n901), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n903), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT104), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n917), .A2(new_n902), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n644), .B(new_n475), .ZN(new_n923));
  XOR2_X1   g498(.A(new_n923), .B(G162), .Z(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n903), .A2(new_n917), .A3(new_n926), .A4(new_n919), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n921), .A2(new_n922), .A3(new_n925), .A4(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n917), .B(new_n902), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n924), .ZN(new_n930));
  INV_X1    g505(.A(G37), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g508(.A1(new_n881), .A2(G868), .ZN(new_n934));
  XOR2_X1   g509(.A(new_n634), .B(new_n888), .Z(new_n935));
  NAND2_X1  g510(.A1(new_n620), .A2(new_n629), .ZN(new_n936));
  NAND4_X1  g511(.A1(G299), .A2(new_n617), .A3(new_n613), .A4(new_n619), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT41), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n936), .A2(new_n937), .A3(KEYINPUT41), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(G290), .A2(G166), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(G290), .A2(G166), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n601), .A2(G288), .ZN(new_n948));
  INV_X1    g523(.A(G288), .ZN(new_n949));
  NOR2_X1   g524(.A1(G305), .A2(new_n949), .ZN(new_n950));
  OAI22_X1  g525(.A1(new_n946), .A2(new_n947), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n947), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n950), .A2(new_n948), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(new_n945), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n955), .B(KEYINPUT42), .ZN(new_n956));
  OAI221_X1 g531(.A(new_n939), .B1(new_n935), .B2(new_n944), .C1(new_n956), .C2(KEYINPUT105), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(KEYINPUT105), .ZN(new_n958));
  XOR2_X1   g533(.A(new_n957), .B(new_n958), .Z(new_n959));
  AOI21_X1  g534(.A(new_n934), .B1(new_n959), .B2(G868), .ZN(G295));
  AOI21_X1  g535(.A(new_n934), .B1(new_n959), .B2(G868), .ZN(G331));
  NAND3_X1  g536(.A1(new_n562), .A2(G89), .A3(new_n563), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT106), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n535), .A2(new_n536), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n964), .B1(G63), .B2(new_n532), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n963), .B1(new_n962), .B2(new_n965), .ZN(new_n967));
  OAI21_X1  g542(.A(G171), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT106), .B1(new_n531), .B2(new_n537), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n969), .A2(G301), .A3(new_n970), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n885), .A2(new_n887), .A3(new_n968), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n968), .A2(new_n971), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n886), .A2(KEYINPUT76), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n559), .A2(new_n543), .A3(new_n564), .A4(new_n565), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n880), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n887), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n973), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n972), .A2(new_n938), .A3(new_n978), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n972), .A2(new_n978), .B1(new_n941), .B2(new_n942), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT107), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n973), .A2(new_n976), .A3(new_n977), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n885), .A2(new_n887), .B1(new_n968), .B2(new_n971), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n943), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT107), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n981), .A2(new_n955), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT108), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n984), .A2(KEYINPUT109), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n980), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n972), .A2(new_n978), .A3(new_n938), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT110), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n972), .A2(new_n978), .A3(KEYINPUT110), .A4(new_n938), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n989), .A2(new_n991), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n955), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n981), .A2(new_n999), .A3(new_n955), .A4(new_n986), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n988), .A2(new_n998), .A3(new_n931), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT43), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n985), .B1(new_n984), .B2(new_n992), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n972), .A2(new_n978), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT107), .B1(new_n1005), .B2(new_n943), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n997), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n988), .A2(new_n931), .A3(new_n1000), .A4(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n1008), .A2(new_n1002), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n1003), .A2(new_n1009), .A3(KEYINPUT44), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n984), .A2(new_n992), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1006), .B1(new_n1012), .B2(KEYINPUT107), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n999), .B1(new_n1013), .B2(new_n955), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1000), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1016), .A2(KEYINPUT43), .A3(new_n931), .A4(new_n998), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1008), .A2(new_n1002), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1011), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT111), .B1(new_n1010), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1018), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1022));
  OAI21_X1  g597(.A(KEYINPUT44), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT111), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1025), .B(new_n1011), .C1(new_n1002), .C2(new_n1008), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1020), .A2(new_n1027), .ZN(G397));
  INV_X1    g603(.A(G290), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n823), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1030), .B(KEYINPUT113), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n870), .B(G2067), .ZN(new_n1033));
  XNOR2_X1  g608(.A(new_n723), .B(G1996), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n835), .A2(new_n838), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n835), .A2(new_n838), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1035), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1032), .B(new_n1038), .C1(new_n823), .C2(new_n1029), .ZN(new_n1039));
  OR3_X1    g614(.A1(G164), .A2(KEYINPUT112), .A3(G1384), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT45), .ZN(new_n1041));
  OAI21_X1  g616(.A(KEYINPUT112), .B1(G164), .B2(G1384), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n470), .A2(G40), .A3(new_n474), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1039), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n601), .A2(new_n706), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n596), .A2(new_n597), .ZN(new_n1048));
  OAI21_X1  g623(.A(G1981), .B1(new_n595), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT49), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(KEYINPUT115), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(G164), .B2(G1384), .ZN(new_n1054));
  INV_X1    g629(.A(G1384), .ZN(new_n1055));
  OAI211_X1 g630(.A(KEYINPUT114), .B(new_n1055), .C1(new_n492), .C2(new_n496), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1044), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G8), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1051), .A2(KEYINPUT115), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1047), .A2(new_n1049), .A3(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1052), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n949), .A2(G1976), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1059), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT52), .ZN(new_n1065));
  INV_X1    g640(.A(G1976), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT52), .B1(G288), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1059), .A2(new_n1063), .A3(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1062), .A2(new_n1065), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(G164), .A2(G1384), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1044), .B1(new_n1071), .B2(KEYINPUT45), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1041), .B1(G164), .B2(G1384), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1971), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT50), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT50), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1071), .A2(new_n1078), .ZN(new_n1079));
  OR3_X1    g654(.A1(new_n1077), .A2(new_n1044), .A3(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1076), .B1(new_n1080), .B2(G2090), .ZN(new_n1081));
  NAND2_X1  g656(.A1(G303), .A2(G8), .ZN(new_n1082));
  XOR2_X1   g657(.A(new_n1082), .B(KEYINPUT55), .Z(new_n1083));
  NAND3_X1  g658(.A1(new_n1081), .A2(G8), .A3(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1054), .A2(KEYINPUT50), .A3(new_n1056), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1044), .B1(new_n1071), .B2(new_n1078), .ZN(new_n1086));
  INV_X1    g661(.A(G2090), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1058), .B1(new_n1076), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1089), .A2(new_n1083), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1090), .A2(KEYINPUT116), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1089), .A2(new_n1083), .A3(new_n1092), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1070), .B(new_n1084), .C1(new_n1091), .C2(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT123), .B(KEYINPUT53), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1074), .B2(G2078), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1054), .A2(new_n1041), .A3(new_n1056), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n1072), .ZN(new_n1098));
  INV_X1    g673(.A(G2078), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT53), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1077), .A2(new_n1079), .A3(new_n1044), .ZN(new_n1101));
  OAI221_X1 g676(.A(new_n1096), .B1(new_n1098), .B2(new_n1100), .C1(G1961), .C2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n1103));
  AND3_X1   g678(.A1(new_n1102), .A2(new_n1103), .A3(G171), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1103), .B1(new_n1102), .B2(G171), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1094), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1098), .A2(new_n727), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  NOR4_X1   g684(.A1(new_n1077), .A2(new_n1079), .A3(G2084), .A4(new_n1044), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT122), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(G2084), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1101), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT122), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(new_n1114), .A3(new_n1108), .ZN(new_n1115));
  AND3_X1   g690(.A1(new_n1111), .A2(new_n1115), .A3(G168), .ZN(new_n1116));
  NAND2_X1  g691(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1058), .B1(new_n1113), .B2(new_n1108), .ZN(new_n1118));
  OAI22_X1  g693(.A1(new_n1116), .A2(new_n1117), .B1(KEYINPUT51), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1111), .A2(new_n1115), .ZN(new_n1121));
  OAI211_X1 g696(.A(G8), .B(G286), .C1(new_n1121), .C2(new_n1117), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1119), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT126), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1107), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1124), .B1(new_n1107), .B2(new_n1123), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1120), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(G1348), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1080), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1057), .A2(new_n873), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT117), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1057), .A2(KEYINPUT117), .A3(new_n873), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1130), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n624), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n625), .A2(KEYINPUT121), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1136), .A2(KEYINPUT60), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1130), .A2(new_n1135), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT60), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1137), .B(new_n624), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1140), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(G1956), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1147));
  XNOR2_X1  g722(.A(KEYINPUT56), .B(G2072), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g724(.A(G299), .B(KEYINPUT57), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1152), .A2(KEYINPUT120), .A3(new_n1153), .ZN(new_n1154));
  XOR2_X1   g729(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n1155));
  OAI21_X1  g730(.A(new_n1154), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT119), .ZN(new_n1157));
  XOR2_X1   g732(.A(KEYINPUT118), .B(G1996), .Z(new_n1158));
  NOR2_X1   g733(.A1(new_n1074), .A2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(KEYINPUT58), .B(G1341), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1057), .A2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1157), .B(new_n568), .C1(new_n1159), .C2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT59), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1145), .A2(new_n1156), .A3(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1136), .A2(new_n624), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1165), .B1(new_n1166), .B2(new_n1152), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1094), .B1(new_n1164), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1080), .A2(new_n768), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1169), .A2(new_n1096), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1043), .A2(KEYINPUT53), .A3(new_n1099), .A4(new_n1072), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT125), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1170), .A2(G301), .A3(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT54), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1106), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1170), .A2(G171), .A3(new_n1172), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1174), .B1(new_n1102), .B2(G301), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI22_X1  g754(.A1(new_n1176), .A2(new_n1179), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1168), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1062), .A2(new_n1066), .A3(new_n949), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n1047), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(new_n1059), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1118), .A2(G168), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1083), .B1(new_n1081), .B2(G8), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1185), .A2(new_n1186), .A3(new_n1069), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT63), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1184), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1118), .A2(new_n1188), .A3(G168), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1084), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1189), .B1(new_n1070), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1181), .A2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1046), .B1(new_n1128), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1045), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT46), .ZN(new_n1197));
  OR3_X1    g772(.A1(new_n1196), .A2(new_n1197), .A3(G1996), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1033), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1045), .B1(new_n1199), .B2(new_n894), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1197), .B1(new_n1196), .B2(G1996), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1198), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1202), .B(KEYINPUT127), .ZN(new_n1203));
  XNOR2_X1  g778(.A(new_n1203), .B(KEYINPUT47), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n870), .A2(new_n873), .ZN(new_n1205));
  INV_X1    g780(.A(new_n1037), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1205), .B1(new_n1206), .B2(new_n1035), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1207), .A2(new_n1045), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1031), .A2(new_n1045), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1209), .B(KEYINPUT48), .ZN(new_n1210));
  OAI21_X1  g785(.A(new_n1210), .B1(new_n1196), .B2(new_n1038), .ZN(new_n1211));
  AND3_X1   g786(.A1(new_n1204), .A2(new_n1208), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1195), .A2(new_n1212), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g788(.A1(new_n1003), .A2(new_n1009), .ZN(new_n1215));
  INV_X1    g789(.A(G229), .ZN(new_n1216));
  NAND3_X1  g790(.A1(new_n1215), .A2(G319), .A3(new_n1216), .ZN(new_n1217));
  NAND3_X1  g791(.A1(new_n932), .A2(new_n671), .A3(new_n687), .ZN(new_n1218));
  NOR2_X1   g792(.A1(new_n1217), .A2(new_n1218), .ZN(G308));
  AND3_X1   g793(.A1(new_n932), .A2(new_n671), .A3(new_n687), .ZN(new_n1220));
  NAND4_X1  g794(.A1(new_n1220), .A2(G319), .A3(new_n1216), .A4(new_n1215), .ZN(G225));
endmodule


