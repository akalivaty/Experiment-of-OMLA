//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 0 1 1 1 0 0 0 0 1 0 1 0 1 1 1 1 0 0 0 0 1 1 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:36 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n561, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n575, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT65), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  OR2_X1    g028(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT67), .Z(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n457), .A2(KEYINPUT68), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n458), .B1(new_n451), .B2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(KEYINPUT68), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(KEYINPUT69), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g044(.A(KEYINPUT69), .B1(new_n465), .B2(new_n467), .ZN(new_n470));
  OAI21_X1  g045(.A(G125), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n463), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n464), .A2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G101), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(new_n466), .A3(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(KEYINPUT70), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n463), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(G137), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n475), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n473), .A2(new_n482), .ZN(G160));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n485));
  INV_X1    g060(.A(G136), .ZN(new_n486));
  INV_X1    g061(.A(G124), .ZN(new_n487));
  OAI211_X1 g062(.A(G2105), .B(new_n477), .C1(new_n478), .C2(new_n479), .ZN(new_n488));
  OAI221_X1 g063(.A(new_n485), .B1(new_n480), .B2(new_n486), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  INV_X1    g065(.A(G126), .ZN(new_n491));
  NOR2_X1   g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(new_n463), .B2(G114), .ZN(new_n493));
  OAI22_X1  g068(.A1(new_n488), .A2(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n465), .A2(new_n467), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(new_n468), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT71), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  AOI211_X1 g078(.A(new_n499), .B(G2105), .C1(new_n501), .C2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n498), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT4), .B1(new_n480), .B2(new_n499), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n494), .B1(new_n505), .B2(new_n506), .ZN(G164));
  NAND2_X1  g082(.A1(G75), .A2(G543), .ZN(new_n508));
  AND3_X1   g083(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n509));
  AOI21_X1  g084(.A(KEYINPUT5), .B1(KEYINPUT72), .B2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G62), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n508), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G651), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n517), .A2(new_n519), .A3(G543), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n517), .A2(new_n519), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n511), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT72), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT5), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT6), .B(G651), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n528), .A2(KEYINPUT73), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n523), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G88), .ZN(new_n532));
  OAI221_X1 g107(.A(new_n514), .B1(new_n515), .B2(new_n520), .C1(new_n531), .C2(new_n532), .ZN(G303));
  INV_X1    g108(.A(G303), .ZN(G166));
  AND2_X1   g109(.A1(new_n528), .A2(G63), .ZN(new_n535));
  INV_X1    g110(.A(new_n520), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n535), .A2(G651), .B1(new_n536), .B2(G51), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n523), .A2(G89), .A3(new_n530), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  AND3_X1   g115(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(G168));
  NAND3_X1  g116(.A1(new_n523), .A2(G90), .A3(new_n530), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n536), .A2(G52), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n528), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n545));
  NOR3_X1   g120(.A1(new_n544), .A2(new_n545), .A3(new_n516), .ZN(new_n546));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G64), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n511), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g124(.A(KEYINPUT74), .B1(new_n549), .B2(G651), .ZN(new_n550));
  OAI211_X1 g125(.A(new_n542), .B(new_n543), .C1(new_n546), .C2(new_n550), .ZN(G301));
  INV_X1    g126(.A(G301), .ZN(G171));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n511), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n555), .A2(G651), .B1(G43), .B2(new_n536), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n523), .A2(G81), .A3(new_n530), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(G188));
  INV_X1    g140(.A(G53), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n520), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n523), .A2(G91), .A3(new_n530), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n528), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(new_n516), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(G299));
  NAND3_X1  g148(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(G286));
  INV_X1    g149(.A(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n511), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n576), .A2(G651), .B1(new_n536), .B2(G49), .ZN(new_n577));
  INV_X1    g152(.A(G87), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n531), .B2(new_n578), .ZN(G288));
  INV_X1    g154(.A(KEYINPUT75), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n528), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n581), .B2(new_n516), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G61), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n511), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n585), .A2(KEYINPUT75), .A3(G651), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n536), .A2(G48), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n523), .A2(G86), .A3(new_n530), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n591), .A2(new_n516), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n523), .A2(G85), .A3(new_n530), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n536), .A2(G47), .ZN(new_n594));
  AND3_X1   g169(.A1(new_n593), .A2(KEYINPUT76), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g170(.A(KEYINPUT76), .B1(new_n593), .B2(new_n594), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  INV_X1    g174(.A(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n511), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G651), .B1(G54), .B2(new_n536), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g178(.A1(new_n523), .A2(G92), .A3(new_n530), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(KEYINPUT77), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT77), .ZN(new_n606));
  NAND4_X1  g181(.A1(new_n523), .A2(new_n606), .A3(new_n530), .A4(G92), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(KEYINPUT10), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n605), .A2(new_n610), .A3(new_n607), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n603), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n598), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n598), .B1(new_n612), .B2(G868), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  XOR2_X1   g190(.A(G299), .B(KEYINPUT78), .Z(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G297));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G280));
  XOR2_X1   g193(.A(KEYINPUT79), .B(G559), .Z(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(G860), .B2(new_n619), .ZN(G148));
  NAND2_X1  g195(.A1(new_n612), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n621), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n498), .A2(new_n474), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT12), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2100), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n465), .A2(new_n476), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(new_n467), .ZN(new_n630));
  NAND4_X1  g205(.A1(new_n630), .A2(G123), .A3(G2105), .A4(new_n477), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT80), .ZN(new_n632));
  INV_X1    g207(.A(new_n480), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(G135), .ZN(new_n634));
  NOR2_X1   g209(.A1(G99), .A2(G2105), .ZN(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(new_n463), .B2(G111), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n632), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n628), .A2(new_n638), .ZN(G156));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  XOR2_X1   g217(.A(new_n642), .B(G2438), .Z(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT82), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT14), .ZN(new_n647));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT81), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT16), .Z(new_n650));
  OR2_X1    g225(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2443), .B(G2446), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n647), .A2(new_n650), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n651), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n653), .B1(new_n651), .B2(new_n654), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n641), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n651), .A2(new_n654), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(new_n652), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n660), .A2(new_n640), .A3(new_n655), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n658), .A2(new_n661), .A3(G14), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G401));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2084), .B(G2090), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(new_n668), .A3(KEYINPUT17), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT18), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2072), .B(G2078), .Z(new_n672));
  AOI21_X1  g247(.A(new_n672), .B1(new_n667), .B2(KEYINPUT18), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2096), .B(G2100), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n674), .B(new_n675), .Z(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1956), .B(G2474), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n682), .A2(KEYINPUT83), .ZN(new_n683));
  XOR2_X1   g258(.A(G1971), .B(G1976), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(KEYINPUT83), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n683), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT20), .ZN(new_n688));
  OR2_X1    g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n680), .A2(new_n681), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  OR3_X1    g266(.A1(new_n685), .A2(new_n682), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n687), .A2(new_n688), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n685), .A2(new_n691), .ZN(new_n694));
  NAND4_X1  g269(.A1(new_n689), .A2(new_n692), .A3(new_n693), .A4(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT84), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1991), .B(G1996), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n698), .A2(new_n699), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n679), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n698), .A2(new_n699), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n704), .A2(new_n678), .A3(new_n700), .ZN(new_n705));
  AND2_X1   g280(.A1(new_n703), .A2(new_n705), .ZN(G229));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  NOR2_X1   g282(.A1(G164), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G27), .B2(new_n707), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n710), .A2(G2078), .ZN(new_n711));
  NAND2_X1  g286(.A1(G168), .A2(G16), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G16), .B2(G21), .ZN(new_n713));
  INV_X1    g288(.A(G1966), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT93), .Z(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT31), .B(G11), .ZN(new_n717));
  NAND2_X1  g292(.A1(G171), .A2(G16), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G5), .B2(G16), .ZN(new_n719));
  INV_X1    g294(.A(G1961), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT30), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n722), .A2(G28), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n707), .B1(new_n722), .B2(G28), .ZN(new_n724));
  OAI22_X1  g299(.A1(new_n637), .A2(new_n707), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n714), .B2(new_n713), .ZN(new_n726));
  NAND4_X1  g301(.A1(new_n716), .A2(new_n717), .A3(new_n721), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT94), .ZN(new_n728));
  INV_X1    g303(.A(G16), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G20), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(KEYINPUT23), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT23), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G299), .B2(G16), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n731), .B1(new_n733), .B2(new_n730), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT95), .B(G1956), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT96), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n734), .B(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT88), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G4), .B2(G16), .ZN(new_n739));
  OR3_X1    g314(.A1(new_n738), .A2(G4), .A3(G16), .ZN(new_n740));
  INV_X1    g315(.A(new_n612), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n739), .B(new_n740), .C1(new_n741), .C2(new_n729), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(G1348), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n707), .A2(G26), .ZN(new_n744));
  INV_X1    g319(.A(G128), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n488), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT89), .ZN(new_n747));
  OR2_X1    g322(.A1(G104), .A2(G2105), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n748), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n633), .A2(G140), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n747), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n744), .B1(new_n752), .B2(new_n707), .ZN(new_n753));
  MUX2_X1   g328(.A(new_n744), .B(new_n753), .S(KEYINPUT28), .Z(new_n754));
  INV_X1    g329(.A(G2067), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(G160), .A2(G29), .ZN(new_n757));
  XNOR2_X1  g332(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G34), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n757), .B1(G29), .B2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(G2084), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AND2_X1   g337(.A1(new_n707), .A2(G33), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n633), .A2(G139), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n474), .A2(G103), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT25), .Z(new_n766));
  AOI22_X1  g341(.A1(new_n498), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n764), .B(new_n766), .C1(new_n767), .C2(new_n463), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n763), .B1(new_n768), .B2(G29), .ZN(new_n769));
  INV_X1    g344(.A(G2072), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n760), .A2(new_n761), .ZN(new_n772));
  NOR2_X1   g347(.A1(G29), .A2(G32), .ZN(new_n773));
  NAND3_X1  g348(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT91), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT26), .Z(new_n776));
  NAND2_X1  g351(.A1(new_n474), .A2(G105), .ZN(new_n777));
  INV_X1    g352(.A(G141), .ZN(new_n778));
  INV_X1    g353(.A(G129), .ZN(new_n779));
  OAI221_X1 g354(.A(new_n777), .B1(new_n480), .B2(new_n778), .C1(new_n779), .C2(new_n488), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n773), .B1(new_n781), .B2(G29), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT27), .B(G1996), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT92), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n762), .A2(new_n771), .A3(new_n772), .A4(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n729), .A2(G19), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n559), .B2(new_n729), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1341), .ZN(new_n789));
  OAI22_X1  g364(.A1(new_n782), .A2(new_n784), .B1(new_n769), .B2(new_n770), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n707), .A2(G35), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G162), .B2(new_n707), .ZN(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT29), .B(G2090), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR4_X1   g369(.A1(new_n786), .A2(new_n789), .A3(new_n790), .A4(new_n794), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n720), .A2(new_n719), .B1(new_n710), .B2(G2078), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n756), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g372(.A1(new_n728), .A2(new_n737), .A3(new_n743), .A4(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(G288), .B(KEYINPUT86), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(G16), .ZN(new_n800));
  INV_X1    g375(.A(G23), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(G16), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT33), .B(G1976), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n729), .A2(G22), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G166), .B2(new_n729), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n802), .A2(new_n804), .B1(G1971), .B2(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n807), .A2(G1971), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n729), .A2(G6), .ZN(new_n810));
  INV_X1    g385(.A(G305), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(new_n729), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT32), .B(G1981), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n805), .A2(new_n808), .A3(new_n809), .A4(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT87), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n815), .A2(new_n816), .A3(KEYINPUT34), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n816), .B1(new_n815), .B2(KEYINPUT34), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT36), .ZN(new_n821));
  OR2_X1    g396(.A1(G95), .A2(G2105), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n822), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n823));
  INV_X1    g398(.A(G131), .ZN(new_n824));
  INV_X1    g399(.A(G119), .ZN(new_n825));
  OAI221_X1 g400(.A(new_n823), .B1(new_n480), .B2(new_n824), .C1(new_n825), .C2(new_n488), .ZN(new_n826));
  MUX2_X1   g401(.A(G25), .B(new_n826), .S(G29), .Z(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT85), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT35), .B(G1991), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n815), .A2(KEYINPUT34), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n729), .A2(G24), .ZN(new_n832));
  INV_X1    g407(.A(G290), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(new_n729), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(G1986), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n831), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n820), .A2(new_n821), .A3(new_n830), .A4(new_n836), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n836), .B(new_n830), .C1(new_n819), .C2(new_n818), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT36), .ZN(new_n839));
  AOI211_X1 g414(.A(new_n711), .B(new_n798), .C1(new_n837), .C2(new_n839), .ZN(G311));
  AOI21_X1  g415(.A(new_n798), .B1(new_n837), .B2(new_n839), .ZN(new_n841));
  INV_X1    g416(.A(new_n711), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(G150));
  NAND2_X1  g418(.A1(G80), .A2(G543), .ZN(new_n844));
  INV_X1    g419(.A(G67), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n844), .B1(new_n511), .B2(new_n845), .ZN(new_n846));
  AOI22_X1  g421(.A1(new_n846), .A2(G651), .B1(G55), .B2(new_n536), .ZN(new_n847));
  INV_X1    g422(.A(G93), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(new_n848), .B2(new_n531), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT100), .B(KEYINPUT37), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n612), .A2(G559), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n531), .A2(new_n848), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n846), .A2(G651), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n536), .A2(G55), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g432(.A(KEYINPUT98), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT98), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n847), .B(new_n859), .C1(new_n848), .C2(new_n531), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(new_n559), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n849), .A2(KEYINPUT98), .A3(new_n558), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n853), .B(new_n863), .ZN(new_n864));
  XOR2_X1   g439(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n866), .A2(KEYINPUT39), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n867), .A2(KEYINPUT99), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(KEYINPUT99), .ZN(new_n869));
  OR3_X1    g444(.A1(new_n868), .A2(new_n869), .A3(G860), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n866), .A2(KEYINPUT39), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n852), .B1(new_n870), .B2(new_n871), .ZN(G145));
  NAND2_X1  g447(.A1(new_n633), .A2(G142), .ZN(new_n873));
  INV_X1    g448(.A(G130), .ZN(new_n874));
  NOR2_X1   g449(.A1(G106), .A2(G2105), .ZN(new_n875));
  OAI21_X1  g450(.A(G2104), .B1(new_n463), .B2(G118), .ZN(new_n876));
  OAI221_X1 g451(.A(new_n873), .B1(new_n874), .B2(new_n488), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n826), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n878), .A2(new_n879), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(new_n626), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n626), .ZN(new_n884));
  INV_X1    g459(.A(new_n882), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n884), .B1(new_n885), .B2(new_n880), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n630), .A2(G138), .A3(new_n463), .A4(new_n477), .ZN(new_n887));
  AOI22_X1  g462(.A1(new_n887), .A2(KEYINPUT4), .B1(new_n498), .B2(new_n504), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n888), .A2(new_n889), .A3(new_n494), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n505), .A2(new_n506), .ZN(new_n891));
  INV_X1    g466(.A(new_n494), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT102), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n781), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n894), .A2(new_n895), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n752), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n898), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n900), .A2(new_n896), .A3(new_n751), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT103), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n768), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n899), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n768), .B(KEYINPUT103), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n907), .B1(new_n899), .B2(new_n901), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n883), .B(new_n886), .C1(new_n905), .C2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n899), .A2(new_n901), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n906), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n886), .A2(new_n883), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(new_n912), .A3(new_n904), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n909), .A2(KEYINPUT105), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n489), .B(KEYINPUT101), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(G160), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n916), .B(new_n637), .ZN(new_n917));
  INV_X1    g492(.A(new_n912), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n918), .B(new_n919), .C1(new_n905), .C2(new_n908), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n914), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G37), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n917), .B1(new_n913), .B2(new_n923), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT106), .A4(new_n904), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n924), .A2(new_n909), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n921), .A2(new_n922), .A3(new_n926), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g503(.A1(G290), .A2(G166), .ZN(new_n929));
  OAI211_X1 g504(.A(G303), .B(new_n592), .C1(new_n595), .C2(new_n596), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n799), .ZN(new_n932));
  INV_X1    g507(.A(new_n799), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(new_n929), .A3(new_n930), .ZN(new_n934));
  AND3_X1   g509(.A1(new_n932), .A2(new_n811), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n811), .B1(new_n932), .B2(new_n934), .ZN(new_n936));
  OR2_X1    g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(new_n938), .A3(KEYINPUT42), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n935), .A2(new_n936), .ZN(new_n940));
  OR2_X1    g515(.A1(new_n938), .A2(KEYINPUT42), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n938), .A2(KEYINPUT42), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n569), .A2(KEYINPUT107), .A3(new_n570), .A4(new_n572), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n605), .A2(new_n610), .A3(new_n607), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n610), .B1(new_n605), .B2(new_n607), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n602), .B(new_n945), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n949));
  NAND2_X1  g524(.A1(G299), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n609), .A2(new_n611), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n953), .A2(new_n602), .A3(new_n950), .A4(new_n945), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n952), .A2(new_n954), .A3(KEYINPUT108), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n621), .B(new_n863), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT108), .B1(new_n952), .B2(new_n954), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n956), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT41), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n950), .B1(new_n612), .B2(new_n945), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n948), .A2(new_n951), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n952), .A2(new_n954), .A3(KEYINPUT41), .ZN(new_n965));
  AND2_X1   g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n960), .B1(new_n966), .B2(new_n957), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n944), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n939), .A2(new_n967), .A3(new_n943), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(G868), .ZN(new_n972));
  INV_X1    g547(.A(G868), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n849), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(G295));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n972), .A2(new_n976), .A3(new_n974), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n973), .B1(new_n969), .B2(new_n970), .ZN(new_n978));
  INV_X1    g553(.A(new_n974), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT110), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n980), .ZN(G331));
  NAND2_X1  g556(.A1(G301), .A2(G168), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n545), .B1(new_n544), .B2(new_n516), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n549), .A2(KEYINPUT74), .A3(G651), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g560(.A1(G286), .A2(new_n985), .A3(new_n542), .A4(new_n543), .ZN(new_n986));
  AND2_X1   g561(.A1(new_n982), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n863), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n982), .A2(new_n986), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n989), .A2(new_n862), .A3(new_n861), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n991), .B1(new_n955), .B2(new_n958), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT114), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n987), .A2(new_n863), .A3(KEYINPUT112), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT112), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n988), .A2(new_n990), .A3(new_n995), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n964), .A2(new_n994), .A3(new_n965), .A4(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT114), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n998), .B(new_n991), .C1(new_n955), .C2(new_n958), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n993), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n1000), .A2(new_n937), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n988), .A2(new_n990), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n964), .A2(new_n965), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(KEYINPUT111), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n996), .A2(new_n994), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(new_n952), .A3(new_n954), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n964), .A2(new_n1007), .A3(new_n965), .A4(new_n1002), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1004), .A2(new_n1006), .A3(new_n940), .A4(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n922), .ZN(new_n1010));
  OAI21_X1  g585(.A(KEYINPUT43), .B1(new_n1001), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1011), .A2(KEYINPUT115), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1004), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1013));
  OAI21_X1  g588(.A(KEYINPUT113), .B1(new_n935), .B2(new_n936), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT43), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1004), .A2(new_n1014), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1016), .A2(new_n1017), .A3(new_n922), .A4(new_n1018), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n1019), .A2(KEYINPUT44), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n1021));
  OAI211_X1 g596(.A(new_n1021), .B(KEYINPUT43), .C1(new_n1001), .C2(new_n1010), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1012), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1000), .A2(new_n937), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1024), .A2(new_n1017), .A3(new_n922), .A4(new_n1009), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1016), .A2(new_n922), .A3(new_n1018), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1025), .B1(new_n1026), .B2(new_n1017), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT44), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1023), .A2(new_n1029), .ZN(G397));
  NOR2_X1   g605(.A1(G164), .A2(G1384), .ZN(new_n1031));
  INV_X1    g606(.A(G40), .ZN(new_n1032));
  NOR3_X1   g607(.A1(new_n473), .A2(new_n1032), .A3(new_n482), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g609(.A(KEYINPUT58), .B(G1341), .Z(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1384), .ZN(new_n1037));
  OAI211_X1 g612(.A(KEYINPUT45), .B(new_n1037), .C1(new_n890), .C2(new_n893), .ZN(new_n1038));
  INV_X1    g613(.A(new_n482), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n498), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n1040));
  OAI211_X1 g615(.A(G40), .B(new_n1039), .C1(new_n1040), .C2(new_n463), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1037), .B1(new_n888), .B2(new_n494), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT45), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1041), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1038), .A2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1036), .B1(new_n1045), .B2(G1996), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n559), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT59), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1046), .A2(new_n1049), .A3(new_n559), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1034), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1053));
  XOR2_X1   g628(.A(KEYINPUT116), .B(KEYINPUT50), .Z(new_n1054));
  OAI211_X1 g629(.A(new_n1037), .B(new_n1054), .C1(new_n888), .C2(new_n494), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1053), .A2(new_n1055), .A3(new_n1033), .ZN(new_n1056));
  INV_X1    g631(.A(G1348), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1052), .A2(new_n755), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1059), .A2(new_n612), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1058), .A2(new_n741), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT60), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OR3_X1    g637(.A1(new_n1059), .A2(KEYINPUT60), .A3(new_n741), .ZN(new_n1063));
  XNOR2_X1  g638(.A(KEYINPUT56), .B(G2072), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1038), .A2(new_n1044), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1956), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1033), .B1(new_n1042), .B2(KEYINPUT50), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1031), .A2(new_n1054), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1066), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1065), .A2(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g645(.A(G299), .B(KEYINPUT57), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1071), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1065), .A2(new_n1073), .A3(new_n1069), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1072), .A2(KEYINPUT61), .A3(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1051), .A2(new_n1062), .A3(new_n1063), .A4(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1074), .A2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1073), .A2(new_n1065), .A3(new_n1069), .A4(KEYINPUT120), .ZN(new_n1079));
  AND2_X1   g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT61), .B1(new_n1080), .B2(new_n1072), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1061), .B1(new_n1071), .B2(new_n1070), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1083));
  OAI22_X1  g658(.A1(new_n1076), .A2(new_n1081), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G2078), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1038), .A2(new_n1085), .A3(new_n1044), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1086), .A2(new_n1087), .B1(new_n720), .B2(new_n1056), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(G2078), .ZN(new_n1089));
  OAI211_X1 g664(.A(KEYINPUT45), .B(new_n1037), .C1(new_n888), .C2(new_n494), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1044), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT54), .B1(new_n1092), .B2(G171), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n482), .A2(KEYINPUT123), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1032), .B1(new_n482), .B2(KEYINPUT123), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1038), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n473), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1043), .B1(new_n894), .B2(G1384), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1089), .ZN(new_n1099));
  AOI21_X1  g674(.A(G301), .B1(new_n1099), .B2(new_n1088), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1093), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT50), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1041), .B1(new_n1031), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G2090), .ZN(new_n1105));
  OAI211_X1 g680(.A(new_n1104), .B(new_n1105), .C1(new_n1031), .C2(new_n1054), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1038), .A2(new_n1044), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1102), .B(new_n1106), .C1(new_n1107), .C2(G1971), .ZN(new_n1108));
  AOI21_X1  g683(.A(G1971), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1109));
  NOR3_X1   g684(.A1(new_n1067), .A2(new_n1068), .A3(G2090), .ZN(new_n1110));
  OAI21_X1  g685(.A(KEYINPUT119), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1108), .A2(new_n1111), .A3(G8), .ZN(new_n1112));
  NAND2_X1  g687(.A1(G303), .A2(G8), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1113), .B(KEYINPUT55), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1114), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1056), .A2(G2090), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1117), .B(G8), .C1(new_n1109), .C2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(KEYINPUT117), .B1(new_n1034), .B2(G8), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n1121));
  INV_X1    g696(.A(G8), .ZN(new_n1122));
  AOI211_X1 g697(.A(new_n1121), .B(new_n1122), .C1(new_n1031), .C2(new_n1033), .ZN(new_n1123));
  INV_X1    g698(.A(G1976), .ZN(new_n1124));
  OAI22_X1  g699(.A1(new_n1120), .A2(new_n1123), .B1(new_n1124), .B2(new_n799), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT52), .ZN(new_n1126));
  OAI21_X1  g701(.A(G8), .B1(new_n1042), .B2(new_n1041), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(new_n1121), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1034), .A2(KEYINPUT117), .A3(G8), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(G305), .A2(G1981), .ZN(new_n1131));
  INV_X1    g706(.A(G1981), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n587), .A2(new_n1132), .A3(new_n588), .A4(new_n589), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1131), .A2(KEYINPUT49), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT49), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AOI211_X1 g713(.A(KEYINPUT118), .B(KEYINPUT49), .C1(new_n1131), .C2(new_n1133), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1130), .B(new_n1134), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT52), .B1(G288), .B2(new_n1124), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1130), .B(new_n1141), .C1(new_n1124), .C2(new_n799), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1119), .A2(new_n1126), .A3(new_n1140), .A4(new_n1142), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1101), .A2(new_n1116), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1092), .A2(G171), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1099), .A2(new_n1088), .A3(G301), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT54), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1043), .B1(G164), .B2(G1384), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1148), .A2(new_n1090), .A3(new_n1033), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n714), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1053), .A2(new_n1055), .A3(new_n1033), .A4(new_n761), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT51), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1152), .A2(new_n1153), .A3(G8), .ZN(new_n1154));
  NOR2_X1   g729(.A1(G168), .A2(new_n1122), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1154), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT121), .B1(new_n1152), .B2(G8), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n1160));
  AOI211_X1 g735(.A(new_n1160), .B(new_n1122), .C1(new_n1150), .C2(new_n1151), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1155), .A2(KEYINPUT122), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1159), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1158), .B1(new_n1164), .B2(new_n1153), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1147), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1084), .A2(new_n1144), .A3(new_n1167), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n1154), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1152), .A2(G8), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n1160), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1152), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1171), .A2(new_n1162), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1169), .B1(new_n1173), .B2(KEYINPUT51), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1166), .ZN(new_n1175));
  OAI21_X1  g750(.A(KEYINPUT62), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT62), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1165), .A2(new_n1177), .A3(new_n1166), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1116), .A2(new_n1143), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1145), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1176), .A2(new_n1178), .A3(new_n1179), .A4(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(G288), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1140), .A2(new_n1124), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(new_n1133), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(new_n1130), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1119), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1186), .A2(new_n1126), .A3(new_n1140), .A4(new_n1142), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  AND4_X1   g763(.A1(new_n1119), .A2(new_n1126), .A3(new_n1140), .A4(new_n1142), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1170), .A2(G286), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1189), .A2(new_n1115), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT63), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  OAI21_X1  g768(.A(G8), .B1(new_n1109), .B2(new_n1118), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1192), .B1(new_n1194), .B2(new_n1114), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1189), .A2(new_n1190), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1188), .B1(new_n1193), .B2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1168), .A2(new_n1181), .A3(new_n1197), .ZN(new_n1198));
  OAI211_X1 g773(.A(new_n1043), .B(new_n1033), .C1(new_n894), .C2(G1384), .ZN(new_n1199));
  INV_X1    g774(.A(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n751), .B(G2067), .ZN(new_n1201));
  INV_X1    g776(.A(G1996), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n781), .B(new_n1202), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1201), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n826), .A2(new_n829), .ZN(new_n1205));
  OR2_X1    g780(.A1(new_n826), .A2(new_n829), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(new_n1207), .ZN(new_n1208));
  INV_X1    g783(.A(G1986), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1208), .B1(new_n1209), .B2(new_n833), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n833), .A2(new_n1209), .ZN(new_n1211));
  INV_X1    g786(.A(new_n1211), .ZN(new_n1212));
  OAI21_X1  g787(.A(new_n1200), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1198), .A2(new_n1213), .ZN(new_n1214));
  OR3_X1    g789(.A1(new_n1208), .A2(KEYINPUT125), .A3(new_n1199), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1200), .A2(new_n1212), .ZN(new_n1216));
  XNOR2_X1  g791(.A(new_n1216), .B(KEYINPUT48), .ZN(new_n1217));
  OAI21_X1  g792(.A(KEYINPUT125), .B1(new_n1208), .B2(new_n1199), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n1215), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  OAI211_X1 g794(.A(new_n1200), .B(new_n1202), .C1(KEYINPUT124), .C2(KEYINPUT46), .ZN(new_n1220));
  XNOR2_X1  g795(.A(KEYINPUT124), .B(KEYINPUT46), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1221), .B1(new_n1199), .B2(G1996), .ZN(new_n1222));
  OAI21_X1  g797(.A(new_n1200), .B1(new_n895), .B2(new_n1201), .ZN(new_n1223));
  NAND3_X1  g798(.A1(new_n1220), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  XNOR2_X1  g799(.A(new_n1224), .B(KEYINPUT47), .ZN(new_n1225));
  INV_X1    g800(.A(new_n1204), .ZN(new_n1226));
  OAI22_X1  g801(.A1(new_n1226), .A2(new_n1206), .B1(G2067), .B2(new_n751), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1227), .A2(new_n1200), .ZN(new_n1228));
  NAND3_X1  g803(.A1(new_n1219), .A2(new_n1225), .A3(new_n1228), .ZN(new_n1229));
  XNOR2_X1  g804(.A(new_n1229), .B(KEYINPUT126), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1214), .A2(new_n1230), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g806(.A(new_n461), .B1(new_n703), .B2(new_n705), .ZN(new_n1233));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n1234));
  AND2_X1   g808(.A1(new_n662), .A2(new_n676), .ZN(new_n1235));
  AND3_X1   g809(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  AOI21_X1  g810(.A(new_n1234), .B1(new_n1233), .B2(new_n1235), .ZN(new_n1237));
  OR2_X1    g811(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  AND3_X1   g812(.A1(new_n1238), .A2(new_n1027), .A3(new_n927), .ZN(G308));
  NAND3_X1  g813(.A1(new_n1238), .A2(new_n1027), .A3(new_n927), .ZN(G225));
endmodule


