//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT0), .Z(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G116), .A2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n214), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(KEYINPUT65), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AND2_X1   g0020(.A1(new_n218), .A2(new_n219), .ZN(new_n221));
  AOI211_X1 g0021(.A(new_n220), .B(new_n221), .C1(G107), .C2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(G58), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  INV_X1    g0024(.A(G87), .ZN(new_n225));
  INV_X1    g0025(.A(G250), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G97), .ZN(new_n228));
  INV_X1    g0028(.A(G257), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n210), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT1), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  INV_X1    g0033(.A(G20), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n204), .A2(G50), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  AOI211_X1 g0037(.A(new_n213), .B(new_n232), .C1(new_n235), .C2(new_n237), .ZN(G361));
  XOR2_X1   g0038(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n239));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G226), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G250), .B(G257), .Z(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G68), .B(G77), .Z(new_n251));
  XNOR2_X1  g0051(.A(G50), .B(G58), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n250), .B(new_n253), .ZN(G351));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n233), .ZN(new_n256));
  XOR2_X1   g0056(.A(KEYINPUT8), .B(G58), .Z(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n257), .A2(new_n259), .B1(G150), .B2(new_n260), .ZN(new_n261));
  XNOR2_X1  g0061(.A(new_n261), .B(KEYINPUT68), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n205), .A2(new_n234), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n256), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(new_n216), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n255), .A2(new_n233), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n269), .B1(G1), .B2(new_n234), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G50), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n264), .A2(new_n268), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT9), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n264), .A2(KEYINPUT9), .A3(new_n268), .A4(new_n272), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n265), .B(G274), .C1(G41), .C2(G45), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  OAI211_X1 g0078(.A(G1), .B(G13), .C1(new_n258), .C2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n277), .B1(new_n281), .B2(new_n217), .ZN(new_n282));
  OR2_X1    g0082(.A1(new_n282), .A2(KEYINPUT67), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT3), .B(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G222), .A2(G1698), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(G223), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n284), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n279), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n288), .B(new_n289), .C1(G77), .C2(new_n284), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n282), .A2(KEYINPUT67), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n283), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G200), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n275), .A2(new_n276), .A3(new_n293), .A4(new_n295), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n296), .A2(KEYINPUT10), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(KEYINPUT10), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OR3_X1    g0099(.A1(new_n292), .A2(KEYINPUT69), .A3(G179), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n292), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT69), .B1(new_n292), .B2(G179), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n300), .A2(new_n273), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n257), .A2(new_n260), .B1(G20), .B2(G77), .ZN(new_n305));
  INV_X1    g0105(.A(new_n259), .ZN(new_n306));
  XOR2_X1   g0106(.A(KEYINPUT15), .B(G87), .Z(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n305), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n309), .A2(new_n256), .B1(new_n206), .B2(new_n267), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(new_n206), .B2(new_n270), .ZN(new_n311));
  NOR2_X1   g0111(.A1(G232), .A2(G1698), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n286), .A2(G238), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n284), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n314), .B(new_n289), .C1(G107), .C2(new_n284), .ZN(new_n315));
  INV_X1    g0115(.A(G244), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n315), .B(new_n277), .C1(new_n316), .C2(new_n281), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n311), .B1(G200), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n318), .B1(new_n294), .B2(new_n317), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n299), .A2(new_n304), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT14), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT70), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n277), .B(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G238), .ZN(new_n324));
  NOR2_X1   g0124(.A1(G226), .A2(G1698), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n325), .B1(new_n224), .B2(G1698), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n326), .A2(new_n284), .B1(G33), .B2(G97), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n323), .B1(new_n281), .B2(new_n324), .C1(new_n327), .C2(new_n279), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n328), .A2(KEYINPUT13), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(KEYINPUT13), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n321), .B1(new_n331), .B2(G169), .ZN(new_n332));
  AOI211_X1 g0132(.A(KEYINPUT14), .B(new_n301), .C1(new_n329), .C2(new_n330), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G179), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G68), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n267), .A2(KEYINPUT12), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT12), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n341), .B1(new_n266), .B2(G68), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n340), .B(new_n342), .C1(new_n270), .C2(new_n339), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT71), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n343), .B(new_n344), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n259), .A2(G77), .B1(G20), .B2(new_n339), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n260), .A2(G50), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n269), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  XOR2_X1   g0148(.A(new_n348), .B(KEYINPUT11), .Z(new_n349));
  INV_X1    g0149(.A(KEYINPUT72), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n345), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n350), .B1(new_n345), .B2(new_n349), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n338), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n317), .A2(new_n301), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n311), .B(new_n356), .C1(G179), .C2(new_n317), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n331), .A2(G200), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n329), .A2(G190), .A3(new_n330), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n359), .B(new_n360), .C1(new_n352), .C2(new_n353), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  AND2_X1   g0162(.A1(G58), .A2(G68), .ZN(new_n363));
  OAI21_X1  g0163(.A(G20), .B1(new_n363), .B2(new_n203), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT74), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n260), .A2(G159), .ZN(new_n367));
  OAI211_X1 g0167(.A(KEYINPUT74), .B(G20), .C1(new_n363), .C2(new_n203), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT3), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT73), .B1(new_n371), .B2(G33), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(G33), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n371), .A2(KEYINPUT73), .A3(G33), .ZN(new_n375));
  AOI21_X1  g0175(.A(G20), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT7), .ZN(new_n377));
  OAI21_X1  g0177(.A(G68), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n371), .A2(KEYINPUT73), .A3(G33), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n379), .B1(new_n373), .B2(new_n372), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n380), .A2(KEYINPUT7), .A3(G20), .ZN(new_n381));
  OAI211_X1 g0181(.A(KEYINPUT16), .B(new_n370), .C1(new_n378), .C2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT75), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT16), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n377), .B1(new_n284), .B2(G20), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n373), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n388), .A2(KEYINPUT7), .A3(new_n234), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n339), .B1(new_n386), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n385), .B1(new_n390), .B2(new_n369), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT7), .B1(new_n380), .B2(G20), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n376), .A2(new_n377), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(new_n393), .A3(G68), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n394), .A2(KEYINPUT75), .A3(KEYINPUT16), .A4(new_n370), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n384), .A2(new_n256), .A3(new_n391), .A4(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n257), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n266), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n271), .B2(new_n397), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n286), .A2(G223), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT73), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(KEYINPUT3), .B2(new_n258), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n375), .B(new_n401), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT76), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G33), .A2(G87), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT76), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n374), .A2(new_n408), .A3(new_n375), .A4(new_n401), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n374), .A2(G226), .A3(G1698), .A4(new_n375), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n406), .A2(new_n407), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n289), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT77), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT78), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n281), .B2(new_n224), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n279), .A2(KEYINPUT78), .A3(G232), .A4(new_n280), .ZN(new_n417));
  AND3_X1   g0217(.A1(new_n416), .A2(new_n277), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n411), .A2(KEYINPUT77), .A3(new_n289), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n414), .A2(new_n335), .A3(new_n418), .A4(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n412), .A2(new_n418), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n301), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(KEYINPUT18), .B1(new_n400), .B2(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n414), .A2(new_n294), .A3(new_n418), .A4(new_n419), .ZN(new_n425));
  INV_X1    g0225(.A(G200), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n421), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n400), .A2(KEYINPUT17), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT17), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n425), .A2(new_n427), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n396), .A2(new_n399), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n420), .A2(new_n422), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT18), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(new_n435), .A3(new_n432), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n424), .A2(new_n429), .A3(new_n433), .A4(new_n436), .ZN(new_n437));
  NOR4_X1   g0237(.A1(new_n320), .A2(new_n358), .A3(new_n362), .A4(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n387), .A2(new_n373), .A3(G250), .A4(G1698), .ZN(new_n439));
  XNOR2_X1  g0239(.A(new_n439), .B(KEYINPUT82), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G33), .A2(G283), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT81), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT81), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n443), .A2(G33), .A3(G283), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT4), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n316), .A2(G1698), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n374), .A2(new_n446), .A3(new_n375), .A4(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n447), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT4), .B1(new_n388), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n440), .A2(new_n445), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n289), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT86), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n265), .A2(G45), .A3(G274), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT83), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT5), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G41), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n455), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT84), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT83), .B1(new_n457), .B2(G41), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n457), .A2(G41), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n459), .A2(new_n460), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n455), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n456), .A2(new_n278), .A3(KEYINPUT5), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n464), .A2(new_n461), .A3(new_n465), .A4(new_n462), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT84), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n462), .A2(new_n265), .A3(G45), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n279), .B(G257), .C1(new_n469), .C2(new_n458), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n453), .A2(new_n454), .A3(new_n471), .ZN(new_n472));
  AOI22_X1  g0272(.A1(new_n448), .A2(new_n450), .B1(new_n444), .B2(new_n442), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n279), .B1(new_n473), .B2(new_n440), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n468), .A2(new_n470), .ZN(new_n475));
  OAI21_X1  g0275(.A(KEYINPUT86), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(KEYINPUT85), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT85), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n468), .A2(new_n479), .A3(new_n470), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n453), .A3(new_n480), .ZN(new_n481));
  AOI22_X1  g0281(.A1(new_n477), .A2(G190), .B1(G200), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n228), .A2(KEYINPUT79), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT79), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G97), .ZN(new_n485));
  INV_X1    g0285(.A(G107), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n483), .A2(new_n485), .A3(KEYINPUT6), .A4(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT80), .ZN(new_n488));
  XNOR2_X1  g0288(.A(KEYINPUT79), .B(G97), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT80), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT6), .A4(new_n486), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT6), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n228), .A2(new_n486), .ZN(new_n493));
  NOR2_X1   g0293(.A1(G97), .A2(G107), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n488), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G20), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n284), .A2(new_n377), .A3(G20), .ZN(new_n499));
  AOI21_X1  g0299(.A(KEYINPUT7), .B1(new_n388), .B2(new_n234), .ZN(new_n500));
  OAI21_X1  g0300(.A(G107), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n260), .A2(G77), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n256), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n269), .B(new_n266), .C1(G1), .C2(new_n258), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G97), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n266), .A2(G97), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n504), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n478), .A2(new_n453), .A3(new_n335), .A4(new_n480), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n472), .A2(new_n476), .A3(new_n301), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n482), .A2(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n374), .A2(new_n234), .A3(G87), .A4(new_n375), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT22), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT22), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n284), .A2(new_n518), .A3(new_n234), .A4(G87), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n234), .A2(G33), .A3(G116), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n234), .A2(G107), .ZN(new_n522));
  XNOR2_X1  g0322(.A(new_n522), .B(KEYINPUT23), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT24), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n520), .A2(KEYINPUT24), .A3(new_n521), .A4(new_n523), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n256), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n506), .A2(G107), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n267), .A2(new_n486), .ZN(new_n530));
  XNOR2_X1  g0330(.A(new_n530), .B(KEYINPUT25), .ZN(new_n531));
  INV_X1    g0331(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n528), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n463), .A2(new_n467), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n226), .A2(new_n286), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n229), .A2(G1698), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n374), .A2(new_n375), .A3(new_n536), .A4(new_n537), .ZN(new_n538));
  XOR2_X1   g0338(.A(KEYINPUT92), .B(G294), .Z(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G33), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n279), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n279), .B(G264), .C1(new_n469), .C2(new_n458), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n535), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G190), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n541), .A2(new_n543), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n468), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G200), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n534), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n515), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT89), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n505), .A2(new_n308), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT87), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n484), .A2(G97), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n228), .A2(KEYINPUT79), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n225), .B(new_n486), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n234), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT19), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n259), .A2(new_n483), .A3(new_n485), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n556), .A2(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n374), .A2(new_n234), .A3(G68), .A4(new_n375), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n269), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n307), .A2(new_n266), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n553), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n556), .A2(new_n558), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n560), .A2(new_n559), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n566), .A2(new_n562), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n256), .ZN(new_n569));
  INV_X1    g0369(.A(new_n564), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(KEYINPUT87), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n552), .B1(new_n565), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n374), .A2(new_n375), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n316), .A2(G1698), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(G238), .B2(G1698), .ZN(new_n575));
  INV_X1    g0375(.A(G116), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n573), .A2(new_n575), .B1(new_n258), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n289), .ZN(new_n578));
  INV_X1    g0378(.A(G45), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n279), .B(G250), .C1(G1), .C2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n455), .A3(new_n580), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n581), .A2(new_n301), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n581), .A2(G179), .ZN(new_n583));
  NOR3_X1   g0383(.A1(new_n572), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n565), .A2(new_n571), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n578), .A2(G190), .A3(new_n455), .A4(new_n580), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n506), .A2(G87), .ZN(new_n587));
  XNOR2_X1  g0387(.A(new_n587), .B(KEYINPUT88), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n581), .A2(G200), .ZN(new_n589));
  AND4_X1   g0389(.A1(new_n585), .A2(new_n586), .A3(new_n588), .A4(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n551), .B1(new_n584), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n552), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n585), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n582), .ZN(new_n594));
  INV_X1    g0394(.A(new_n583), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n585), .A2(new_n586), .A3(new_n588), .A4(new_n589), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(KEYINPUT89), .A3(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n591), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n266), .A2(G116), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n505), .A2(new_n576), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n576), .A2(G20), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n256), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(G20), .B1(new_n442), .B2(new_n444), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n483), .A2(new_n485), .A3(new_n258), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n606), .A2(KEYINPUT90), .A3(KEYINPUT20), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT90), .B1(new_n606), .B2(KEYINPUT20), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n606), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT91), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT20), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(KEYINPUT91), .B1(new_n606), .B2(KEYINPUT20), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI211_X1 g0415(.A(new_n600), .B(new_n601), .C1(new_n609), .C2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n388), .A2(G303), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n380), .B1(G257), .B2(G1698), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n286), .A2(G264), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n289), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n279), .B(G270), .C1(new_n469), .C2(new_n458), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n621), .A2(new_n468), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(G200), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n616), .B(new_n624), .C1(new_n294), .C2(new_n623), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT21), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n623), .A2(G169), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n626), .B1(new_n616), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n600), .B1(new_n609), .B2(new_n615), .ZN(new_n629));
  INV_X1    g0429(.A(new_n601), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n535), .B1(new_n620), .B2(new_n289), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n301), .B1(new_n632), .B2(new_n622), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n631), .A2(KEYINPUT21), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n623), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n631), .A2(G179), .A3(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n625), .A2(new_n628), .A3(new_n634), .A4(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT93), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n638), .B1(new_n544), .B2(new_n301), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n547), .A2(KEYINPUT93), .A3(G169), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n544), .A2(G179), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n533), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n637), .A2(new_n644), .ZN(new_n645));
  AND4_X1   g0445(.A1(new_n438), .A2(new_n550), .A3(new_n599), .A4(new_n645), .ZN(G372));
  AND2_X1   g0446(.A1(new_n429), .A2(new_n433), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n358), .A2(new_n647), .A3(new_n361), .ZN(new_n648));
  XNOR2_X1  g0448(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n434), .A2(KEYINPUT95), .A3(new_n432), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT95), .B1(new_n434), .B2(new_n432), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n653), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n655), .A2(new_n651), .A3(new_n649), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n648), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n299), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(new_n304), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n472), .A2(new_n476), .A3(new_n301), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n510), .A2(new_n512), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n591), .A2(new_n663), .A3(new_n598), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT26), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n643), .A2(new_n628), .A3(new_n634), .A4(new_n636), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n666), .A2(new_n515), .A3(new_n549), .A4(new_n597), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n584), .A2(new_n590), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT94), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n661), .B2(new_n662), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT26), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n514), .A2(KEYINPUT94), .A3(new_n512), .A4(new_n510), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n668), .A2(new_n670), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n665), .A2(new_n667), .A3(new_n596), .A4(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n438), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n660), .B1(new_n675), .B2(new_n676), .ZN(G369));
  AND2_X1   g0477(.A1(new_n549), .A2(new_n643), .ZN(new_n678));
  INV_X1    g0478(.A(G13), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(G20), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n265), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n678), .B1(new_n534), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n644), .A2(new_n686), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n628), .A2(new_n634), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n686), .B1(new_n691), .B2(new_n636), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n636), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n616), .A2(new_n687), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n637), .B2(new_n695), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n693), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n686), .B(KEYINPUT97), .ZN(new_n700));
  AOI22_X1  g0500(.A1(new_n692), .A2(new_n678), .B1(new_n644), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g0502(.A(new_n702), .B(KEYINPUT98), .Z(G399));
  INV_X1    g0503(.A(new_n211), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(G41), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G1), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n556), .A2(G116), .ZN(new_n708));
  OAI22_X1  g0508(.A1(new_n707), .A2(new_n708), .B1(new_n236), .B2(new_n706), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n709), .B(KEYINPUT28), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n674), .A2(new_n700), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(KEYINPUT29), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n668), .A2(new_n670), .A3(new_n672), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT26), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n591), .A2(new_n598), .A3(new_n671), .A4(new_n663), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n667), .A2(new_n715), .A3(new_n596), .A4(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n713), .B1(new_n717), .B2(new_n687), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n712), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n550), .A2(new_n645), .A3(new_n599), .A4(new_n700), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT31), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n481), .A2(new_n335), .A3(new_n547), .A4(new_n581), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n635), .ZN(new_n723));
  INV_X1    g0523(.A(new_n581), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n477), .A2(new_n546), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n635), .A2(G179), .ZN(new_n726));
  OR3_X1    g0526(.A1(new_n725), .A2(new_n726), .A3(KEYINPUT30), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT30), .B1(new_n725), .B2(new_n726), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n723), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n721), .B1(new_n729), .B2(new_n687), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n727), .A2(new_n728), .ZN(new_n731));
  INV_X1    g0531(.A(new_n723), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XOR2_X1   g0533(.A(KEYINPUT99), .B(KEYINPUT31), .Z(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n720), .B(new_n730), .C1(new_n735), .C2(new_n700), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G330), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n719), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n710), .B1(new_n739), .B2(G1), .ZN(G364));
  NOR3_X1   g0540(.A1(new_n679), .A2(new_n579), .A3(G20), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n741), .A2(KEYINPUT100), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(KEYINPUT100), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n742), .A2(G1), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n705), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n237), .A2(new_n579), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n380), .A2(new_n704), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n747), .B(new_n748), .C1(new_n253), .C2(new_n579), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n284), .A2(G355), .A3(new_n211), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n749), .B(new_n750), .C1(G116), .C2(new_n211), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G13), .A2(G33), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n233), .B1(G20), .B2(new_n301), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT101), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n746), .B1(new_n751), .B2(new_n759), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT102), .Z(new_n761));
  NOR2_X1   g0561(.A1(new_n234), .A2(new_n294), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n335), .A2(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n234), .A2(G190), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G179), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(G322), .A2(new_n765), .B1(new_n769), .B2(G329), .ZN(new_n770));
  INV_X1    g0570(.A(G326), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n335), .A2(new_n426), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n762), .A2(new_n772), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n770), .B(new_n388), .C1(new_n771), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n426), .A2(G179), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n766), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n774), .B1(G283), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n762), .A2(new_n775), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G303), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n234), .B1(new_n767), .B2(G190), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n539), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n772), .A2(new_n766), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(KEYINPUT33), .B(G317), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n766), .A2(new_n763), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n786), .A2(new_n787), .B1(new_n789), .B2(G311), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n778), .A2(new_n781), .A3(new_n784), .A4(new_n790), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n764), .B(KEYINPUT103), .Z(new_n792));
  INV_X1    g0592(.A(new_n773), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n792), .A2(G58), .B1(G50), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n284), .B1(new_n785), .B2(new_n339), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n788), .A2(new_n206), .B1(new_n782), .B2(new_n228), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n795), .B(new_n796), .C1(G87), .C2(new_n780), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n777), .A2(G107), .ZN(new_n798));
  INV_X1    g0598(.A(G159), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n768), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT104), .B(KEYINPUT32), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n794), .A2(new_n797), .A3(new_n798), .A4(new_n802), .ZN(new_n803));
  AND2_X1   g0603(.A1(new_n791), .A2(new_n803), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n761), .B1(new_n757), .B2(new_n804), .C1(new_n697), .C2(new_n755), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n698), .A2(new_n746), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n697), .A2(G330), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(G396));
  NAND2_X1  g0608(.A1(new_n311), .A2(new_n686), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n319), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n357), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n357), .A2(new_n686), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n711), .B(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n737), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT106), .Z(new_n819));
  AOI21_X1  g0619(.A(new_n745), .B1(new_n817), .B2(new_n737), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n814), .A2(new_n752), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n756), .A2(new_n752), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n745), .B1(G77), .B2(new_n824), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n825), .A2(KEYINPUT105), .ZN(new_n826));
  INV_X1    g0626(.A(G283), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n785), .A2(new_n827), .B1(new_n782), .B2(new_n228), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n828), .B1(G116), .B2(new_n789), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n388), .B1(new_n779), .B2(new_n486), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(G311), .B2(new_n769), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n765), .A2(G294), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G303), .A2(new_n793), .B1(new_n777), .B2(G87), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n829), .A2(new_n831), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G137), .A2(new_n793), .B1(new_n786), .B2(G150), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n799), .B2(new_n788), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G143), .B2(new_n792), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT34), .Z(new_n838));
  NOR2_X1   g0638(.A1(new_n776), .A2(new_n339), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(G50), .B2(new_n780), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n573), .B1(G132), .B2(new_n769), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n838), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n782), .A2(new_n223), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n834), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n756), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n825), .A2(KEYINPUT105), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n822), .A2(new_n826), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n821), .A2(new_n847), .ZN(G384));
  NAND2_X1  g0648(.A1(new_n394), .A2(new_n370), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n385), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n850), .A2(new_n384), .A3(new_n256), .A4(new_n395), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n851), .A2(new_n399), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(new_n423), .B2(new_n684), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n431), .A2(new_n432), .ZN(new_n854));
  OAI21_X1  g0654(.A(KEYINPUT37), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT37), .B1(new_n434), .B2(new_n432), .ZN(new_n856));
  INV_X1    g0656(.A(new_n854), .ZN(new_n857));
  INV_X1    g0657(.A(new_n684), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n432), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT108), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n852), .A2(new_n684), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n437), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n862), .B1(new_n437), .B2(new_n863), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n861), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI211_X1 g0668(.A(KEYINPUT38), .B(new_n861), .C1(new_n864), .C2(new_n865), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n733), .A2(KEYINPUT31), .A3(new_n686), .ZN(new_n871));
  INV_X1    g0671(.A(new_n734), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n729), .B2(new_n687), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n871), .A2(new_n720), .A3(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT107), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n338), .A2(new_n354), .A3(new_n687), .ZN(new_n876));
  INV_X1    g0676(.A(new_n353), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(new_n351), .A3(new_n686), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n361), .A2(new_n878), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n332), .A2(new_n333), .A3(new_n336), .ZN(new_n880));
  INV_X1    g0680(.A(new_n354), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n875), .B1(new_n876), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n876), .A2(new_n882), .A3(new_n875), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n874), .A2(new_n886), .A3(new_n815), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT40), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n870), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n654), .A2(new_n656), .A3(new_n647), .ZN(new_n890));
  INV_X1    g0690(.A(new_n859), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n655), .A2(new_n857), .A3(new_n651), .A4(new_n859), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT37), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n890), .A2(new_n891), .B1(new_n893), .B2(new_n860), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n869), .B1(new_n894), .B2(KEYINPUT38), .ZN(new_n895));
  AND2_X1   g0695(.A1(new_n887), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n889), .B1(new_n896), .B2(new_n888), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(G330), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n438), .A2(new_n874), .A3(G330), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n438), .A2(new_n874), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n898), .A2(new_n899), .B1(new_n901), .B2(new_n897), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n437), .A2(new_n863), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT108), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n437), .A2(new_n862), .A3(new_n863), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT38), .B1(new_n906), .B2(new_n861), .ZN(new_n907));
  INV_X1    g0707(.A(new_n869), .ZN(new_n908));
  OAI21_X1  g0708(.A(KEYINPUT39), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT39), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n869), .B(new_n910), .C1(new_n894), .C2(KEYINPUT38), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n876), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n876), .A2(new_n882), .A3(new_n875), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n913), .A2(new_n883), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n674), .A2(new_n700), .A3(new_n815), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n914), .B1(new_n915), .B2(new_n813), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n907), .B2(new_n908), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n657), .A2(new_n858), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n912), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n902), .B(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n438), .B1(new_n712), .B2(new_n718), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n660), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n922), .B(new_n924), .Z(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n265), .B2(new_n680), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n576), .B1(new_n496), .B2(KEYINPUT35), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n927), .B(new_n235), .C1(KEYINPUT35), .C2(new_n496), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT36), .ZN(new_n929));
  NOR3_X1   g0729(.A1(new_n236), .A2(new_n206), .A3(new_n363), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n202), .A2(new_n339), .ZN(new_n931));
  OAI211_X1 g0731(.A(G1), .B(new_n679), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n926), .A2(new_n929), .A3(new_n932), .ZN(G367));
  NAND2_X1  g0733(.A1(new_n585), .A2(new_n588), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n686), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n668), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n584), .A2(new_n934), .A3(new_n686), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n746), .B1(new_n939), .B2(new_n754), .ZN(new_n940));
  INV_X1    g0740(.A(new_n748), .ZN(new_n941));
  OAI221_X1 g0741(.A(new_n759), .B1(new_n211), .B2(new_n308), .C1(new_n246), .C2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n380), .B1(G311), .B2(new_n793), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n786), .A2(new_n539), .B1(new_n789), .B2(G283), .ZN(new_n944));
  INV_X1    g0744(.A(new_n489), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n943), .B(new_n944), .C1(new_n945), .C2(new_n776), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n792), .A2(G303), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n780), .A2(G116), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT46), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n948), .A2(new_n949), .B1(new_n783), .B2(G107), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n947), .B(new_n950), .C1(new_n949), .C2(new_n948), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n946), .B(new_n951), .C1(G317), .C2(new_n769), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT110), .ZN(new_n953));
  AOI22_X1  g0753(.A1(G58), .A2(new_n780), .B1(new_n769), .B2(G137), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT112), .Z(new_n955));
  OAI21_X1  g0755(.A(new_n284), .B1(new_n785), .B2(new_n799), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n776), .A2(new_n206), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n793), .A2(G143), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n789), .A2(new_n202), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n782), .A2(new_n339), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(G150), .B2(new_n765), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT111), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n953), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT47), .Z(new_n966));
  OAI211_X1 g0766(.A(new_n940), .B(new_n942), .C1(new_n966), .C2(new_n757), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n515), .B1(new_n511), .B2(new_n700), .ZN(new_n968));
  INV_X1    g0768(.A(new_n663), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n969), .A2(new_n700), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n692), .A2(new_n678), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT42), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n969), .B1(new_n968), .B2(new_n643), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT109), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n700), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n974), .A2(new_n977), .B1(KEYINPUT43), .B2(new_n938), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n978), .B(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n699), .A2(new_n971), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n980), .B(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n971), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n701), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT45), .Z(new_n985));
  NOR2_X1   g0785(.A1(new_n983), .A2(new_n701), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT44), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n985), .A2(new_n699), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n693), .A2(new_n698), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n699), .A2(new_n972), .A3(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n988), .A2(new_n739), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n739), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n705), .B(KEYINPUT41), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n744), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n967), .B1(new_n982), .B2(new_n995), .ZN(G387));
  NAND2_X1  g0796(.A1(new_n991), .A2(new_n739), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n706), .B1(new_n990), .B2(new_n738), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n764), .A2(new_n216), .B1(new_n776), .B2(new_n228), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n308), .A2(new_n782), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(G159), .C2(new_n793), .ZN(new_n1002));
  XOR2_X1   g0802(.A(KEYINPUT113), .B(G150), .Z(new_n1003));
  NAND2_X1  g0803(.A1(new_n769), .A2(new_n1003), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n779), .A2(new_n206), .B1(new_n788), .B2(new_n339), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n257), .B2(new_n786), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1002), .A2(new_n380), .A3(new_n1004), .A4(new_n1006), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G311), .A2(new_n786), .B1(new_n789), .B2(G303), .ZN(new_n1008));
  INV_X1    g0808(.A(G322), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1008), .B1(new_n1009), .B2(new_n773), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(G317), .B2(new_n792), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT48), .Z(new_n1012));
  NAND2_X1  g0812(.A1(new_n780), .A2(new_n539), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(new_n827), .C2(new_n782), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT49), .Z(new_n1015));
  OAI221_X1 g0815(.A(new_n573), .B1(new_n576), .B2(new_n776), .C1(new_n771), .C2(new_n768), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1007), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n756), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n257), .A2(new_n216), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT50), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n339), .A2(new_n206), .ZN(new_n1021));
  NOR4_X1   g0821(.A1(new_n1020), .A2(G45), .A3(new_n1021), .A4(new_n708), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n748), .B1(new_n243), .B2(new_n579), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n708), .A2(new_n211), .A3(new_n284), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1022), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n211), .A2(G107), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n759), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n688), .A2(new_n689), .A3(new_n754), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1018), .A2(new_n745), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n744), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n999), .B(new_n1029), .C1(new_n1030), .C2(new_n990), .ZN(G393));
  NAND2_X1  g0831(.A1(new_n971), .A2(new_n754), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G317), .A2(new_n793), .B1(new_n765), .B2(G311), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT52), .Z(new_n1034));
  NAND2_X1  g0834(.A1(new_n789), .A2(G294), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n786), .A2(G303), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n779), .A2(new_n827), .B1(new_n768), .B2(new_n1009), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G116), .B2(new_n783), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1038), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n284), .B(new_n1039), .C1(G107), .C2(new_n777), .ZN(new_n1040));
  INV_X1    g0840(.A(G150), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n773), .A2(new_n1041), .B1(new_n764), .B2(new_n799), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT51), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n782), .A2(new_n206), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G68), .B2(new_n780), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n573), .B1(G143), .B2(new_n769), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n257), .A2(new_n789), .B1(new_n777), .B2(G87), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1043), .A2(new_n1045), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n202), .B2(new_n786), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n756), .B1(new_n1040), .B2(new_n1049), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n759), .B1(new_n211), .B2(new_n945), .C1(new_n250), .C2(new_n941), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1032), .A2(new_n745), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n985), .A2(new_n987), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(new_n699), .Z(new_n1054));
  NAND3_X1  g0854(.A1(new_n1054), .A2(KEYINPUT114), .A3(new_n997), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n705), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1054), .A2(new_n997), .B1(KEYINPUT114), .B2(new_n992), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1052), .B1(new_n1030), .B2(new_n1054), .C1(new_n1056), .C2(new_n1057), .ZN(G390));
  INV_X1    g0858(.A(new_n911), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n910), .B1(new_n868), .B2(new_n869), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n752), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G128), .A2(new_n793), .B1(new_n765), .B2(G132), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT116), .Z(new_n1064));
  XOR2_X1   g0864(.A(KEYINPUT54), .B(G143), .Z(new_n1065));
  AOI21_X1  g0865(.A(new_n1064), .B1(new_n789), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n786), .A2(G137), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n780), .A2(new_n1003), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT53), .Z(new_n1069));
  OAI22_X1  g0869(.A1(new_n776), .A2(new_n201), .B1(new_n782), .B2(new_n799), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n388), .B(new_n1070), .C1(G125), .C2(new_n769), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1066), .A2(new_n1067), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n945), .A2(new_n788), .B1(new_n785), .B2(new_n486), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT117), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1044), .B(new_n839), .C1(G283), .C2(new_n793), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n388), .B1(new_n779), .B2(new_n225), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT118), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n769), .A2(G294), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1073), .A2(new_n1074), .B1(G116), .B2(new_n765), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1076), .A2(new_n1078), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1072), .B1(new_n1075), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n756), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n823), .A2(new_n397), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n1062), .A2(new_n745), .A3(new_n1083), .A4(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n717), .A2(new_n687), .A3(new_n811), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n813), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n886), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1088), .A2(new_n876), .A3(new_n895), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n736), .A2(G330), .A3(new_n886), .A4(new_n815), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n909), .A2(new_n911), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n876), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n916), .A2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1089), .B(new_n1090), .C1(new_n1091), .C2(new_n1093), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n1088), .A2(new_n876), .A3(new_n895), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n915), .A2(new_n813), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n886), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n876), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1095), .B1(new_n1061), .B2(new_n1098), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n815), .A2(G330), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n874), .A2(new_n886), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1094), .B1(new_n1099), .B2(new_n1102), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1103), .A2(new_n1030), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n886), .B1(new_n736), .B2(new_n1100), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1096), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1087), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n874), .A2(new_n1100), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1090), .B(new_n1107), .C1(new_n1108), .C2(new_n886), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n923), .A2(new_n899), .A3(new_n660), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1098), .A2(new_n909), .A3(new_n911), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n1114), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1102), .B1(new_n1114), .B2(new_n1089), .ZN(new_n1116));
  OAI211_X1 g0916(.A(KEYINPUT115), .B(new_n1113), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1111), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1118), .B(new_n1094), .C1(new_n1099), .C2(new_n1102), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1117), .A2(new_n705), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(KEYINPUT115), .B1(new_n1103), .B2(new_n1113), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1085), .B(new_n1104), .C1(new_n1120), .C2(new_n1121), .ZN(G378));
  OAI21_X1  g0922(.A(new_n304), .B1(new_n297), .B2(new_n298), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n273), .A2(new_n858), .ZN(new_n1124));
  AND2_X1   g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  OR3_X1    g0928(.A1(new_n1125), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1128), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n912), .A2(new_n920), .A3(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1092), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n918), .B1(new_n870), .B2(new_n916), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1131), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n898), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1132), .B1(new_n912), .B2(new_n920), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1134), .A2(new_n1135), .A3(new_n1131), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1138), .A2(new_n1139), .A3(G330), .A4(new_n897), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n744), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n824), .A2(new_n202), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n776), .A2(new_n223), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(G77), .A2(new_n780), .B1(new_n765), .B2(G107), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n576), .B2(new_n773), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1144), .B(new_n1146), .C1(new_n307), .C2(new_n789), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n573), .A2(new_n278), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n962), .B(new_n1148), .C1(G283), .C2(new_n769), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1147), .B(new_n1149), .C1(new_n228), .C2(new_n785), .ZN(new_n1150));
  XOR2_X1   g0950(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1151));
  XNOR2_X1  g0951(.A(new_n1150), .B(new_n1151), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1148), .B(new_n216), .C1(G33), .C2(G41), .ZN(new_n1153));
  AOI211_X1 g0953(.A(G33), .B(G41), .C1(new_n769), .C2(G124), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n799), .B2(new_n776), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G132), .A2(new_n786), .B1(new_n789), .B2(G137), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n793), .A2(G125), .B1(new_n783), .B2(G150), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n780), .A2(new_n1065), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n765), .A2(G128), .ZN(new_n1159));
  NAND4_X1  g0959(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .A4(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT59), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1152), .B(new_n1153), .C1(new_n1155), .C2(new_n1161), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n746), .B(new_n1143), .C1(new_n1162), .C2(new_n756), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n1131), .B2(new_n753), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT120), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1142), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1119), .A2(new_n1112), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1141), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n706), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1137), .A2(new_n1140), .B1(new_n1119), .B2(new_n1112), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(KEYINPUT57), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1169), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(G375));
  NAND2_X1  g0977(.A1(new_n914), .A2(new_n752), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1001), .B1(G303), .B2(new_n769), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n228), .B2(new_n779), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n957), .B(new_n1180), .C1(G283), .C2(new_n765), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n793), .A2(G294), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n789), .A2(G107), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n284), .B1(new_n786), .B2(G116), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n779), .A2(new_n799), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n786), .A2(new_n1065), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n1144), .B(new_n1187), .C1(G132), .C2(new_n793), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n792), .A2(G137), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n788), .A2(new_n1041), .B1(new_n782), .B2(new_n216), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n573), .B(new_n1190), .C1(G128), .C2(new_n769), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1188), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1185), .B1(new_n1186), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n756), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n823), .A2(new_n339), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1178), .A2(new_n745), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1196), .B1(new_n1197), .B2(new_n1030), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT121), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n994), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1199), .B1(new_n1118), .B2(new_n1200), .ZN(G381));
  NAND2_X1  g1001(.A1(new_n1103), .A2(new_n1113), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT115), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1204), .A2(new_n705), .A3(new_n1119), .A4(new_n1117), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1205), .A2(KEYINPUT122), .A3(new_n1085), .A4(new_n1104), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT122), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(G378), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1206), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1210), .A2(G375), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(G390), .A2(G387), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(G393), .A2(G396), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  OR3_X1    g1014(.A1(new_n1214), .A2(G384), .A3(G381), .ZN(G407));
  NAND2_X1  g1015(.A1(new_n685), .A2(G213), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT123), .Z(new_n1217));
  INV_X1    g1017(.A(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1211), .A2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(G407), .A2(G213), .A3(new_n1219), .ZN(G409));
  XNOR2_X1  g1020(.A(G393), .B(G396), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(G390), .A2(G387), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1222), .B1(new_n1224), .B2(new_n1212), .ZN(new_n1225));
  OR2_X1    g1025(.A1(G390), .A2(G387), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1226), .A2(new_n1221), .A3(new_n1223), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1168), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1166), .B(new_n1229), .C1(new_n1141), .C2(new_n744), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n994), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1230), .B1(new_n1231), .B2(new_n1171), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1209), .A2(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT124), .B1(new_n1176), .B2(G378), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n705), .B1(new_n1174), .B2(KEYINPUT57), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1141), .A2(KEYINPUT57), .A3(new_n1170), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G378), .B(new_n1230), .C1(new_n1235), .C2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT124), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1233), .B1(new_n1234), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT125), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT60), .B1(new_n1197), .B2(new_n1111), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1241), .B1(new_n1242), .B2(new_n1118), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1244));
  OAI211_X1 g1044(.A(KEYINPUT125), .B(new_n1113), .C1(new_n1244), .C2(KEYINPUT60), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(KEYINPUT60), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1243), .A2(new_n705), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1247), .A2(G384), .A3(new_n1199), .ZN(new_n1248));
  AOI21_X1  g1048(.A(G384), .B1(new_n1247), .B2(new_n1199), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1240), .A2(new_n1216), .A3(new_n1250), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1176), .A2(KEYINPUT124), .A3(G378), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1218), .B1(new_n1255), .B2(new_n1233), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1250), .A2(KEYINPUT62), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1251), .A2(new_n1252), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT61), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1247), .A2(new_n1199), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(new_n821), .A3(new_n847), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1216), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1247), .A2(G384), .A3(new_n1199), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1261), .A2(G2897), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1218), .A2(G2897), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1264), .A2(new_n1266), .A3(KEYINPUT126), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT126), .B1(new_n1264), .B2(new_n1266), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1259), .B1(new_n1270), .B2(new_n1256), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1228), .B1(new_n1258), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT63), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n1248), .A2(new_n1249), .A3(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1228), .B1(new_n1256), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1240), .A2(new_n1216), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT126), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1267), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1273), .B1(new_n1276), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1251), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1259), .B(new_n1275), .C1(new_n1281), .C2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1272), .A2(new_n1283), .ZN(G405));
  OAI21_X1  g1084(.A(new_n1255), .B1(new_n1176), .B2(new_n1210), .ZN(new_n1285));
  OR2_X1    g1085(.A1(new_n1285), .A2(new_n1250), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1250), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1228), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1286), .A2(new_n1225), .A3(new_n1227), .A4(new_n1287), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(G402));
endmodule


