

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578;

  OR2_X1 U321 ( .A1(n565), .A2(n537), .ZN(n343) );
  OR2_X1 U322 ( .A1(n379), .A2(n378), .ZN(n380) );
  XNOR2_X1 U323 ( .A(n328), .B(KEYINPUT31), .ZN(n329) );
  INV_X1 U324 ( .A(KEYINPUT113), .ZN(n381) );
  XNOR2_X1 U325 ( .A(n434), .B(n329), .ZN(n330) );
  XNOR2_X1 U326 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U327 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U328 ( .A(n405), .B(n305), .Z(n551) );
  XNOR2_X1 U329 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U330 ( .A(n451), .B(n450), .ZN(G1349GAT) );
  XOR2_X1 U331 ( .A(KEYINPUT85), .B(KEYINPUT17), .Z(n290) );
  XNOR2_X1 U332 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n289) );
  XNOR2_X1 U333 ( .A(n290), .B(n289), .ZN(n291) );
  XNOR2_X1 U334 ( .A(KEYINPUT19), .B(n291), .ZN(n405) );
  XOR2_X1 U335 ( .A(G176GAT), .B(KEYINPUT20), .Z(n293) );
  XNOR2_X1 U336 ( .A(G169GAT), .B(KEYINPUT84), .ZN(n292) );
  XNOR2_X1 U337 ( .A(n293), .B(n292), .ZN(n304) );
  XOR2_X1 U338 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n295) );
  XOR2_X1 U339 ( .A(G190GAT), .B(G134GAT), .Z(n345) );
  XOR2_X1 U340 ( .A(G120GAT), .B(G71GAT), .Z(n334) );
  XNOR2_X1 U341 ( .A(n345), .B(n334), .ZN(n294) );
  XNOR2_X1 U342 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U343 ( .A(n296), .B(G99GAT), .Z(n302) );
  XNOR2_X1 U344 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n297), .B(G127GAT), .ZN(n420) );
  XOR2_X1 U346 ( .A(n420), .B(G15GAT), .Z(n299) );
  NAND2_X1 U347 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U348 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U349 ( .A(G43GAT), .B(n300), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U351 ( .A(n304), .B(n303), .Z(n305) );
  INV_X1 U352 ( .A(n551), .ZN(n455) );
  XNOR2_X1 U353 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n306) );
  XNOR2_X1 U354 ( .A(n306), .B(G29GAT), .ZN(n307) );
  XOR2_X1 U355 ( .A(n307), .B(KEYINPUT8), .Z(n309) );
  XNOR2_X1 U356 ( .A(G43GAT), .B(G50GAT), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n358) );
  XOR2_X1 U358 ( .A(G169GAT), .B(G8GAT), .Z(n394) );
  XOR2_X1 U359 ( .A(G15GAT), .B(G1GAT), .Z(n364) );
  XOR2_X1 U360 ( .A(n394), .B(n364), .Z(n311) );
  NAND2_X1 U361 ( .A1(G229GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U363 ( .A(G141GAT), .B(G22GAT), .Z(n440) );
  XOR2_X1 U364 ( .A(n312), .B(n440), .Z(n320) );
  XOR2_X1 U365 ( .A(KEYINPUT72), .B(KEYINPUT29), .Z(n314) );
  XNOR2_X1 U366 ( .A(G113GAT), .B(G197GAT), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U368 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n316) );
  XNOR2_X1 U369 ( .A(KEYINPUT71), .B(KEYINPUT69), .ZN(n315) );
  XNOR2_X1 U370 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n358), .B(n321), .ZN(n565) );
  XNOR2_X1 U374 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n341) );
  XOR2_X1 U375 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n323) );
  XNOR2_X1 U376 ( .A(KEYINPUT75), .B(KEYINPUT32), .ZN(n322) );
  XOR2_X1 U377 ( .A(n323), .B(n322), .Z(n340) );
  XOR2_X1 U378 ( .A(KEYINPUT33), .B(KEYINPUT80), .Z(n325) );
  XNOR2_X1 U379 ( .A(KEYINPUT76), .B(KEYINPUT77), .ZN(n324) );
  XNOR2_X1 U380 ( .A(n325), .B(n324), .ZN(n331) );
  XOR2_X1 U381 ( .A(G78GAT), .B(G148GAT), .Z(n327) );
  XNOR2_X1 U382 ( .A(G106GAT), .B(G204GAT), .ZN(n326) );
  XNOR2_X1 U383 ( .A(n327), .B(n326), .ZN(n434) );
  AND2_X1 U384 ( .A1(G230GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n338) );
  XNOR2_X1 U386 ( .A(G57GAT), .B(KEYINPUT74), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n332), .B(KEYINPUT13), .ZN(n363) );
  XNOR2_X1 U388 ( .A(G176GAT), .B(G92GAT), .ZN(n333) );
  XNOR2_X1 U389 ( .A(n333), .B(G64GAT), .ZN(n395) );
  XNOR2_X1 U390 ( .A(n363), .B(n395), .ZN(n336) );
  XOR2_X1 U391 ( .A(G99GAT), .B(G85GAT), .Z(n344) );
  XOR2_X1 U392 ( .A(n334), .B(n344), .Z(n335) );
  XNOR2_X1 U393 ( .A(n340), .B(n339), .ZN(n385) );
  XOR2_X1 U394 ( .A(n341), .B(n385), .Z(n537) );
  XOR2_X1 U395 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n342) );
  XNOR2_X1 U396 ( .A(n343), .B(n342), .ZN(n379) );
  XOR2_X1 U397 ( .A(KEYINPUT9), .B(KEYINPUT81), .Z(n347) );
  XNOR2_X1 U398 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U399 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U400 ( .A(n348), .B(KEYINPUT11), .Z(n353) );
  XOR2_X1 U401 ( .A(G92GAT), .B(KEYINPUT10), .Z(n350) );
  XNOR2_X1 U402 ( .A(G162GAT), .B(G106GAT), .ZN(n349) );
  XNOR2_X1 U403 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U404 ( .A(G218GAT), .B(n351), .ZN(n352) );
  XNOR2_X1 U405 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U406 ( .A(KEYINPUT66), .B(KEYINPUT82), .Z(n355) );
  NAND2_X1 U407 ( .A1(G232GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U408 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U409 ( .A(n357), .B(n356), .ZN(n360) );
  XNOR2_X1 U410 ( .A(n358), .B(KEYINPUT67), .ZN(n359) );
  XNOR2_X1 U411 ( .A(n360), .B(n359), .ZN(n544) );
  XOR2_X1 U412 ( .A(G78GAT), .B(G155GAT), .Z(n362) );
  XNOR2_X1 U413 ( .A(G22GAT), .B(G183GAT), .ZN(n361) );
  XNOR2_X1 U414 ( .A(n362), .B(n361), .ZN(n377) );
  XOR2_X1 U415 ( .A(n363), .B(G71GAT), .Z(n366) );
  XNOR2_X1 U416 ( .A(n364), .B(G127GAT), .ZN(n365) );
  XNOR2_X1 U417 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U418 ( .A(KEYINPUT12), .B(KEYINPUT83), .Z(n368) );
  NAND2_X1 U419 ( .A1(G231GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U420 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U421 ( .A(n370), .B(n369), .Z(n375) );
  XOR2_X1 U422 ( .A(KEYINPUT14), .B(G64GAT), .Z(n372) );
  XNOR2_X1 U423 ( .A(G8GAT), .B(G211GAT), .ZN(n371) );
  XNOR2_X1 U424 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U425 ( .A(n373), .B(KEYINPUT15), .ZN(n374) );
  XNOR2_X1 U426 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U427 ( .A(n377), .B(n376), .ZN(n550) );
  INV_X1 U428 ( .A(n550), .ZN(n573) );
  NAND2_X1 U429 ( .A1(n544), .A2(n573), .ZN(n378) );
  XNOR2_X1 U430 ( .A(n380), .B(KEYINPUT47), .ZN(n382) );
  XNOR2_X1 U431 ( .A(n382), .B(n381), .ZN(n390) );
  XNOR2_X1 U432 ( .A(KEYINPUT73), .B(n565), .ZN(n546) );
  XNOR2_X1 U433 ( .A(KEYINPUT36), .B(KEYINPUT103), .ZN(n383) );
  XOR2_X1 U434 ( .A(n544), .B(n383), .Z(n576) );
  NOR2_X1 U435 ( .A1(n573), .A2(n576), .ZN(n384) );
  XNOR2_X1 U436 ( .A(KEYINPUT45), .B(n384), .ZN(n386) );
  NAND2_X1 U437 ( .A1(n386), .A2(n385), .ZN(n387) );
  NOR2_X1 U438 ( .A1(n546), .A2(n387), .ZN(n388) );
  XNOR2_X1 U439 ( .A(KEYINPUT114), .B(n388), .ZN(n389) );
  NOR2_X1 U440 ( .A1(n390), .A2(n389), .ZN(n391) );
  XNOR2_X1 U441 ( .A(KEYINPUT48), .B(n391), .ZN(n519) );
  XOR2_X1 U442 ( .A(KEYINPUT97), .B(G204GAT), .Z(n393) );
  XNOR2_X1 U443 ( .A(G36GAT), .B(G190GAT), .ZN(n392) );
  XNOR2_X1 U444 ( .A(n393), .B(n392), .ZN(n404) );
  XOR2_X1 U445 ( .A(n395), .B(n394), .Z(n397) );
  NAND2_X1 U446 ( .A1(G226GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U447 ( .A(n397), .B(n396), .ZN(n398) );
  XOR2_X1 U448 ( .A(n398), .B(KEYINPUT95), .Z(n402) );
  XOR2_X1 U449 ( .A(G211GAT), .B(KEYINPUT21), .Z(n400) );
  XNOR2_X1 U450 ( .A(G197GAT), .B(G218GAT), .ZN(n399) );
  XNOR2_X1 U451 ( .A(n400), .B(n399), .ZN(n439) );
  XNOR2_X1 U452 ( .A(n439), .B(KEYINPUT96), .ZN(n401) );
  XNOR2_X1 U453 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U454 ( .A(n404), .B(n403), .ZN(n406) );
  XOR2_X1 U455 ( .A(n406), .B(n405), .Z(n511) );
  INV_X1 U456 ( .A(n511), .ZN(n407) );
  NOR2_X1 U457 ( .A1(n519), .A2(n407), .ZN(n408) );
  XNOR2_X1 U458 ( .A(n408), .B(KEYINPUT54), .ZN(n430) );
  XOR2_X1 U459 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n410) );
  XNOR2_X1 U460 ( .A(KEYINPUT94), .B(G57GAT), .ZN(n409) );
  XNOR2_X1 U461 ( .A(n410), .B(n409), .ZN(n424) );
  XOR2_X1 U462 ( .A(G148GAT), .B(G120GAT), .Z(n412) );
  XNOR2_X1 U463 ( .A(G29GAT), .B(G141GAT), .ZN(n411) );
  XNOR2_X1 U464 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U465 ( .A(KEYINPUT93), .B(KEYINPUT6), .Z(n414) );
  XNOR2_X1 U466 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n413) );
  XNOR2_X1 U467 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U468 ( .A(n416), .B(n415), .Z(n422) );
  XOR2_X1 U469 ( .A(G85GAT), .B(G134GAT), .Z(n418) );
  NAND2_X1 U470 ( .A1(G225GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U471 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U472 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U473 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U474 ( .A(n424), .B(n423), .ZN(n429) );
  XOR2_X1 U475 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n426) );
  XNOR2_X1 U476 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n425) );
  XNOR2_X1 U477 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U478 ( .A(G162GAT), .B(KEYINPUT3), .Z(n427) );
  XOR2_X1 U479 ( .A(n428), .B(n427), .Z(n446) );
  XOR2_X1 U480 ( .A(n429), .B(n446), .Z(n463) );
  NAND2_X1 U481 ( .A1(n430), .A2(n463), .ZN(n431) );
  XNOR2_X1 U482 ( .A(n431), .B(KEYINPUT65), .ZN(n564) );
  XOR2_X1 U483 ( .A(KEYINPUT23), .B(KEYINPUT89), .Z(n433) );
  XNOR2_X1 U484 ( .A(KEYINPUT88), .B(KEYINPUT24), .ZN(n432) );
  XNOR2_X1 U485 ( .A(n433), .B(n432), .ZN(n438) );
  XOR2_X1 U486 ( .A(n434), .B(KEYINPUT22), .Z(n436) );
  NAND2_X1 U487 ( .A1(G228GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U488 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n438), .B(n437), .ZN(n444) );
  XOR2_X1 U490 ( .A(n439), .B(KEYINPUT92), .Z(n442) );
  XNOR2_X1 U491 ( .A(G50GAT), .B(n440), .ZN(n441) );
  XNOR2_X1 U492 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U493 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U494 ( .A(n446), .B(n445), .ZN(n458) );
  AND2_X1 U495 ( .A1(n564), .A2(n458), .ZN(n447) );
  XNOR2_X1 U496 ( .A(n447), .B(KEYINPUT55), .ZN(n553) );
  NOR2_X1 U497 ( .A1(n455), .A2(n553), .ZN(n560) );
  INV_X1 U498 ( .A(n537), .ZN(n524) );
  NAND2_X1 U499 ( .A1(n560), .A2(n524), .ZN(n451) );
  XOR2_X1 U500 ( .A(G176GAT), .B(KEYINPUT57), .Z(n449) );
  XOR2_X1 U501 ( .A(KEYINPUT56), .B(KEYINPUT121), .Z(n448) );
  NAND2_X1 U502 ( .A1(n546), .A2(n385), .ZN(n483) );
  INV_X1 U503 ( .A(n544), .ZN(n559) );
  NOR2_X1 U504 ( .A1(n559), .A2(n573), .ZN(n452) );
  XNOR2_X1 U505 ( .A(KEYINPUT16), .B(n452), .ZN(n468) );
  XOR2_X1 U506 ( .A(KEYINPUT68), .B(KEYINPUT28), .Z(n453) );
  XNOR2_X1 U507 ( .A(n458), .B(n453), .ZN(n522) );
  INV_X1 U508 ( .A(n463), .ZN(n509) );
  XNOR2_X1 U509 ( .A(KEYINPUT27), .B(n511), .ZN(n460) );
  NAND2_X1 U510 ( .A1(n509), .A2(n460), .ZN(n518) );
  NOR2_X1 U511 ( .A1(n522), .A2(n518), .ZN(n454) );
  NAND2_X1 U512 ( .A1(n455), .A2(n454), .ZN(n466) );
  NAND2_X1 U513 ( .A1(n511), .A2(n551), .ZN(n456) );
  NAND2_X1 U514 ( .A1(n458), .A2(n456), .ZN(n457) );
  XOR2_X1 U515 ( .A(KEYINPUT25), .B(n457), .Z(n462) );
  NOR2_X1 U516 ( .A1(n458), .A2(n551), .ZN(n459) );
  XNOR2_X1 U517 ( .A(n459), .B(KEYINPUT26), .ZN(n563) );
  NAND2_X1 U518 ( .A1(n563), .A2(n460), .ZN(n461) );
  NAND2_X1 U519 ( .A1(n462), .A2(n461), .ZN(n464) );
  NAND2_X1 U520 ( .A1(n464), .A2(n463), .ZN(n465) );
  NAND2_X1 U521 ( .A1(n466), .A2(n465), .ZN(n467) );
  XNOR2_X1 U522 ( .A(KEYINPUT98), .B(n467), .ZN(n480) );
  NAND2_X1 U523 ( .A1(n468), .A2(n480), .ZN(n495) );
  NOR2_X1 U524 ( .A1(n483), .A2(n495), .ZN(n469) );
  XOR2_X1 U525 ( .A(KEYINPUT99), .B(n469), .Z(n478) );
  NAND2_X1 U526 ( .A1(n478), .A2(n509), .ZN(n470) );
  XNOR2_X1 U527 ( .A(n470), .B(KEYINPUT34), .ZN(n471) );
  XNOR2_X1 U528 ( .A(G1GAT), .B(n471), .ZN(G1324GAT) );
  NAND2_X1 U529 ( .A1(n478), .A2(n511), .ZN(n472) );
  XNOR2_X1 U530 ( .A(n472), .B(KEYINPUT100), .ZN(n473) );
  XNOR2_X1 U531 ( .A(G8GAT), .B(n473), .ZN(G1325GAT) );
  XOR2_X1 U532 ( .A(KEYINPUT35), .B(KEYINPUT102), .Z(n475) );
  NAND2_X1 U533 ( .A1(n478), .A2(n551), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n475), .B(n474), .ZN(n477) );
  XOR2_X1 U535 ( .A(G15GAT), .B(KEYINPUT101), .Z(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(G1326GAT) );
  NAND2_X1 U537 ( .A1(n478), .A2(n522), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n479), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n487) );
  NAND2_X1 U540 ( .A1(n573), .A2(n480), .ZN(n481) );
  NOR2_X1 U541 ( .A1(n576), .A2(n481), .ZN(n482) );
  XNOR2_X1 U542 ( .A(KEYINPUT37), .B(n482), .ZN(n508) );
  NOR2_X1 U543 ( .A1(n508), .A2(n483), .ZN(n485) );
  XNOR2_X1 U544 ( .A(KEYINPUT104), .B(KEYINPUT38), .ZN(n484) );
  XNOR2_X1 U545 ( .A(n485), .B(n484), .ZN(n492) );
  NAND2_X1 U546 ( .A1(n492), .A2(n509), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U548 ( .A(G29GAT), .B(n488), .Z(G1328GAT) );
  NAND2_X1 U549 ( .A1(n492), .A2(n511), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n489), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U551 ( .A1(n551), .A2(n492), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n490), .B(KEYINPUT40), .ZN(n491) );
  XNOR2_X1 U553 ( .A(G43GAT), .B(n491), .ZN(G1330GAT) );
  NAND2_X1 U554 ( .A1(n492), .A2(n522), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n493), .B(KEYINPUT106), .ZN(n494) );
  XNOR2_X1 U556 ( .A(G50GAT), .B(n494), .ZN(G1331GAT) );
  XNOR2_X1 U557 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n497) );
  NAND2_X1 U558 ( .A1(n524), .A2(n565), .ZN(n507) );
  NOR2_X1 U559 ( .A1(n495), .A2(n507), .ZN(n503) );
  NAND2_X1 U560 ( .A1(n509), .A2(n503), .ZN(n496) );
  XNOR2_X1 U561 ( .A(n497), .B(n496), .ZN(G1332GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n499) );
  NAND2_X1 U563 ( .A1(n503), .A2(n511), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U565 ( .A(G64GAT), .B(n500), .ZN(G1333GAT) );
  XOR2_X1 U566 ( .A(G71GAT), .B(KEYINPUT109), .Z(n502) );
  NAND2_X1 U567 ( .A1(n503), .A2(n551), .ZN(n501) );
  XNOR2_X1 U568 ( .A(n502), .B(n501), .ZN(G1334GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT43), .B(KEYINPUT110), .Z(n505) );
  NAND2_X1 U570 ( .A1(n503), .A2(n522), .ZN(n504) );
  XNOR2_X1 U571 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U572 ( .A(G78GAT), .B(n506), .ZN(G1335GAT) );
  NOR2_X1 U573 ( .A1(n508), .A2(n507), .ZN(n514) );
  NAND2_X1 U574 ( .A1(n509), .A2(n514), .ZN(n510) );
  XNOR2_X1 U575 ( .A(G85GAT), .B(n510), .ZN(G1336GAT) );
  NAND2_X1 U576 ( .A1(n514), .A2(n511), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n512), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U578 ( .A1(n551), .A2(n514), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n513), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n516) );
  NAND2_X1 U581 ( .A1(n514), .A2(n522), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U583 ( .A(G106GAT), .B(n517), .ZN(G1339GAT) );
  NOR2_X1 U584 ( .A1(n519), .A2(n518), .ZN(n535) );
  NAND2_X1 U585 ( .A1(n535), .A2(n551), .ZN(n520) );
  XOR2_X1 U586 ( .A(KEYINPUT115), .B(n520), .Z(n521) );
  NOR2_X1 U587 ( .A1(n522), .A2(n521), .ZN(n531) );
  NAND2_X1 U588 ( .A1(n531), .A2(n546), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n523), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n526) );
  NAND2_X1 U591 ( .A1(n531), .A2(n524), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n526), .B(n525), .ZN(n528) );
  XOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT116), .Z(n527) );
  XNOR2_X1 U594 ( .A(n528), .B(n527), .ZN(G1341GAT) );
  NAND2_X1 U595 ( .A1(n550), .A2(n531), .ZN(n529) );
  XNOR2_X1 U596 ( .A(n529), .B(KEYINPUT50), .ZN(n530) );
  XNOR2_X1 U597 ( .A(G127GAT), .B(n530), .ZN(G1342GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT51), .B(KEYINPUT118), .Z(n533) );
  NAND2_X1 U599 ( .A1(n531), .A2(n559), .ZN(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U601 ( .A(G134GAT), .B(n534), .ZN(G1343GAT) );
  NAND2_X1 U602 ( .A1(n535), .A2(n563), .ZN(n543) );
  NOR2_X1 U603 ( .A1(n565), .A2(n543), .ZN(n536) );
  XOR2_X1 U604 ( .A(G141GAT), .B(n536), .Z(G1344GAT) );
  NOR2_X1 U605 ( .A1(n537), .A2(n543), .ZN(n539) );
  XNOR2_X1 U606 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(n540), .ZN(G1345GAT) );
  NOR2_X1 U609 ( .A1(n573), .A2(n543), .ZN(n542) );
  XNOR2_X1 U610 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n541) );
  XNOR2_X1 U611 ( .A(n542), .B(n541), .ZN(G1346GAT) );
  NOR2_X1 U612 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U613 ( .A(G162GAT), .B(n545), .Z(G1347GAT) );
  NAND2_X1 U614 ( .A1(n551), .A2(n546), .ZN(n547) );
  OR2_X1 U615 ( .A1(n553), .A2(n547), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n548), .B(KEYINPUT120), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n549), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  OR2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n554), .B(KEYINPUT122), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n557) );
  XNOR2_X1 U623 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U625 ( .A(KEYINPUT123), .B(n558), .Z(n562) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1351GAT) );
  NAND2_X1 U628 ( .A1(n564), .A2(n563), .ZN(n575) );
  NOR2_X1 U629 ( .A1(n565), .A2(n575), .ZN(n570) );
  XOR2_X1 U630 ( .A(KEYINPUT127), .B(KEYINPUT60), .Z(n567) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(KEYINPUT126), .B(n568), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  NOR2_X1 U635 ( .A1(n385), .A2(n575), .ZN(n572) );
  XNOR2_X1 U636 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1353GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n575), .ZN(n574) );
  XOR2_X1 U639 ( .A(G211GAT), .B(n574), .Z(G1354GAT) );
  NOR2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT62), .B(n577), .Z(n578) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(n578), .ZN(G1355GAT) );
endmodule

