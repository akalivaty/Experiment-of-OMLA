//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 1 1 0 1 1 0 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035;
  INV_X1    g000(.A(KEYINPUT81), .ZN(new_n187));
  XOR2_X1   g001(.A(G110), .B(G140), .Z(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT76), .ZN(new_n189));
  INV_X1    g003(.A(G227), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G953), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n189), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT77), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n193), .A2(KEYINPUT77), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G104), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n194), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G101), .ZN(new_n199));
  INV_X1    g013(.A(G104), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G107), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n193), .A2(new_n196), .A3(KEYINPUT77), .A4(G104), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n198), .A2(new_n199), .A3(new_n201), .A4(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n197), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G101), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT79), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT65), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n209), .A2(new_n211), .A3(G143), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n208), .A2(G143), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G128), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n212), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n215), .B1(new_n212), .B2(KEYINPUT1), .ZN(new_n218));
  INV_X1    g032(.A(G143), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n209), .A2(new_n211), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(new_n219), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n217), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT79), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n203), .A2(new_n224), .A3(new_n205), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n207), .A2(KEYINPUT10), .A3(new_n223), .A4(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G137), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT11), .A3(G134), .ZN(new_n228));
  INV_X1    g042(.A(G134), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G137), .ZN(new_n230));
  AOI21_X1  g044(.A(KEYINPUT11), .B1(new_n227), .B2(G134), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n228), .B(new_n230), .C1(new_n231), .C2(KEYINPUT66), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n227), .A2(G134), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT11), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(KEYINPUT66), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(G131), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n228), .A2(new_n230), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n229), .A2(G137), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(KEYINPUT11), .ZN(new_n241));
  INV_X1    g055(.A(G131), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n238), .A2(new_n241), .A3(new_n242), .A4(new_n235), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n237), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT77), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n200), .A2(G107), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n202), .A2(new_n201), .ZN(new_n251));
  OAI21_X1  g065(.A(G101), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(KEYINPUT4), .A3(new_n203), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n210), .A2(G146), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n208), .A2(KEYINPUT65), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n219), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n220), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  NOR2_X1   g073(.A1(KEYINPUT0), .A2(G128), .ZN(new_n260));
  OR2_X1    g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT65), .B(G146), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n213), .B1(new_n263), .B2(G143), .ZN(new_n264));
  AOI22_X1  g078(.A1(new_n258), .A2(new_n262), .B1(new_n264), .B2(new_n259), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n266), .B(G101), .C1(new_n250), .C2(new_n251), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n253), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n212), .A2(new_n214), .A3(new_n216), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT1), .B1(new_n219), .B2(G146), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n212), .A2(new_n214), .B1(G128), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n269), .B1(new_n273), .B2(new_n206), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n226), .A2(new_n245), .A3(new_n268), .A4(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n223), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n203), .A2(new_n224), .A3(new_n205), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n224), .B1(new_n203), .B2(new_n205), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OR2_X1    g093(.A1(new_n273), .A2(new_n206), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n245), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT12), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n275), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  AOI211_X1 g097(.A(KEYINPUT12), .B(new_n245), .C1(new_n279), .C2(new_n280), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n192), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n226), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n268), .A2(new_n274), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n244), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n192), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n275), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT80), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT80), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n285), .A2(new_n293), .A3(new_n290), .ZN(new_n294));
  AOI21_X1  g108(.A(G902), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G469), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n187), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n285), .A2(new_n293), .A3(new_n290), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n293), .B1(new_n285), .B2(new_n290), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(KEYINPUT81), .A3(G469), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n223), .B1(new_n207), .B2(new_n225), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n273), .A2(new_n206), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n244), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(KEYINPUT12), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n281), .A2(new_n282), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n306), .A2(new_n307), .A3(new_n275), .A4(new_n289), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n268), .A2(new_n274), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n245), .B1(new_n309), .B2(new_n226), .ZN(new_n310));
  INV_X1    g124(.A(new_n275), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n192), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(G902), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n296), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n297), .A2(new_n302), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT72), .ZN(new_n316));
  INV_X1    g130(.A(G125), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(G140), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(G140), .ZN(new_n319));
  INV_X1    g133(.A(G140), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(KEYINPUT72), .A3(G125), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n318), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n322), .A2(KEYINPUT16), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT16), .B1(new_n320), .B2(G125), .ZN(new_n324));
  OAI21_X1  g138(.A(G146), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT88), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n324), .B1(new_n322), .B2(KEYINPUT16), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n208), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n325), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n327), .A2(new_n208), .ZN(new_n330));
  AOI211_X1 g144(.A(G146), .B(new_n324), .C1(new_n322), .C2(KEYINPUT16), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT88), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(G237), .A2(G953), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(G214), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n219), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n333), .A2(G143), .A3(G214), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G131), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT17), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n335), .A2(new_n242), .A3(new_n336), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n337), .A2(KEYINPUT17), .A3(G131), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n329), .A2(new_n332), .A3(new_n341), .A4(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(G113), .B(G122), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(new_n200), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n337), .A2(KEYINPUT18), .A3(G131), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n322), .A2(G146), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n320), .A2(G125), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n263), .A2(new_n348), .A3(new_n319), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(KEYINPUT18), .A2(G131), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n335), .A2(new_n336), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n346), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n343), .A2(new_n345), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n322), .A2(KEYINPUT19), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT19), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n348), .A2(new_n319), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n355), .A2(new_n263), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT86), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n338), .A2(new_n340), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT86), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n355), .A2(new_n361), .A3(new_n263), .A4(new_n357), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n359), .A2(new_n325), .A3(new_n360), .A4(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(KEYINPUT87), .A3(new_n353), .ZN(new_n364));
  INV_X1    g178(.A(new_n345), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT87), .B1(new_n363), .B2(new_n353), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n354), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT89), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(G475), .A2(G902), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n354), .B(KEYINPUT89), .C1(new_n366), .C2(new_n367), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NOR3_X1   g187(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n373), .A2(KEYINPUT20), .B1(new_n368), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n345), .B1(new_n343), .B2(new_n353), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(G902), .B1(new_n377), .B2(new_n354), .ZN(new_n378));
  INV_X1    g192(.A(G475), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G122), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G116), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n196), .B1(new_n383), .B2(KEYINPUT14), .ZN(new_n384));
  XNOR2_X1  g198(.A(G116), .B(G122), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n384), .B(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n219), .A2(G128), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n215), .A2(G143), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n389), .A2(KEYINPUT90), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT90), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n391), .B1(new_n387), .B2(new_n388), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n390), .A2(new_n229), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n389), .A2(KEYINPUT90), .ZN(new_n394));
  XNOR2_X1  g208(.A(G128), .B(G143), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n391), .ZN(new_n396));
  AOI21_X1  g210(.A(G134), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n386), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n229), .B1(new_n390), .B2(new_n392), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(KEYINPUT13), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n400), .B(G134), .C1(KEYINPUT13), .C2(new_n387), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n385), .B(new_n196), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(KEYINPUT9), .B(G234), .ZN(new_n404));
  INV_X1    g218(.A(G217), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n404), .A2(new_n405), .A3(G953), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n398), .A2(new_n403), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n406), .B1(new_n398), .B2(new_n403), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n298), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT91), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n398), .A2(new_n403), .ZN(new_n412));
  INV_X1    g226(.A(new_n406), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n398), .A2(new_n403), .A3(new_n406), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT91), .A3(new_n298), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT15), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G478), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n409), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n420), .B1(new_n422), .B2(KEYINPUT91), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(G952), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(G953), .ZN(new_n427));
  INV_X1    g241(.A(G234), .ZN(new_n428));
  INV_X1    g242(.A(G237), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n427), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  OAI211_X1 g245(.A(G902), .B(G953), .C1(new_n428), .C2(new_n429), .ZN(new_n432));
  XOR2_X1   g246(.A(new_n432), .B(KEYINPUT92), .Z(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(G898), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n425), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n381), .A2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G210), .B1(G237), .B2(G902), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(G110), .B(G122), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(G116), .B(G119), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT5), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT5), .ZN(new_n445));
  INV_X1    g259(.A(G119), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n446), .A3(G116), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT82), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n445), .A2(new_n446), .A3(KEYINPUT82), .A4(G116), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n444), .A2(G113), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  XOR2_X1   g265(.A(G116), .B(G119), .Z(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT2), .B(G113), .ZN(new_n453));
  OR2_X1    g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n451), .A2(new_n454), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n277), .A2(new_n278), .A3(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n452), .B(new_n453), .ZN(new_n457));
  AND3_X1   g271(.A1(new_n253), .A2(new_n267), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n442), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n451), .A2(new_n454), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n207), .A2(new_n460), .A3(new_n225), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n253), .A2(new_n267), .A3(new_n457), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n441), .A3(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n459), .A2(KEYINPUT6), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n465), .B(new_n442), .C1(new_n456), .C2(new_n458), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n261), .B1(new_n256), .B2(new_n257), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n212), .A2(new_n214), .A3(new_n259), .ZN(new_n468));
  OAI21_X1  g282(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n317), .B(new_n217), .C1(new_n218), .C2(new_n222), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G953), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G224), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT83), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n471), .B(new_n474), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n464), .A2(new_n466), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n455), .A2(new_n206), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n461), .A2(new_n477), .ZN(new_n478));
  XOR2_X1   g292(.A(new_n441), .B(KEYINPUT8), .Z(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT7), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n474), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n469), .B(new_n470), .C1(KEYINPUT84), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n469), .A2(KEYINPUT84), .ZN(new_n485));
  INV_X1    g299(.A(new_n483), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n471), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n481), .A2(new_n463), .A3(new_n484), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n298), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n440), .B1(new_n476), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n487), .A2(new_n484), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n479), .B1(new_n461), .B2(new_n477), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(G902), .B1(new_n493), .B2(new_n463), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n464), .A2(new_n466), .A3(new_n475), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(new_n439), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(G214), .B1(G237), .B2(G902), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(KEYINPUT85), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT85), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n497), .A2(new_n502), .A3(new_n499), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(G221), .B1(new_n404), .B2(G902), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(KEYINPUT75), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n315), .A2(new_n438), .A3(new_n504), .A4(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n405), .B1(G234), .B2(new_n298), .ZN(new_n509));
  XNOR2_X1  g323(.A(KEYINPUT22), .B(G137), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n472), .A2(G221), .A3(G234), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT23), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n513), .B1(new_n446), .B2(G128), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n215), .A2(KEYINPUT23), .A3(G119), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n514), .B(new_n515), .C1(G119), .C2(new_n215), .ZN(new_n516));
  XNOR2_X1  g330(.A(G119), .B(G128), .ZN(new_n517));
  XOR2_X1   g331(.A(KEYINPUT24), .B(G110), .Z(new_n518));
  OAI22_X1  g332(.A1(new_n516), .A2(G110), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n325), .A2(new_n349), .A3(new_n519), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n516), .A2(G110), .B1(new_n517), .B2(new_n518), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n521), .B1(new_n330), .B2(new_n331), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT73), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g338(.A(KEYINPUT73), .B(new_n521), .C1(new_n330), .C2(new_n331), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n520), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n512), .B1(new_n526), .B2(KEYINPUT74), .ZN(new_n527));
  INV_X1    g341(.A(new_n520), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n325), .A2(new_n328), .ZN(new_n529));
  AOI21_X1  g343(.A(KEYINPUT73), .B1(new_n529), .B2(new_n521), .ZN(new_n530));
  INV_X1    g344(.A(new_n525), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT74), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n527), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n532), .A2(new_n533), .A3(new_n512), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT25), .B1(new_n537), .B2(new_n298), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT25), .ZN(new_n539));
  AOI211_X1 g353(.A(new_n539), .B(G902), .C1(new_n535), .C2(new_n536), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n509), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n509), .A2(G902), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT32), .ZN(new_n545));
  XOR2_X1   g359(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n546));
  NAND2_X1  g360(.A1(new_n333), .A2(G210), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(KEYINPUT26), .B(G101), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n548), .B(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT67), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n230), .B1(new_n240), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n233), .A2(KEYINPUT67), .ZN(new_n553));
  OAI21_X1  g367(.A(G131), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n223), .A2(new_n243), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n212), .A2(new_n214), .A3(new_n259), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n556), .B1(new_n222), .B2(new_n261), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n557), .B1(new_n237), .B2(new_n243), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n457), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n244), .A2(new_n265), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n223), .A2(new_n243), .A3(new_n554), .ZN(new_n561));
  INV_X1    g375(.A(new_n457), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT28), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n243), .A2(new_n554), .ZN(new_n566));
  AOI22_X1  g380(.A1(new_n566), .A2(new_n223), .B1(new_n244), .B2(new_n265), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT28), .B1(new_n567), .B2(new_n562), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n550), .B1(new_n565), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT31), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT68), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n572), .B1(new_n567), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n573), .ZN(new_n575));
  OAI211_X1 g389(.A(KEYINPUT68), .B(new_n575), .C1(new_n555), .C2(new_n558), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n567), .A2(KEYINPUT30), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n574), .A2(new_n457), .A3(new_n576), .A4(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n563), .ZN(new_n579));
  INV_X1    g393(.A(new_n550), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n571), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n578), .A2(new_n571), .A3(new_n581), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(KEYINPUT70), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT70), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n578), .A2(new_n585), .A3(new_n571), .A4(new_n581), .ZN(new_n586));
  AOI211_X1 g400(.A(new_n570), .B(new_n582), .C1(new_n584), .C2(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(G472), .A2(G902), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n545), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n565), .A2(KEYINPUT29), .A3(new_n550), .A4(new_n569), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT71), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n568), .B1(new_n564), .B2(KEYINPUT28), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT71), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n593), .A2(new_n594), .A3(KEYINPUT29), .A4(new_n550), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n550), .B1(new_n578), .B2(new_n563), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT29), .B1(new_n593), .B2(new_n550), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n596), .A2(new_n600), .A3(new_n298), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n584), .A2(new_n586), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n582), .A2(new_n570), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n589), .A2(new_n545), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n601), .A2(G472), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n544), .B1(new_n590), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n508), .A2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(new_n199), .ZN(G3));
  AOI21_X1  g424(.A(G902), .B1(new_n602), .B2(new_n603), .ZN(new_n611));
  INV_X1    g425(.A(G472), .ZN(new_n612));
  OAI22_X1  g426(.A1(new_n611), .A2(new_n612), .B1(new_n587), .B2(new_n589), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(new_n544), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(new_n507), .A3(new_n315), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n298), .A2(G478), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n416), .A2(KEYINPUT33), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT33), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n414), .A2(new_n618), .A3(new_n415), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n616), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(KEYINPUT94), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT94), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n622), .B1(new_n422), .B2(G478), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n621), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n625), .B1(new_n375), .B2(new_n380), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT95), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT95), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n625), .B(new_n628), .C1(new_n375), .C2(new_n380), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT93), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n490), .A2(new_n631), .A3(new_n496), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n439), .B1(new_n494), .B2(new_n495), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n500), .B1(new_n633), .B2(KEYINPUT93), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n635), .A2(new_n435), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n630), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n615), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT34), .B(G104), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  AND3_X1   g454(.A1(new_n614), .A2(new_n507), .A3(new_n315), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n373), .A2(KEYINPUT20), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT20), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n370), .A2(new_n643), .A3(new_n371), .A4(new_n372), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  AOI22_X1  g459(.A1(new_n411), .A2(new_n417), .B1(new_n419), .B2(G478), .ZN(new_n646));
  OAI22_X1  g460(.A1(new_n646), .A2(new_n423), .B1(new_n378), .B2(new_n379), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n649), .A2(new_n635), .A3(new_n435), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n641), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  INV_X1    g467(.A(KEYINPUT96), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT36), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n512), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n526), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n542), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n541), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n589), .B1(new_n602), .B2(new_n603), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g475(.A(G472), .B1(new_n587), .B2(G902), .ZN(new_n662));
  AND4_X1   g476(.A1(new_n654), .A2(new_n659), .A3(new_n661), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n604), .A2(new_n298), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n660), .B1(new_n664), .B2(G472), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n654), .B1(new_n665), .B2(new_n659), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n667), .A2(new_n508), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT37), .B(G110), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT97), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n668), .B(new_n670), .ZN(G12));
  AND2_X1   g485(.A1(new_n302), .A2(new_n314), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n506), .B1(new_n672), .B2(new_n297), .ZN(new_n673));
  INV_X1    g487(.A(G900), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n431), .B1(new_n433), .B2(new_n674), .ZN(new_n675));
  AOI211_X1 g489(.A(new_n675), .B(new_n647), .C1(new_n642), .C2(new_n644), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT98), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n632), .A2(new_n634), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n675), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n645), .A2(new_n648), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g495(.A(KEYINPUT98), .B1(new_n681), .B2(new_n635), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  AOI22_X1  g497(.A1(new_n606), .A2(new_n590), .B1(new_n541), .B2(new_n658), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n673), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G128), .ZN(G30));
  XOR2_X1   g500(.A(new_n675), .B(KEYINPUT39), .Z(new_n687));
  NAND2_X1  g501(.A1(new_n673), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(KEYINPUT40), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n604), .A2(new_n605), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n578), .A2(new_n581), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n612), .B1(new_n564), .B2(new_n580), .ZN(new_n693));
  AOI22_X1  g507(.A1(new_n692), .A2(new_n693), .B1(G472), .B2(G902), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT99), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(new_n696));
  OAI211_X1 g510(.A(new_n691), .B(new_n696), .C1(KEYINPUT32), .C2(new_n660), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT38), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n497), .B(new_n698), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n425), .B1(new_n375), .B2(new_n380), .ZN(new_n700));
  NOR4_X1   g514(.A1(new_n699), .A2(new_n659), .A3(new_n700), .A4(new_n500), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n689), .A2(new_n690), .A3(new_n697), .A4(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G143), .ZN(G45));
  INV_X1    g517(.A(KEYINPUT100), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n625), .B(new_n680), .C1(new_n375), .C2(new_n380), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n704), .B1(new_n705), .B2(new_n635), .ZN(new_n706));
  INV_X1    g520(.A(new_n705), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(KEYINPUT100), .A3(new_n678), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n673), .A2(new_n684), .A3(new_n706), .A4(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  AND2_X1   g524(.A1(new_n592), .A2(new_n595), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n565), .A2(new_n550), .A3(new_n569), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT29), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n298), .B1(new_n714), .B2(new_n597), .ZN(new_n715));
  OAI21_X1  g529(.A(G472), .B1(new_n711), .B2(new_n715), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n716), .B(new_n691), .C1(KEYINPUT32), .C2(new_n660), .ZN(new_n717));
  INV_X1    g531(.A(new_n544), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT101), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n313), .B2(new_n296), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n283), .A2(new_n284), .A3(new_n192), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n289), .B1(new_n288), .B2(new_n275), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n298), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(G469), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n723), .A2(new_n719), .A3(G469), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n506), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n717), .A2(new_n718), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n637), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g543(.A(KEYINPUT41), .B(G113), .Z(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G15));
  NAND4_X1  g545(.A1(new_n650), .A2(new_n717), .A3(new_n718), .A4(new_n727), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G116), .ZN(G18));
  NAND2_X1  g547(.A1(new_n725), .A2(new_n726), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n734), .A2(new_n678), .A3(new_n507), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n684), .A2(new_n735), .A3(new_n438), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G119), .ZN(G21));
  NOR2_X1   g551(.A1(new_n700), .A2(new_n635), .ZN(new_n738));
  AOI211_X1 g552(.A(new_n506), .B(new_n435), .C1(new_n725), .C2(new_n726), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n614), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  XOR2_X1   g554(.A(KEYINPUT102), .B(G122), .Z(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G24));
  NAND2_X1  g556(.A1(new_n665), .A2(new_n659), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n727), .A2(new_n678), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n743), .A2(new_n744), .A3(new_n705), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n317), .ZN(G27));
  INV_X1    g560(.A(KEYINPUT42), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n490), .A2(new_n499), .A3(new_n496), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT104), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n290), .A2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n288), .A2(KEYINPUT104), .A3(new_n275), .A4(new_n289), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n750), .A2(new_n285), .A3(G469), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(G469), .A2(G902), .ZN(new_n753));
  XOR2_X1   g567(.A(new_n753), .B(KEYINPUT103), .Z(new_n754));
  NAND3_X1  g568(.A1(new_n314), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n748), .A2(new_n755), .A3(new_n507), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n717), .A2(new_n718), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n747), .B1(new_n757), .B2(new_n705), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n607), .A2(KEYINPUT42), .A3(new_n707), .A4(new_n756), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(new_n242), .ZN(G33));
  INV_X1    g575(.A(KEYINPUT105), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n681), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n645), .A2(KEYINPUT105), .A3(new_n648), .A4(new_n680), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n757), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(KEYINPUT106), .B(G134), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(G36));
  NAND2_X1  g582(.A1(new_n381), .A2(new_n625), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT43), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n658), .ZN(new_n772));
  AOI21_X1  g586(.A(G902), .B1(new_n535), .B2(new_n536), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT25), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n772), .B1(new_n774), .B2(new_n509), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n665), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n771), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n771), .A2(KEYINPUT44), .A3(new_n776), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(new_n748), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT45), .B1(new_n292), .B2(new_n294), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n750), .A2(new_n285), .A3(KEYINPUT45), .A4(new_n751), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(G469), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(KEYINPUT46), .A3(new_n754), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT107), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n785), .A2(KEYINPUT107), .A3(KEYINPUT46), .A4(new_n754), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT46), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n782), .A2(new_n784), .ZN(new_n791));
  INV_X1    g605(.A(new_n754), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n788), .A2(new_n314), .A3(new_n789), .A4(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n507), .A3(new_n687), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n781), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(KEYINPUT108), .B(G137), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n796), .B(new_n797), .ZN(G39));
  NAND2_X1  g612(.A1(new_n794), .A2(new_n507), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT47), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n794), .A2(KEYINPUT47), .A3(new_n507), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n748), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n717), .A2(new_n718), .A3(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n803), .A2(new_n707), .A3(new_n805), .ZN(new_n806));
  XOR2_X1   g620(.A(KEYINPUT109), .B(G140), .Z(new_n807));
  XNOR2_X1  g621(.A(new_n806), .B(new_n807), .ZN(G42));
  XOR2_X1   g622(.A(new_n734), .B(KEYINPUT49), .Z(new_n809));
  NAND4_X1  g623(.A1(new_n718), .A2(new_n507), .A3(new_n699), .A4(new_n499), .ZN(new_n810));
  OR4_X1    g624(.A1(new_n697), .A2(new_n809), .A3(new_n769), .A4(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n743), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(new_n707), .A3(new_n735), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n709), .A2(new_n685), .A3(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n541), .A2(new_n658), .A3(new_n680), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n755), .A2(new_n507), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n738), .A2(new_n815), .A3(new_n697), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT114), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n659), .A2(new_n816), .A3(new_n675), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT114), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(new_n821), .A3(new_n697), .A4(new_n738), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT52), .B1(new_n814), .B2(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n315), .A2(new_n507), .A3(new_n717), .A4(new_n659), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n745), .B1(new_n826), .B2(new_n683), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n819), .A2(new_n822), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n827), .A2(new_n828), .A3(new_n709), .A4(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n824), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n508), .B1(new_n667), .B2(new_n608), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n435), .B1(new_n501), .B2(new_n503), .ZN(new_n833));
  INV_X1    g647(.A(new_n375), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT110), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(new_n835), .A3(new_n648), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT110), .B1(new_n375), .B2(new_n647), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n836), .A2(new_n626), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n833), .A2(new_n838), .ZN(new_n839));
  OAI22_X1  g653(.A1(new_n615), .A2(new_n839), .B1(new_n637), .B2(new_n728), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n736), .A2(new_n732), .A3(new_n740), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n832), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n354), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n298), .B1(new_n843), .B2(new_n376), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(G475), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n421), .A3(new_n424), .A4(new_n680), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n645), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n804), .B1(new_n848), .B2(KEYINPUT111), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(KEYINPUT111), .B2(new_n848), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT112), .B1(new_n825), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n846), .B1(new_n642), .B2(new_n644), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT111), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n748), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n848), .A2(KEYINPUT111), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT112), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n673), .A2(new_n856), .A3(new_n857), .A4(new_n684), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n851), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n707), .A2(new_n665), .A3(new_n756), .A4(new_n659), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n860), .B1(new_n757), .B2(new_n765), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n759), .B2(new_n758), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n842), .A2(KEYINPUT113), .A3(new_n859), .A4(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT113), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n859), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n833), .A2(new_n838), .ZN(new_n866));
  AOI211_X1 g680(.A(new_n435), .B(new_n635), .C1(new_n627), .C2(new_n629), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n717), .A2(new_n718), .A3(new_n727), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n641), .A2(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n736), .A2(new_n732), .A3(new_n740), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n437), .B1(new_n503), .B2(new_n501), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT96), .B1(new_n775), .B2(new_n613), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n665), .A2(new_n654), .A3(new_n659), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n673), .B(new_n871), .C1(new_n874), .C2(new_n607), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n869), .A2(new_n870), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n864), .B1(new_n865), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n831), .B1(new_n863), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT53), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n863), .A2(new_n877), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n879), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n824), .A2(KEYINPUT115), .A3(new_n830), .ZN(new_n882));
  AOI21_X1  g696(.A(KEYINPUT115), .B1(new_n824), .B2(new_n830), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI221_X1 g698(.A(KEYINPUT54), .B1(new_n878), .B2(new_n879), .C1(new_n881), .C2(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n842), .A2(KEYINPUT53), .A3(new_n859), .A4(new_n862), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n887), .B1(new_n882), .B2(new_n883), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT54), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n888), .B(new_n889), .C1(KEYINPUT53), .C2(new_n878), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n771), .A2(new_n431), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AND3_X1   g706(.A1(new_n699), .A2(new_n727), .A3(new_n500), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n892), .A2(new_n614), .A3(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT117), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n895), .A3(KEYINPUT50), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n727), .A2(new_n748), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  NOR4_X1   g712(.A1(new_n897), .A2(new_n697), .A3(new_n430), .A4(new_n544), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n375), .A2(new_n625), .A3(new_n380), .ZN(new_n900));
  AOI22_X1  g714(.A1(new_n898), .A2(new_n812), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT50), .B1(new_n894), .B2(new_n895), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT118), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(new_n903), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT118), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n905), .A2(new_n906), .A3(new_n896), .A4(new_n901), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n734), .A2(new_n506), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n801), .A2(new_n802), .A3(new_n908), .ZN(new_n909));
  NOR4_X1   g723(.A1(new_n891), .A2(new_n544), .A3(new_n613), .A4(new_n804), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n904), .A2(new_n907), .A3(KEYINPUT51), .A4(new_n911), .ZN(new_n912));
  XNOR2_X1  g726(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n905), .A2(new_n896), .A3(new_n901), .ZN(new_n914));
  INV_X1    g728(.A(new_n911), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n892), .A2(new_n614), .A3(new_n735), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n899), .A2(new_n630), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n917), .A2(new_n427), .A3(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT119), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n898), .A2(new_n607), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT48), .ZN(new_n924));
  OR2_X1    g738(.A1(new_n923), .A2(KEYINPUT48), .ZN(new_n925));
  AOI22_X1  g739(.A1(new_n921), .A2(new_n922), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n916), .A2(new_n926), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n885), .A2(new_n890), .A3(new_n912), .A4(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT120), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n426), .A2(new_n472), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n928), .A2(new_n929), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n811), .B1(new_n932), .B2(new_n933), .ZN(G75));
  OAI21_X1  g748(.A(new_n888), .B1(KEYINPUT53), .B2(new_n878), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n935), .A2(G902), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(G210), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n464), .A2(new_n466), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(new_n475), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT55), .Z(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n942), .A2(KEYINPUT56), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n937), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n941), .B1(new_n937), .B2(new_n943), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n472), .A2(G952), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(G51));
  INV_X1    g761(.A(new_n831), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT53), .B1(new_n880), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT115), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n831), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n824), .A2(KEYINPUT115), .A3(new_n830), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n886), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(KEYINPUT54), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n890), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n754), .B(KEYINPUT57), .ZN(new_n957));
  OAI22_X1  g771(.A1(new_n956), .A2(new_n957), .B1(new_n722), .B2(new_n721), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n936), .A2(new_n791), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n946), .B1(new_n958), .B2(new_n959), .ZN(G54));
  NAND3_X1  g774(.A1(new_n936), .A2(KEYINPUT58), .A3(G475), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n370), .A2(new_n372), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n963), .A2(new_n964), .A3(new_n946), .ZN(G60));
  INV_X1    g779(.A(new_n946), .ZN(new_n966));
  INV_X1    g780(.A(new_n617), .ZN(new_n967));
  INV_X1    g781(.A(new_n619), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(G478), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT59), .Z(new_n971));
  NOR2_X1   g785(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(KEYINPUT122), .B1(new_n955), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT122), .ZN(new_n974));
  INV_X1    g788(.A(new_n972), .ZN(new_n975));
  AOI211_X1 g789(.A(new_n974), .B(new_n975), .C1(new_n954), .C2(new_n890), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n966), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n971), .B1(new_n885), .B2(new_n890), .ZN(new_n978));
  INV_X1    g792(.A(new_n969), .ZN(new_n979));
  OAI21_X1  g793(.A(KEYINPUT123), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OR3_X1    g794(.A1(new_n978), .A2(KEYINPUT123), .A3(new_n979), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n977), .B1(new_n980), .B2(new_n981), .ZN(G63));
  INV_X1    g796(.A(KEYINPUT61), .ZN(new_n983));
  NAND2_X1  g797(.A1(G217), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT60), .Z(new_n985));
  NAND3_X1  g799(.A1(new_n935), .A2(new_n657), .A3(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n983), .B1(new_n987), .B2(KEYINPUT124), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n986), .A2(new_n966), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n537), .B1(new_n935), .B2(new_n985), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n988), .B(new_n991), .ZN(G66));
  INV_X1    g806(.A(G224), .ZN(new_n993));
  OAI21_X1  g807(.A(G953), .B1(new_n434), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n994), .B1(new_n842), .B2(G953), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n938), .B1(G898), .B2(new_n472), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n995), .B(new_n996), .ZN(G69));
  NAND3_X1  g811(.A1(new_n574), .A2(new_n577), .A3(new_n576), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n355), .A2(new_n357), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT125), .Z(new_n1000));
  XNOR2_X1  g814(.A(new_n998), .B(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1001), .B1(new_n674), .B2(new_n472), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n806), .A2(new_n796), .ZN(new_n1003));
  NOR4_X1   g817(.A1(new_n795), .A2(new_n608), .A3(new_n635), .A4(new_n700), .ZN(new_n1004));
  NOR4_X1   g818(.A1(new_n1004), .A2(new_n760), .A3(new_n766), .A4(new_n814), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1002), .B1(new_n1007), .B2(new_n472), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n702), .A2(new_n709), .A3(new_n827), .ZN(new_n1009));
  OR2_X1    g823(.A1(new_n1009), .A2(KEYINPUT62), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n607), .A2(new_n748), .A3(new_n838), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n688), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1012), .B1(new_n1009), .B2(KEYINPUT62), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1010), .A2(new_n1003), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1001), .B1(new_n1014), .B2(new_n472), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n1008), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(G953), .B1(new_n190), .B2(new_n674), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1016), .B(new_n1017), .ZN(G72));
  NAND2_X1  g832(.A1(G472), .A2(G902), .ZN(new_n1019));
  XOR2_X1   g833(.A(new_n1019), .B(KEYINPUT63), .Z(new_n1020));
  OAI21_X1  g834(.A(new_n1020), .B1(new_n1006), .B2(new_n876), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n578), .A2(new_n563), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1022), .B(KEYINPUT126), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n1023), .A2(new_n550), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n946), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  OAI22_X1  g839(.A1(new_n881), .A2(new_n884), .B1(new_n878), .B2(new_n879), .ZN(new_n1026));
  INV_X1    g840(.A(new_n692), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1020), .B1(new_n1027), .B2(new_n597), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1025), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1023), .A2(new_n550), .ZN(new_n1030));
  OR2_X1    g844(.A1(new_n1014), .A2(new_n876), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1030), .B1(new_n1031), .B2(new_n1020), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT127), .ZN(new_n1033));
  OR2_X1    g847(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1029), .B1(new_n1034), .B2(new_n1035), .ZN(G57));
endmodule


