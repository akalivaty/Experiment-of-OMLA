//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1222, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  AND2_X1   g0006(.A1(G107), .A2(G264), .ZN(new_n207));
  INV_X1    g0007(.A(G87), .ZN(new_n208));
  INV_X1    g0008(.A(G250), .ZN(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  OAI22_X1  g0011(.A1(new_n208), .A2(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI211_X1 g0012(.A(new_n207), .B(new_n212), .C1(G68), .C2(G238), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G50), .A2(G226), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G77), .A2(G244), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G116), .A2(G270), .ZN(new_n216));
  NAND4_X1  g0016(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n203), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(G50), .B1(G58), .B2(G68), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n206), .B(new_n222), .C1(new_n225), .C2(new_n227), .ZN(G361));
  XNOR2_X1  g0028(.A(G250), .B(G257), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G264), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(G270), .Z(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(new_n219), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n231), .B(new_n235), .Z(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G58), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G13), .ZN(new_n244));
  NOR3_X1   g0044(.A1(new_n244), .A2(new_n224), .A3(G1), .ZN(new_n245));
  INV_X1    g0045(.A(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n223), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT67), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT67), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n248), .A2(new_n251), .A3(new_n223), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(G1), .B2(new_n224), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n247), .B1(new_n255), .B2(new_n246), .ZN(new_n256));
  XOR2_X1   g0056(.A(KEYINPUT8), .B(G58), .Z(new_n257));
  INV_X1    g0057(.A(KEYINPUT68), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(new_n224), .A3(G33), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  OAI21_X1  g0060(.A(KEYINPUT68), .B1(new_n260), .B2(G20), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n257), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G58), .A2(G68), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n224), .B1(new_n263), .B2(new_n246), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G20), .A2(G33), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n264), .B1(G150), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n254), .B1(new_n262), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n256), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G1), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT64), .B(G41), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n269), .B(G274), .C1(new_n270), .C2(G45), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  AOI21_X1  g0075(.A(G1), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  AND2_X1   g0077(.A1(new_n277), .A2(G226), .ZN(new_n278));
  XNOR2_X1  g0078(.A(KEYINPUT3), .B(G33), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G222), .A2(G1698), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(G223), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n279), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(G77), .B2(new_n279), .ZN(new_n284));
  XOR2_X1   g0084(.A(new_n284), .B(KEYINPUT65), .Z(new_n285));
  NAND2_X1  g0085(.A1(new_n273), .A2(KEYINPUT66), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT66), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n260), .A2(new_n274), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n287), .B1(new_n288), .B2(new_n223), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AOI211_X1 g0091(.A(new_n272), .B(new_n278), .C1(new_n285), .C2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G169), .ZN(new_n293));
  INV_X1    g0093(.A(G179), .ZN(new_n294));
  AOI211_X1 g0094(.A(new_n268), .B(new_n293), .C1(new_n294), .C2(new_n292), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n268), .A2(KEYINPUT9), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n296), .B(KEYINPUT73), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n292), .A2(G190), .B1(KEYINPUT9), .B2(new_n268), .ZN(new_n298));
  INV_X1    g0098(.A(G200), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n297), .B(new_n298), .C1(new_n299), .C2(new_n292), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n300), .A2(KEYINPUT10), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(KEYINPUT10), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n295), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G68), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G20), .ZN(new_n305));
  INV_X1    g0105(.A(new_n265), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n261), .A2(new_n259), .ZN(new_n307));
  INV_X1    g0107(.A(G77), .ZN(new_n308));
  OAI221_X1 g0108(.A(new_n305), .B1(new_n246), .B2(new_n306), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n253), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT11), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n269), .A2(new_n304), .A3(G13), .A4(G20), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT12), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n313), .A2(KEYINPUT77), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n311), .B(new_n315), .C1(new_n304), .C2(new_n255), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n313), .A2(KEYINPUT77), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n312), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT3), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G33), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n321), .A2(new_n323), .A3(G232), .A4(G1698), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT74), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT74), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n279), .A2(new_n326), .A3(G232), .A4(G1698), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n279), .A2(G226), .A3(new_n281), .ZN(new_n329));
  NAND2_X1  g0129(.A1(G33), .A2(G97), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(KEYINPUT75), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT75), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n328), .A2(new_n333), .A3(new_n329), .A4(new_n330), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n291), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT13), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n272), .B1(G238), .B2(new_n277), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n336), .B1(new_n335), .B2(new_n337), .ZN(new_n339));
  OAI21_X1  g0139(.A(G169), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT14), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n335), .A2(new_n337), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(KEYINPUT13), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT14), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(new_n346), .A3(G169), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n343), .A2(KEYINPUT76), .A3(new_n344), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT76), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n338), .B1(new_n339), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n294), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n320), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n349), .A2(new_n351), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G190), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n345), .A2(G200), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(new_n319), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G159), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n306), .A2(KEYINPUT80), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT80), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n363), .B1(new_n265), .B2(G159), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(G58), .B(G68), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n365), .B1(G20), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n321), .A2(new_n323), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n368), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT78), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n321), .A2(new_n323), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n371), .B1(new_n321), .B2(new_n323), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n224), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT7), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n370), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n376), .A2(KEYINPUT79), .A3(new_n304), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT79), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n322), .A2(G33), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT78), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n321), .A2(new_n323), .A3(new_n371), .ZN(new_n382));
  AOI21_X1  g0182(.A(G20), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n369), .B1(new_n383), .B2(KEYINPUT7), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n378), .B1(new_n384), .B2(G68), .ZN(new_n385));
  OAI211_X1 g0185(.A(KEYINPUT16), .B(new_n367), .C1(new_n377), .C2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT16), .ZN(new_n387));
  INV_X1    g0187(.A(new_n367), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n375), .B1(new_n279), .B2(G20), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n304), .B1(new_n389), .B2(new_n369), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n387), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n386), .A2(new_n391), .A3(new_n253), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n257), .A2(new_n245), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n255), .B2(new_n257), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(G169), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT81), .B1(new_n260), .B2(new_n208), .ZN(new_n398));
  OR3_X1    g0198(.A1(new_n260), .A2(new_n208), .A3(KEYINPUT81), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n279), .B1(G226), .B2(new_n281), .ZN(new_n400));
  NOR2_X1   g0200(.A1(G223), .A2(G1698), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n398), .B(new_n399), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n402), .A2(new_n291), .B1(G232), .B2(new_n277), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n397), .B1(new_n403), .B2(new_n271), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n403), .A2(new_n271), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n404), .B1(G179), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT18), .B1(new_n396), .B2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT18), .ZN(new_n409));
  AOI211_X1 g0209(.A(new_n409), .B(new_n406), .C1(new_n392), .C2(new_n395), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n254), .B(G77), .C1(G1), .C2(new_n224), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT71), .ZN(new_n413));
  XNOR2_X1  g0213(.A(new_n412), .B(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n257), .A2(new_n265), .ZN(new_n415));
  XNOR2_X1  g0215(.A(KEYINPUT15), .B(G87), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT70), .ZN(new_n417));
  OAI221_X1 g0217(.A(new_n415), .B1(new_n224), .B2(new_n308), .C1(new_n417), .C2(new_n307), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n418), .A2(new_n253), .B1(new_n308), .B2(new_n245), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n277), .A2(G244), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G238), .A2(G1698), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n279), .B(new_n422), .C1(new_n219), .C2(G1698), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(G107), .B2(new_n279), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n421), .B(new_n271), .C1(new_n424), .C2(new_n290), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n397), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n420), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT72), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n425), .A2(G179), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n420), .A2(KEYINPUT72), .A3(new_n426), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n420), .B1(G200), .B2(new_n425), .ZN(new_n434));
  INV_X1    g0234(.A(G190), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n425), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT69), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n403), .A2(new_n271), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n299), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(G190), .B2(new_n440), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n392), .A2(new_n395), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT17), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n392), .A2(KEYINPUT17), .A3(new_n395), .A4(new_n442), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n411), .A2(new_n439), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n303), .A2(new_n360), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT84), .ZN(new_n450));
  INV_X1    g0250(.A(G283), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n260), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n321), .A2(new_n323), .A3(G244), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT4), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n454), .A2(KEYINPUT83), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n452), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n455), .B1(new_n279), .B2(G250), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n456), .B1(new_n457), .B2(new_n281), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n279), .A2(G244), .A3(new_n281), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n454), .B1(new_n459), .B2(KEYINPUT83), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n450), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(KEYINPUT83), .B1(new_n453), .B2(G1698), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT4), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n368), .A2(new_n209), .ZN(new_n464));
  OAI21_X1  g0264(.A(G1698), .B1(new_n464), .B2(new_n455), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT84), .A4(new_n456), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n461), .A2(new_n466), .A3(new_n291), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT5), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n269), .B(G45), .C1(new_n468), .C2(G41), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n469), .B1(new_n270), .B2(new_n468), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G274), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n273), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n270), .A2(new_n468), .ZN(new_n474));
  OAI211_X1 g0274(.A(G257), .B(new_n473), .C1(new_n474), .C2(new_n469), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT85), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n470), .A2(new_n273), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n478), .A2(KEYINPUT85), .A3(G257), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n472), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n467), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G200), .ZN(new_n482));
  OAI21_X1  g0282(.A(KEYINPUT82), .B1(new_n306), .B2(new_n308), .ZN(new_n483));
  OR3_X1    g0283(.A1(new_n306), .A2(KEYINPUT82), .A3(new_n308), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT6), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n485), .A2(new_n210), .A3(G107), .ZN(new_n486));
  XNOR2_X1  g0286(.A(G97), .B(G107), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n486), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n483), .B(new_n484), .C1(new_n488), .C2(new_n224), .ZN(new_n489));
  INV_X1    g0289(.A(G107), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n490), .B1(new_n389), .B2(new_n369), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n253), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n245), .A2(new_n210), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n260), .A2(G1), .ZN(new_n494));
  NOR3_X1   g0294(.A1(new_n253), .A2(new_n245), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G97), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n492), .A2(new_n493), .A3(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n482), .B(new_n497), .C1(new_n435), .C2(new_n481), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n492), .A2(new_n493), .A3(new_n496), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT86), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n497), .A2(KEYINPUT86), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n467), .A2(new_n480), .A3(G179), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n397), .B1(new_n467), .B2(new_n480), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n501), .B(new_n502), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n498), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n209), .A2(new_n281), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n211), .A2(G1698), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n321), .A2(new_n507), .A3(new_n323), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(G33), .A2(G294), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n291), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(G264), .B(new_n473), .C1(new_n474), .C2(new_n469), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n512), .A2(new_n435), .A3(new_n513), .A4(new_n471), .ZN(new_n514));
  INV_X1    g0314(.A(new_n511), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n471), .B1(new_n515), .B2(new_n290), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT92), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n478), .A2(KEYINPUT92), .A3(G264), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n516), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n514), .B1(new_n520), .B2(G200), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n495), .A2(G107), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n490), .A2(G20), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n523), .A2(G1), .A3(new_n244), .ZN(new_n524));
  XNOR2_X1  g0324(.A(new_n524), .B(KEYINPUT25), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n321), .A2(new_n323), .A3(new_n224), .A4(G87), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(KEYINPUT22), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT22), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n279), .A2(new_n528), .A3(new_n224), .A4(G87), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  XOR2_X1   g0330(.A(new_n523), .B(KEYINPUT23), .Z(new_n531));
  NAND3_X1  g0331(.A1(new_n224), .A2(G33), .A3(G116), .ZN(new_n532));
  XOR2_X1   g0332(.A(new_n532), .B(KEYINPUT91), .Z(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT24), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n530), .A2(new_n533), .A3(KEYINPUT24), .A4(new_n531), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n536), .A2(new_n253), .A3(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n521), .A2(new_n522), .A3(new_n525), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n518), .A2(new_n519), .ZN(new_n540));
  INV_X1    g0340(.A(new_n516), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n540), .A2(G179), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n512), .A2(new_n471), .A3(new_n513), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(G169), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n538), .A2(new_n522), .A3(new_n525), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n539), .A2(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n478), .A2(G270), .B1(G274), .B2(new_n470), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G264), .A2(G1698), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n279), .B(new_n550), .C1(new_n211), .C2(G1698), .ZN(new_n551));
  INV_X1    g0351(.A(G303), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n368), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n551), .A2(new_n289), .A3(new_n286), .A4(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n397), .B1(new_n549), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(G116), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n248), .A2(new_n223), .B1(G20), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(G20), .B1(G33), .B2(G283), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n260), .A2(G97), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT90), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n560), .B1(new_n558), .B2(new_n559), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n557), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT20), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(KEYINPUT20), .B(new_n557), .C1(new_n561), .C2(new_n562), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n495), .A2(G116), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n245), .A2(new_n556), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n555), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT21), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n549), .A2(new_n554), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(G200), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n567), .A2(new_n568), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n549), .A2(G190), .A3(new_n554), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n569), .A4(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n574), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n579), .A2(G179), .A3(new_n570), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n555), .A2(new_n570), .A3(KEYINPUT21), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n573), .A2(new_n578), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n548), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT89), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n261), .A2(new_n259), .A3(G97), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT19), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(KEYINPUT87), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n224), .B1(new_n330), .B2(new_n586), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n208), .A2(new_n210), .A3(new_n490), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n321), .A2(new_n323), .A3(new_n224), .A4(G68), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT87), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n585), .A2(new_n594), .A3(new_n586), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n588), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT88), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n588), .A2(KEYINPUT88), .A3(new_n593), .A4(new_n595), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n253), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n417), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n495), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n417), .A2(new_n245), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n473), .B(G250), .C1(G1), .C2(new_n275), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n269), .A2(G45), .A3(G274), .ZN(new_n606));
  MUX2_X1   g0406(.A(G238), .B(G244), .S(G1698), .Z(new_n607));
  AOI22_X1  g0407(.A1(new_n607), .A2(new_n279), .B1(G33), .B2(G116), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n605), .B(new_n606), .C1(new_n290), .C2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n397), .ZN(new_n610));
  INV_X1    g0410(.A(new_n609), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n294), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n604), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(G190), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n495), .A2(G87), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n600), .A2(new_n603), .A3(new_n614), .A4(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n611), .A2(new_n299), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n584), .B1(new_n613), .B2(new_n618), .ZN(new_n619));
  OR2_X1    g0419(.A1(new_n616), .A2(new_n617), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n604), .A2(new_n610), .A3(new_n612), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(KEYINPUT89), .A3(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n506), .A2(new_n583), .A3(new_n619), .A4(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n449), .A2(new_n623), .ZN(G372));
  OAI21_X1  g0424(.A(KEYINPUT79), .B1(new_n376), .B2(new_n304), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n384), .A2(new_n378), .A3(G68), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n388), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n254), .B1(new_n627), .B2(KEYINPUT16), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n394), .B1(new_n628), .B2(new_n391), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n409), .B1(new_n629), .B2(new_n406), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n396), .A2(KEYINPUT18), .A3(new_n407), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n433), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n354), .B1(new_n633), .B2(new_n358), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n632), .B1(new_n634), .B2(new_n447), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n301), .A2(new_n302), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n295), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n505), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n619), .A2(new_n622), .A3(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n639), .A2(KEYINPUT26), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n499), .B1(new_n503), .B2(new_n504), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT94), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  OAI211_X1 g0444(.A(KEYINPUT94), .B(new_n499), .C1(new_n503), .C2(new_n504), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n643), .A2(new_n644), .A3(new_n620), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n610), .B(KEYINPUT93), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n647), .A2(new_n604), .A3(new_n612), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n573), .A2(new_n580), .A3(new_n581), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n545), .B2(new_n546), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n620), .A2(new_n498), .A3(new_n505), .A4(new_n539), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n646), .B(new_n648), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n640), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n637), .B1(new_n449), .B2(new_n653), .ZN(G369));
  NOR3_X1   g0454(.A1(new_n244), .A2(G1), .A3(G20), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT27), .ZN(new_n656));
  OR3_X1    g0456(.A1(new_n655), .A2(KEYINPUT95), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G213), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n658), .B1(new_n655), .B2(new_n656), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT95), .B1(new_n655), .B2(new_n656), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT96), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G343), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n576), .B2(new_n569), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n582), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n649), .A2(new_n664), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(G330), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT97), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n663), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n671), .A2(new_n546), .ZN(new_n672));
  OAI22_X1  g0472(.A1(new_n548), .A2(new_n672), .B1(new_n547), .B2(new_n663), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n649), .A2(new_n663), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(new_n548), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n547), .A2(new_n671), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n674), .A2(new_n678), .ZN(G399));
  INV_X1    g0479(.A(new_n270), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n204), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n590), .A2(G116), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G1), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n226), .B2(new_n681), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n663), .B1(new_n640), .B2(new_n652), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT29), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n643), .A2(new_n620), .A3(new_n645), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(KEYINPUT26), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n619), .A2(new_n622), .A3(new_n644), .A4(new_n638), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n648), .B1(new_n651), .B2(new_n650), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n663), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(KEYINPUT29), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n687), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(G330), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT98), .B1(new_n623), .B2(new_n671), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n619), .A2(new_n622), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n498), .A2(new_n505), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n699), .A2(new_n548), .A3(new_n582), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT98), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n698), .A2(new_n700), .A3(new_n701), .A4(new_n663), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n478), .A2(G270), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n704), .A2(G179), .A3(new_n471), .A4(new_n554), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n515), .A2(new_n290), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n705), .A2(new_n609), .A3(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n707), .A2(new_n467), .A3(new_n480), .A4(new_n540), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT30), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n481), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n711), .A2(KEYINPUT30), .A3(new_n540), .A4(new_n707), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n579), .A2(G179), .ZN(new_n713));
  INV_X1    g0513(.A(new_n520), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n713), .A2(new_n481), .A3(new_n609), .A4(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n710), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n671), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT31), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n717), .B(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n696), .B1(new_n703), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n695), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n685), .B1(new_n722), .B2(G1), .ZN(G364));
  INV_X1    g0523(.A(new_n670), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n224), .A2(G13), .A3(G45), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n681), .A2(G1), .A3(new_n725), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n724), .B(new_n726), .C1(G330), .C2(new_n667), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n223), .B1(G20), .B2(new_n397), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT100), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n294), .A2(new_n299), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n224), .A2(G190), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n304), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n299), .A2(G179), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(new_n490), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G179), .A2(G200), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n731), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G159), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT32), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n224), .A2(new_n435), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n730), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n734), .ZN(new_n744));
  OAI22_X1  g0544(.A1(new_n743), .A2(new_n246), .B1(new_n744), .B2(new_n208), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n294), .A2(G200), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n731), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n737), .A2(G190), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n748), .A2(G20), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI221_X1 g0550(.A(new_n279), .B1(new_n747), .B2(new_n308), .C1(new_n750), .C2(new_n210), .ZN(new_n751));
  OR4_X1    g0551(.A1(new_n736), .A2(new_n741), .A3(new_n745), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n742), .A2(new_n746), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n733), .B(new_n752), .C1(G58), .C2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n732), .ZN(new_n756));
  INV_X1    g0556(.A(G317), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(KEYINPUT33), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n757), .A2(KEYINPUT33), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n756), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n743), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G326), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n739), .A2(G329), .ZN(new_n763));
  INV_X1    g0563(.A(new_n735), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G283), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n760), .A2(new_n762), .A3(new_n763), .A4(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(G294), .B2(new_n749), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n279), .B1(new_n754), .B2(G322), .ZN(new_n768));
  OAI211_X1 g0568(.A(new_n767), .B(new_n768), .C1(new_n552), .C2(new_n744), .ZN(new_n769));
  INV_X1    g0569(.A(new_n747), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n769), .B1(G311), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n729), .B1(new_n755), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n726), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n372), .A2(new_n373), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n204), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT99), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n227), .A2(new_n275), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n777), .B(new_n778), .C1(new_n275), .C2(new_n239), .ZN(new_n779));
  INV_X1    g0579(.A(G355), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n279), .A2(new_n204), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n779), .B1(G116), .B2(new_n204), .C1(new_n780), .C2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G13), .A2(G33), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n729), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n772), .A2(new_n773), .A3(new_n787), .ZN(new_n788));
  XOR2_X1   g0588(.A(new_n788), .B(KEYINPUT101), .Z(new_n789));
  INV_X1    g0589(.A(new_n785), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n789), .B1(new_n667), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g0591(.A1(new_n727), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(G396));
  AOI21_X1  g0593(.A(new_n663), .B1(new_n414), .B2(new_n419), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n429), .A2(new_n431), .A3(new_n432), .A4(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n439), .B2(new_n794), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n686), .A2(new_n797), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n663), .B(new_n796), .C1(new_n640), .C2(new_n652), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(new_n721), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n726), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n797), .A2(new_n783), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n729), .A2(new_n783), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n308), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n743), .A2(new_n552), .B1(new_n747), .B2(new_n556), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(G283), .B2(new_n756), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT102), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n279), .B(new_n808), .C1(G294), .C2(new_n754), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n764), .A2(G87), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n739), .A2(G311), .ZN(new_n811));
  INV_X1    g0611(.A(new_n744), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n812), .A2(G107), .B1(new_n749), .B2(G97), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n809), .A2(new_n810), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n775), .B1(G58), .B2(new_n749), .ZN(new_n815));
  AOI22_X1  g0615(.A1(G68), .A2(new_n764), .B1(new_n739), .B2(G132), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n815), .B(new_n816), .C1(new_n246), .C2(new_n744), .ZN(new_n817));
  XOR2_X1   g0617(.A(new_n817), .B(KEYINPUT103), .Z(new_n818));
  AOI22_X1  g0618(.A1(G143), .A2(new_n754), .B1(new_n770), .B2(G159), .ZN(new_n819));
  INV_X1    g0619(.A(G137), .ZN(new_n820));
  INV_X1    g0620(.A(G150), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n819), .B1(new_n820), .B2(new_n743), .C1(new_n821), .C2(new_n732), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT34), .Z(new_n823));
  OAI21_X1  g0623(.A(new_n814), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n729), .ZN(new_n825));
  NAND4_X1  g0625(.A1(new_n803), .A2(new_n773), .A3(new_n805), .A4(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT104), .Z(new_n827));
  NAND2_X1  g0627(.A1(new_n802), .A2(new_n827), .ZN(G384));
  INV_X1    g0628(.A(new_n637), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n449), .B1(new_n687), .B2(new_n694), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT106), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n832), .B1(new_n320), .B2(new_n671), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n832), .B(new_n671), .C1(new_n316), .C2(new_n318), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n353), .B2(new_n358), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n353), .A2(new_n358), .A3(new_n836), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n719), .B1(new_n697), .B2(new_n702), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n840), .A2(new_n841), .A3(new_n797), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT40), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT38), .ZN(new_n844));
  INV_X1    g0644(.A(new_n662), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n392), .A2(new_n395), .B1(new_n406), .B2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT37), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n847), .A2(new_n848), .A3(new_n443), .ZN(new_n849));
  INV_X1    g0649(.A(new_n443), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT37), .B1(new_n850), .B2(new_n846), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n629), .A2(new_n845), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n445), .A2(new_n446), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n855), .B1(new_n856), .B2(new_n632), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n844), .B1(new_n853), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n367), .B1(new_n377), .B2(new_n385), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n387), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n394), .B1(new_n628), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n861), .A2(new_n845), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n411), .B2(new_n447), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n443), .B1(new_n861), .B2(new_n406), .ZN(new_n864));
  OAI21_X1  g0664(.A(KEYINPUT37), .B1(new_n864), .B2(new_n862), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n849), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n863), .A2(new_n866), .A3(KEYINPUT38), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n843), .B1(new_n858), .B2(new_n867), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n840), .A2(new_n841), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n863), .A2(new_n866), .A3(KEYINPUT38), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT38), .B1(new_n863), .B2(new_n866), .ZN(new_n871));
  OAI21_X1  g0671(.A(KEYINPUT107), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NOR3_X1   g0672(.A1(new_n850), .A2(new_n846), .A3(KEYINPUT37), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n628), .A2(new_n860), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n395), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n662), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n407), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(new_n443), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n873), .B1(new_n878), .B2(KEYINPUT37), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n876), .B1(new_n856), .B2(new_n632), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n844), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT107), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(new_n882), .A3(new_n867), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n869), .A2(new_n872), .A3(new_n796), .A4(new_n883), .ZN(new_n884));
  AOI221_X4 g0684(.A(new_n696), .B1(new_n842), .B2(new_n868), .C1(new_n884), .C2(new_n843), .ZN(new_n885));
  NOR3_X1   g0685(.A1(new_n449), .A2(new_n841), .A3(new_n696), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n887), .B(KEYINPUT109), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n884), .A2(new_n843), .B1(new_n842), .B2(new_n868), .ZN(new_n889));
  INV_X1    g0689(.A(new_n449), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n703), .A2(new_n720), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT110), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT108), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n888), .A2(KEYINPUT110), .A3(new_n892), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n896), .B1(new_n895), .B2(new_n897), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n831), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n900), .ZN(new_n902));
  INV_X1    g0702(.A(new_n831), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n902), .A2(new_n903), .A3(new_n898), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n633), .A2(new_n663), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n799), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n839), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(new_n837), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n872), .A2(new_n883), .A3(new_n907), .A4(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT39), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n854), .B1(new_n411), .B2(new_n447), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT38), .B1(new_n912), .B2(new_n852), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n911), .B1(new_n870), .B2(new_n913), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n341), .A2(new_n347), .ZN(new_n915));
  INV_X1    g0715(.A(new_n352), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(new_n320), .A3(new_n663), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n881), .A2(KEYINPUT39), .A3(new_n867), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n914), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n632), .A2(new_n662), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n910), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n905), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(G1), .B1(new_n244), .B2(G20), .ZN(new_n926));
  INV_X1    g0726(.A(new_n924), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n901), .A2(new_n904), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT35), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n488), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(G116), .A3(new_n225), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n932), .B(KEYINPUT105), .Z(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n930), .B2(new_n488), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT36), .ZN(new_n935));
  OAI21_X1  g0735(.A(G77), .B1(new_n218), .B2(new_n304), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n936), .A2(new_n226), .B1(G50), .B2(new_n304), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(G1), .A3(new_n244), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n929), .A2(new_n935), .A3(new_n938), .ZN(G367));
  NAND2_X1  g0739(.A1(new_n725), .A2(G1), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n722), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n497), .A2(new_n663), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n699), .A2(new_n943), .B1(new_n641), .B2(new_n663), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n678), .A2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT45), .Z(new_n946));
  NOR2_X1   g0746(.A1(new_n678), .A2(new_n944), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT44), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT113), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n946), .B(new_n948), .C1(new_n674), .C2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n674), .A2(new_n949), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n950), .B(new_n951), .Z(new_n952));
  INV_X1    g0752(.A(new_n676), .ZN(new_n953));
  INV_X1    g0753(.A(new_n675), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n953), .B1(new_n673), .B2(new_n954), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n670), .B(new_n955), .Z(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n942), .B1(new_n952), .B2(new_n957), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n681), .B(KEYINPUT41), .Z(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n941), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n600), .A2(new_n603), .A3(new_n615), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n671), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n620), .A2(new_n963), .ZN(new_n964));
  MUX2_X1   g0764(.A(new_n963), .B(new_n964), .S(new_n648), .Z(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT43), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n944), .B(KEYINPUT111), .Z(new_n967));
  OR2_X1    g0767(.A1(new_n967), .A2(new_n547), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n671), .B1(new_n968), .B2(new_n505), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n944), .A2(new_n676), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT42), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n966), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(KEYINPUT112), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n969), .A2(new_n971), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT43), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n974), .A2(new_n975), .A3(new_n965), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT112), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n977), .B(new_n966), .C1(new_n969), .C2(new_n971), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n973), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n979), .B1(new_n674), .B2(new_n967), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n674), .A2(new_n967), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n973), .A2(new_n976), .A3(new_n981), .A4(new_n978), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n961), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n726), .B1(new_n965), .B2(new_n785), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n761), .A2(G311), .B1(new_n739), .B2(G317), .ZN(new_n985));
  INV_X1    g0785(.A(G294), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n985), .B1(new_n986), .B2(new_n732), .C1(new_n552), .C2(new_n753), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n987), .B1(G283), .B2(new_n770), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n749), .A2(G107), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n812), .A2(G116), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT46), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n735), .A2(new_n210), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n774), .A2(new_n992), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n988), .A2(new_n989), .A3(new_n991), .A4(new_n993), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n761), .A2(G143), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n744), .A2(new_n218), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n753), .A2(new_n821), .B1(new_n738), .B2(new_n820), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n996), .B(new_n997), .C1(G68), .C2(new_n749), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n756), .A2(G159), .ZN(new_n999));
  AOI22_X1  g0799(.A1(G50), .A2(new_n770), .B1(new_n764), .B2(G77), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n998), .A2(new_n279), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n994), .B1(new_n995), .B2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT47), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n729), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n777), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n786), .B1(new_n204), .B2(new_n417), .C1(new_n1005), .C2(new_n231), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n984), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n983), .A2(new_n1007), .ZN(G387));
  INV_X1    g0808(.A(KEYINPUT117), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n942), .A2(new_n956), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT115), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n681), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1011), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n942), .A2(KEYINPUT116), .A3(new_n956), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT116), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n957), .B2(new_n722), .ZN(new_n1017));
  OAI21_X1  g0817(.A(KEYINPUT115), .B1(new_n1010), .B2(new_n681), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n747), .A2(new_n304), .B1(new_n738), .B2(new_n821), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n992), .B(new_n1020), .C1(G50), .C2(new_n754), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n601), .A2(new_n749), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G77), .A2(new_n812), .B1(new_n756), .B2(new_n257), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n775), .B1(G159), .B2(new_n761), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G322), .A2(new_n761), .B1(new_n756), .B2(G311), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n552), .B2(new_n747), .C1(new_n757), .C2(new_n753), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT48), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n451), .B2(new_n750), .C1(new_n986), .C2(new_n744), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT49), .Z(new_n1030));
  NAND2_X1  g0830(.A1(new_n739), .A2(G326), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n775), .B(new_n1031), .C1(new_n556), .C2(new_n735), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1025), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n729), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1034), .B(new_n773), .C1(new_n673), .C2(new_n790), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1005), .B1(G45), .B2(new_n235), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n682), .B(new_n275), .C1(new_n304), .C2(new_n308), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT114), .Z(new_n1038));
  NAND2_X1  g0838(.A1(new_n257), .A2(new_n246), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT50), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1036), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(G107), .B2(new_n204), .C1(new_n682), .C2(new_n781), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1035), .B1(new_n786), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n957), .B2(new_n940), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1009), .B1(new_n1019), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1019), .A2(new_n1009), .A3(new_n1044), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(G393));
  NAND2_X1  g0848(.A1(new_n967), .A2(new_n785), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n786), .B1(new_n210), .B2(new_n204), .C1(new_n1005), .C2(new_n242), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G317), .A2(new_n761), .B1(new_n754), .B2(G311), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT52), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n750), .A2(new_n556), .B1(new_n986), .B2(new_n747), .ZN(new_n1053));
  INV_X1    g0853(.A(G322), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n368), .B1(new_n738), .B2(new_n1054), .ZN(new_n1055));
  NOR4_X1   g0855(.A1(new_n1052), .A2(new_n736), .A3(new_n1053), .A4(new_n1055), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(new_n451), .B2(new_n744), .C1(new_n552), .C2(new_n732), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G87), .A2(new_n764), .B1(new_n739), .B2(G143), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1058), .B(new_n774), .C1(new_n304), .C2(new_n744), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT118), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n743), .A2(new_n821), .B1(new_n753), .B2(new_n361), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT51), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n756), .A2(G50), .B1(new_n749), .B2(G77), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n257), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1063), .B1(new_n1064), .B2(new_n747), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT119), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1060), .A2(new_n1062), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1057), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n726), .B1(new_n1068), .B2(new_n729), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1049), .A2(new_n1050), .A3(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n950), .B(new_n951), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1070), .B1(new_n1071), .B2(new_n941), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n681), .B1(new_n1011), .B2(new_n1071), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n952), .A2(new_n1010), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1072), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(G390));
  NAND3_X1  g0876(.A1(new_n721), .A2(new_n796), .A3(new_n909), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n907), .A2(new_n909), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n918), .A2(new_n1079), .B1(new_n914), .B2(new_n920), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n918), .A2(KEYINPUT120), .ZN(new_n1081));
  OR3_X1    g0881(.A1(new_n353), .A2(KEYINPUT120), .A3(new_n671), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n858), .A2(new_n867), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n796), .B(new_n663), .C1(new_n691), .C2(new_n692), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n906), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n909), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1078), .B1(new_n1080), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1089));
  AND2_X1   g0889(.A1(new_n914), .A2(new_n920), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n919), .B1(new_n907), .B2(new_n909), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1089), .B(new_n1077), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n940), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1090), .A2(new_n784), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n804), .A2(new_n1064), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n732), .A2(new_n820), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n744), .A2(new_n821), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(KEYINPUT121), .B(KEYINPUT53), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1099), .B(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(G132), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n753), .A2(new_n1102), .B1(new_n735), .B2(new_n246), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(G128), .B2(new_n761), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n749), .A2(G159), .ZN(new_n1105));
  XOR2_X1   g0905(.A(KEYINPUT54), .B(G143), .Z(new_n1106));
  AOI21_X1  g0906(.A(new_n368), .B1(new_n770), .B2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1101), .A2(new_n1104), .A3(new_n1105), .A4(new_n1107), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1098), .B(new_n1108), .C1(G125), .C2(new_n739), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n743), .A2(new_n451), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(G87), .A2(new_n812), .B1(new_n764), .B2(G68), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(G97), .A2(new_n770), .B1(new_n739), .B2(G294), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n756), .A2(G107), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n279), .B1(new_n749), .B2(G77), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1111), .A2(new_n1112), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n1110), .B(new_n1115), .C1(G116), .C2(new_n754), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n729), .B1(new_n1109), .B2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1096), .A2(new_n773), .A3(new_n1097), .A4(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1095), .A2(new_n1118), .ZN(new_n1119));
  NOR3_X1   g0919(.A1(new_n829), .A2(new_n830), .A3(new_n886), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n891), .A2(G330), .A3(new_n796), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n840), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1085), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1123), .A2(new_n1124), .A3(new_n1077), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n1123), .A2(new_n1077), .B1(new_n799), .B2(new_n906), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1121), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n1093), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n681), .B1(new_n1128), .B2(new_n1094), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1119), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(G378));
  OAI21_X1  g0933(.A(new_n1120), .B1(new_n1093), .B2(new_n1127), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n268), .A2(new_n845), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  XOR2_X1   g0936(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n303), .A2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n303), .A2(new_n1138), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1136), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  OR2_X1    g0941(.A1(new_n303), .A2(new_n1138), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n303), .A2(new_n1138), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n1135), .A3(new_n1143), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n924), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1147), .A2(new_n910), .A3(new_n921), .A4(new_n923), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n889), .A2(G330), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n885), .A2(new_n1148), .A3(new_n1146), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1134), .A2(KEYINPUT57), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n1013), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(KEYINPUT124), .ZN(new_n1155));
  AND2_X1   g0955(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n1134), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT57), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT124), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1153), .A2(new_n1160), .A3(new_n1013), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1155), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1156), .A2(new_n940), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n726), .B1(new_n1147), .B2(new_n783), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(G33), .A2(G41), .ZN(new_n1165));
  AOI211_X1 g0965(.A(G50), .B(new_n1165), .C1(new_n775), .C2(new_n680), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n750), .A2(new_n304), .B1(new_n753), .B2(new_n490), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G77), .A2(new_n812), .B1(new_n764), .B2(G58), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n739), .A2(G283), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n1168), .A2(new_n775), .A3(new_n680), .A4(new_n1169), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n1170), .B(KEYINPUT122), .Z(new_n1171));
  AOI211_X1 g0971(.A(new_n1167), .B(new_n1171), .C1(G97), .C2(new_n756), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1172), .B1(new_n556), .B2(new_n743), .C1(new_n417), .C2(new_n747), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT58), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1166), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT123), .Z(new_n1176));
  INV_X1    g0976(.A(G124), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1165), .B1(new_n738), .B2(new_n1177), .C1(new_n361), .C2(new_n735), .ZN(new_n1178));
  INV_X1    g0978(.A(G128), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n753), .A2(new_n1179), .B1(new_n747), .B2(new_n820), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1106), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n750), .A2(new_n821), .B1(new_n1181), .B2(new_n744), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1180), .B(new_n1182), .C1(G125), .C2(new_n761), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n1102), .B2(new_n732), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT59), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1176), .B1(new_n1174), .B2(new_n1173), .C1(new_n1178), .C2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n729), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n804), .A2(new_n246), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1164), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1163), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1162), .A2(new_n1191), .ZN(G375));
  NAND2_X1  g0992(.A1(new_n739), .A2(G303), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n754), .A2(G283), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n279), .B1(new_n812), .B2(G97), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1022), .A2(new_n1193), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n743), .A2(new_n986), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n732), .A2(new_n556), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n308), .A2(new_n735), .B1(new_n747), .B2(new_n490), .ZN(new_n1199));
  NOR4_X1   g0999(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(G159), .A2(new_n812), .B1(new_n770), .B2(G150), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n246), .B2(new_n750), .C1(new_n820), .C2(new_n753), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n761), .A2(G132), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT125), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1181), .A2(new_n732), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n774), .B1(new_n218), .B2(new_n735), .C1(new_n1179), .C2(new_n738), .ZN(new_n1206));
  NOR4_X1   g1006(.A1(new_n1202), .A2(new_n1204), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n729), .B1(new_n1200), .B2(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n773), .B(new_n1208), .C1(new_n909), .C2(new_n784), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(new_n304), .B2(new_n804), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1127), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1210), .B1(new_n1211), .B2(new_n940), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1121), .A2(new_n1127), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n959), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1212), .B1(new_n1214), .B2(new_n1128), .ZN(G381));
  NOR2_X1   g1015(.A1(G375), .A2(G378), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(G381), .A2(G384), .ZN(new_n1217));
  AND3_X1   g1017(.A1(new_n983), .A2(new_n1007), .A3(new_n1075), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1047), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1219), .A2(G396), .A3(new_n1045), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .A4(new_n1220), .ZN(G407));
  INV_X1    g1021(.A(G343), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n658), .B1(new_n1216), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(G407), .ZN(G409));
  OAI21_X1  g1024(.A(G396), .B1(new_n1219), .B2(new_n1045), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1046), .A2(new_n792), .A3(new_n1047), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(G387), .A2(G390), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n983), .A2(new_n1007), .A3(new_n1075), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1227), .A2(new_n1230), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1225), .A2(new_n1226), .A3(new_n1229), .A4(new_n1228), .ZN(new_n1232));
  AND3_X1   g1032(.A1(new_n1231), .A2(new_n1232), .A3(KEYINPUT127), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT127), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1153), .A2(new_n1160), .A3(new_n1013), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1160), .B1(new_n1153), .B2(new_n1013), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT57), .B1(new_n1156), .B2(new_n1134), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(G378), .B1(new_n1239), .B2(new_n1190), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT60), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1213), .A2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1121), .A2(new_n1127), .A3(KEYINPUT60), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1242), .A2(new_n1129), .A3(new_n1013), .A4(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1212), .ZN(new_n1245));
  INV_X1    g1045(.A(G384), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1244), .A2(G384), .A3(new_n1212), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n658), .A2(G343), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1156), .A2(new_n959), .A3(new_n1134), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1191), .A2(new_n1132), .A3(new_n1253), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1240), .A2(new_n1250), .A3(new_n1252), .A4(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(KEYINPUT62), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1251), .B1(G375), .B2(G378), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT62), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1257), .A2(new_n1258), .A3(new_n1250), .A4(new_n1254), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1256), .A2(new_n1259), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1132), .B1(new_n1162), .B2(new_n1191), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1254), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(new_n1262), .A2(new_n1263), .A3(new_n1251), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1251), .A2(G2897), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  XNOR2_X1  g1066(.A(new_n1249), .B(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1261), .B1(new_n1264), .B2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1235), .B1(new_n1260), .B2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT61), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1264), .A2(KEYINPUT63), .A3(new_n1250), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT63), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1240), .A2(new_n1252), .A3(new_n1254), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1249), .B(new_n1265), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1272), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1255), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1270), .B(new_n1271), .C1(new_n1275), .C2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1269), .A2(new_n1277), .ZN(G405));
  NAND2_X1  g1078(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1216), .A2(new_n1262), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1249), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1280), .A2(new_n1249), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1279), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  OR2_X1    g1084(.A1(new_n1216), .A2(new_n1262), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1250), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1286), .A2(new_n1232), .A3(new_n1231), .A4(new_n1281), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1284), .A2(new_n1287), .ZN(G402));
endmodule


