//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 1 0 0 0 1 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n805, new_n806,
    new_n808, new_n809, new_n810, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n876, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936;
  XNOR2_X1  g000(.A(KEYINPUT86), .B(G50gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G228gat), .A2(G233gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(KEYINPUT88), .ZN(new_n208));
  XNOR2_X1  g007(.A(G155gat), .B(G162gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210));
  AOI22_X1  g009(.A1(new_n209), .A2(KEYINPUT77), .B1(KEYINPUT2), .B2(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(G155gat), .B(G162gat), .Z(new_n212));
  INV_X1    g011(.A(KEYINPUT77), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G141gat), .B(G148gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n211), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT78), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n212), .B1(new_n215), .B2(KEYINPUT2), .ZN(new_n220));
  NAND4_X1  g019(.A1(new_n211), .A2(new_n214), .A3(KEYINPUT78), .A4(new_n216), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n224), .A2(KEYINPUT82), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(KEYINPUT82), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT29), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(G197gat), .B(G204gat), .ZN(new_n228));
  XOR2_X1   g027(.A(KEYINPUT75), .B(KEYINPUT22), .Z(new_n229));
  INV_X1    g028(.A(G211gat), .ZN(new_n230));
  INV_X1    g029(.A(G218gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n228), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G211gat), .B(G218gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n235), .B(KEYINPUT76), .Z(new_n236));
  NOR2_X1   g035(.A1(new_n227), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n223), .B1(new_n235), .B2(KEYINPUT29), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n208), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(G22gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(KEYINPUT3), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n235), .A2(KEYINPUT29), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n207), .B1(new_n244), .B2(new_n239), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n243), .B(new_n245), .C1(new_n227), .C2(new_n236), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n241), .A2(new_n242), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT89), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n242), .B1(new_n241), .B2(new_n246), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI211_X1 g050(.A(new_n248), .B(new_n242), .C1(new_n241), .C2(new_n246), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n206), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n206), .B(KEYINPUT87), .Z(new_n254));
  INV_X1    g053(.A(new_n247), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n254), .B1(new_n255), .B2(new_n250), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G227gat), .A2(G233gat), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G120gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G113gat), .ZN(new_n261));
  INV_X1    g060(.A(G113gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G120gat), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT1), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(G127gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G134gat), .ZN(new_n266));
  INV_X1    g065(.A(G127gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n264), .B(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G134gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT69), .ZN(new_n272));
  AND2_X1   g071(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n273));
  NOR2_X1   g072(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n272), .B1(new_n275), .B2(G190gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(KEYINPUT27), .B(G183gat), .ZN(new_n277));
  INV_X1    g076(.A(G190gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(KEYINPUT69), .A3(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n280));
  NAND3_X1  g079(.A1(new_n276), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n277), .A2(KEYINPUT28), .A3(new_n278), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n276), .A2(new_n279), .A3(KEYINPUT71), .A4(new_n280), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n284), .A3(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT66), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT66), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n289), .B1(G169gat), .B2(G176gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT26), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G169gat), .ZN(new_n294));
  INV_X1    g093(.A(G176gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n287), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n296), .B1(KEYINPUT26), .B2(new_n297), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n293), .A2(new_n298), .B1(G183gat), .B2(G190gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT25), .ZN(new_n300));
  NAND3_X1  g099(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT67), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n302), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G183gat), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n303), .A2(KEYINPUT67), .B1(new_n307), .B2(new_n278), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n306), .A2(new_n308), .B1(new_n291), .B2(KEYINPUT23), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT23), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n297), .B1(new_n296), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n300), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n287), .A2(KEYINPUT23), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT65), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n287), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT25), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n301), .A2(KEYINPUT64), .B1(new_n307), .B2(new_n278), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n318), .B(new_n304), .C1(KEYINPUT64), .C2(new_n301), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n317), .A2(new_n319), .A3(new_n311), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT68), .B1(new_n312), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n305), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n322), .A2(new_n308), .A3(new_n301), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n291), .A2(KEYINPUT23), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(new_n311), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT25), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT68), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n317), .A2(new_n319), .A3(new_n311), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  AOI221_X4 g128(.A(new_n271), .B1(new_n286), .B2(new_n299), .C1(new_n321), .C2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n271), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n321), .A2(new_n329), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n286), .A2(new_n299), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n259), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT32), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT33), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G15gat), .B(G43gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(G71gat), .B(G99gat), .ZN(new_n340));
  XOR2_X1   g139(.A(new_n339), .B(new_n340), .Z(new_n341));
  NAND3_X1  g140(.A1(new_n336), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n341), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n335), .B(KEYINPUT32), .C1(new_n337), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  OR3_X1    g145(.A1(new_n330), .A2(new_n334), .A3(new_n259), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n349), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT72), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n342), .A2(new_n352), .A3(new_n344), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n352), .B1(new_n342), .B2(new_n344), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n351), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AND4_X1   g154(.A1(KEYINPUT35), .A2(new_n257), .A3(new_n350), .A4(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT0), .B(G57gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n357), .B(G85gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(G1gat), .B(G29gat), .ZN(new_n359));
  XOR2_X1   g158(.A(new_n358), .B(new_n359), .Z(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n225), .A2(new_n226), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n271), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n266), .A2(new_n270), .A3(KEYINPUT80), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT79), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n243), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n239), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n362), .A2(new_n366), .A3(new_n368), .A4(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT83), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n366), .A2(new_n368), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n373), .A2(KEYINPUT83), .A3(new_n362), .A4(new_n369), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n271), .A2(new_n239), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT4), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT84), .ZN(new_n379));
  INV_X1    g178(.A(new_n376), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(KEYINPUT4), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n380), .A2(KEYINPUT84), .A3(KEYINPUT4), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(G225gat), .A2(G233gat), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n386), .A2(KEYINPUT5), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n375), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n381), .A2(new_n378), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n385), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n391), .B1(new_n372), .B2(new_n374), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n376), .B1(new_n366), .B2(new_n239), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT5), .B1(new_n393), .B2(new_n385), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g194(.A(KEYINPUT6), .B(new_n361), .C1(new_n389), .C2(new_n395), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n388), .B(new_n360), .C1(new_n394), .C2(new_n392), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT6), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OR2_X1    g198(.A1(new_n392), .A2(new_n394), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n360), .B1(new_n400), .B2(new_n388), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n396), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT30), .ZN(new_n403));
  INV_X1    g202(.A(new_n236), .ZN(new_n404));
  AND2_X1   g203(.A1(G226gat), .A2(G233gat), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n333), .A2(new_n326), .A3(new_n328), .A4(new_n405), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n332), .A2(new_n333), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n405), .A2(KEYINPUT29), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n404), .B(new_n406), .C1(new_n407), .C2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n333), .A2(new_n326), .A3(new_n328), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n407), .A2(new_n405), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n410), .B1(new_n412), .B2(new_n404), .ZN(new_n413));
  XOR2_X1   g212(.A(G8gat), .B(G36gat), .Z(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(G64gat), .ZN(new_n415));
  INV_X1    g214(.A(G92gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n403), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n418), .B1(new_n413), .B2(new_n417), .ZN(new_n419));
  INV_X1    g218(.A(new_n413), .ZN(new_n420));
  INV_X1    g219(.A(new_n417), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n403), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n419), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n402), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT35), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n360), .B(KEYINPUT90), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n427), .B1(new_n400), .B2(new_n388), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n396), .B1(new_n399), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n346), .A2(new_n349), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n351), .A2(new_n345), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n257), .A2(new_n429), .A3(new_n432), .A4(new_n423), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n356), .A2(new_n425), .B1(new_n426), .B2(new_n433), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n372), .A2(new_n374), .B1(new_n382), .B2(new_n383), .ZN(new_n435));
  OR3_X1    g234(.A1(new_n435), .A2(KEYINPUT39), .A3(new_n385), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n393), .A2(new_n385), .ZN(new_n437));
  OAI211_X1 g236(.A(KEYINPUT39), .B(new_n437), .C1(new_n435), .C2(new_n385), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n427), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT40), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n428), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n423), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n436), .A2(KEYINPUT40), .A3(new_n427), .A4(new_n438), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n441), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n389), .A2(new_n395), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n398), .B(new_n397), .C1(new_n445), .C2(new_n427), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT37), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n420), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n413), .A2(KEYINPUT37), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n417), .A3(new_n449), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n450), .A2(KEYINPUT38), .B1(new_n420), .B2(new_n421), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT38), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n236), .B(new_n406), .C1(new_n407), .C2(new_n409), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n453), .B(KEYINPUT37), .C1(new_n412), .C2(new_n236), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n448), .A2(new_n452), .A3(new_n417), .A4(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n446), .A2(new_n396), .A3(new_n451), .A4(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n444), .A2(new_n456), .A3(new_n257), .ZN(new_n457));
  INV_X1    g256(.A(new_n257), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n424), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n355), .A2(KEYINPUT36), .A3(new_n350), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT74), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT36), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n462), .B1(new_n430), .B2(new_n431), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT74), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n355), .A2(new_n464), .A3(KEYINPUT36), .A4(new_n350), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n461), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n457), .A2(new_n459), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n434), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(G50gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT93), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT93), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(G50gat), .ZN(new_n472));
  INV_X1    g271(.A(G43gat), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n470), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n469), .A2(G43gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT94), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT15), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n473), .A2(G50gat), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(new_n475), .A3(KEYINPUT15), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(G29gat), .A2(G36gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(KEYINPUT92), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT92), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n485), .A2(G29gat), .A3(G36gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n488));
  OR3_X1    g287(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT15), .B1(new_n474), .B2(new_n475), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n490), .B1(new_n491), .B2(new_n477), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT95), .B1(new_n482), .B2(new_n492), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n490), .A2(new_n481), .ZN(new_n494));
  INV_X1    g293(.A(new_n481), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n495), .B1(new_n491), .B2(new_n477), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT95), .ZN(new_n497));
  INV_X1    g296(.A(new_n475), .ZN(new_n498));
  XNOR2_X1  g297(.A(KEYINPUT93), .B(G50gat), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n498), .B1(new_n499), .B2(new_n473), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT94), .B1(new_n500), .B2(KEYINPUT15), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n496), .A2(new_n497), .A3(new_n490), .A4(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n493), .A2(new_n494), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT17), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT17), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n493), .A2(new_n505), .A3(new_n502), .A4(new_n494), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(G8gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(G15gat), .B(G22gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT16), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n509), .B1(new_n510), .B2(G1gat), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n508), .B1(new_n511), .B2(KEYINPUT96), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n511), .B1(G1gat), .B2(new_n509), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n507), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(G229gat), .A2(G233gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n503), .A2(new_n514), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n516), .A2(KEYINPUT18), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT97), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT18), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n503), .B(new_n514), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n517), .B(KEYINPUT13), .Z(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n518), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n528), .B1(new_n507), .B2(new_n515), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n529), .A2(KEYINPUT97), .A3(KEYINPUT18), .A4(new_n517), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n521), .A2(new_n524), .A3(new_n527), .A4(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G113gat), .B(G141gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G169gat), .B(G197gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n536), .B(KEYINPUT12), .Z(new_n537));
  NAND2_X1  g336(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n522), .A2(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n539));
  INV_X1    g338(.A(new_n537), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n539), .A2(new_n521), .A3(new_n530), .A4(new_n540), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n538), .A2(KEYINPUT98), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT98), .B1(new_n538), .B2(new_n541), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G85gat), .A2(G92gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT7), .ZN(new_n547));
  NAND2_X1  g346(.A1(G99gat), .A2(G106gat), .ZN(new_n548));
  INV_X1    g347(.A(G85gat), .ZN(new_n549));
  AOI22_X1  g348(.A1(KEYINPUT8), .A2(new_n548), .B1(new_n549), .B2(new_n416), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT104), .ZN(new_n552));
  OR2_X1    g351(.A1(G99gat), .A2(G106gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(new_n548), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n552), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n553), .A2(KEYINPUT104), .A3(new_n548), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n556), .A2(new_n547), .A3(new_n557), .A4(new_n550), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n559), .B1(new_n504), .B2(new_n506), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n503), .A2(new_n559), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT41), .ZN(new_n562));
  NAND2_X1  g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G134gat), .B(G162gat), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n565), .B(KEYINPUT103), .Z(new_n566));
  NOR3_X1   g365(.A1(new_n560), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n563), .A2(new_n562), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT102), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(new_n278), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(G218gat), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n566), .B1(new_n560), .B2(new_n564), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n568), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n572), .B1(new_n568), .B2(new_n573), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G127gat), .B(G155gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(new_n230), .ZN(new_n578));
  INV_X1    g377(.A(G71gat), .ZN(new_n579));
  INV_X1    g378(.A(G78gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G71gat), .A2(G78gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G57gat), .B(G64gat), .Z(new_n584));
  AOI21_X1  g383(.A(new_n583), .B1(new_n584), .B2(KEYINPUT9), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT99), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n587), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n588), .A2(new_n584), .A3(new_n583), .A4(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT100), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI22_X1  g391(.A1(new_n582), .A2(new_n581), .B1(new_n586), .B2(new_n587), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n593), .A2(new_n588), .A3(KEYINPUT100), .A4(new_n584), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n585), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT21), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(G183gat), .B1(new_n597), .B2(new_n514), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n515), .A2(new_n307), .A3(new_n596), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(KEYINPUT101), .ZN(new_n601));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT101), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n598), .A2(new_n599), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n601), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n603), .B1(new_n601), .B2(new_n605), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n578), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n601), .A2(new_n605), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n602), .ZN(new_n611));
  INV_X1    g410(.A(new_n578), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(new_n606), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n592), .A2(new_n594), .ZN(new_n614));
  INV_X1    g413(.A(new_n585), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT21), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n618), .B(new_n619), .Z(new_n620));
  NAND3_X1  g419(.A1(new_n609), .A2(new_n613), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n620), .B1(new_n609), .B2(new_n613), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n576), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G120gat), .B(G148gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(new_n295), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n626), .B(G204gat), .Z(new_n627));
  NAND2_X1  g426(.A1(G230gat), .A2(G233gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT106), .ZN(new_n629));
  XNOR2_X1  g428(.A(KEYINPUT105), .B(KEYINPUT10), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n555), .A2(new_n558), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n631), .A2(new_n595), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n595), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n595), .A2(KEYINPUT10), .A3(new_n559), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n629), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n629), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n632), .A2(new_n633), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n627), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n630), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n616), .A2(new_n559), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n631), .A2(new_n595), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n640), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n635), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n637), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n638), .ZN(new_n646));
  INV_X1    g445(.A(new_n627), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n639), .A2(KEYINPUT107), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT107), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n650), .B(new_n627), .C1(new_n636), .C2(new_n638), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n624), .A2(new_n652), .ZN(new_n653));
  AND3_X1   g452(.A1(new_n468), .A2(new_n545), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n402), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g456(.A(KEYINPUT108), .B(G8gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(new_n510), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n654), .A2(new_n442), .A3(new_n659), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n660), .A2(KEYINPUT42), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n660), .A2(KEYINPUT42), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n654), .A2(new_n442), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n663), .A2(KEYINPUT109), .A3(G8gat), .ZN(new_n664));
  AOI21_X1  g463(.A(KEYINPUT109), .B1(new_n663), .B2(G8gat), .ZN(new_n665));
  OAI22_X1  g464(.A1(new_n661), .A2(new_n662), .B1(new_n664), .B2(new_n665), .ZN(G1325gat));
  AOI21_X1  g465(.A(G15gat), .B1(new_n654), .B2(new_n432), .ZN(new_n667));
  INV_X1    g466(.A(new_n466), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n654), .A2(G15gat), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(G1326gat));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n458), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT43), .B(G22gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1327gat));
  AOI21_X1  g472(.A(new_n576), .B1(new_n434), .B2(new_n467), .ZN(new_n674));
  INV_X1    g473(.A(new_n623), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n621), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n652), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n674), .A2(new_n545), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(G29gat), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n678), .A2(new_n679), .A3(new_n655), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT45), .ZN(new_n681));
  INV_X1    g480(.A(new_n576), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n468), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n538), .A2(new_n541), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n674), .A2(KEYINPUT44), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n685), .A2(new_n686), .A3(new_n677), .A4(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(G29gat), .B1(new_n688), .B2(new_n402), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n681), .A2(new_n689), .ZN(G1328gat));
  NOR2_X1   g489(.A1(new_n423), .A2(G36gat), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n674), .A2(new_n545), .A3(new_n677), .A4(new_n691), .ZN(new_n692));
  XOR2_X1   g491(.A(new_n692), .B(KEYINPUT46), .Z(new_n693));
  OAI21_X1  g492(.A(G36gat), .B1(new_n688), .B2(new_n423), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT110), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n693), .A2(new_n694), .A3(KEYINPUT110), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(G1329gat));
  NOR3_X1   g498(.A1(new_n688), .A2(new_n473), .A3(new_n466), .ZN(new_n700));
  AOI21_X1  g499(.A(G43gat), .B1(new_n678), .B2(new_n432), .ZN(new_n701));
  OR3_X1    g500(.A1(new_n700), .A2(KEYINPUT47), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(KEYINPUT47), .B1(new_n700), .B2(new_n701), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(G1330gat));
  INV_X1    g503(.A(new_n499), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n688), .A2(new_n705), .A3(new_n257), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n499), .B1(new_n678), .B2(new_n458), .ZN(new_n707));
  OR3_X1    g506(.A1(new_n706), .A2(KEYINPUT48), .A3(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT48), .B1(new_n706), .B2(new_n707), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(G1331gat));
  INV_X1    g509(.A(new_n652), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n434), .B2(new_n467), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n624), .A2(new_n686), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n402), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT111), .B(G57gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1332gat));
  NOR2_X1   g516(.A1(new_n714), .A2(new_n423), .ZN(new_n718));
  NOR2_X1   g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  AND2_X1   g518(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(new_n718), .B2(new_n719), .ZN(G1333gat));
  INV_X1    g521(.A(new_n432), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n579), .B1(new_n714), .B2(new_n723), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n712), .A2(G71gat), .A3(new_n668), .A4(new_n713), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g526(.A1(new_n714), .A2(new_n257), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(new_n580), .ZN(G1335gat));
  XNOR2_X1  g528(.A(new_n674), .B(new_n684), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n676), .A2(new_n686), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n652), .ZN(new_n732));
  XOR2_X1   g531(.A(new_n732), .B(KEYINPUT112), .Z(new_n733));
  NAND2_X1  g532(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n734), .A2(new_n549), .A3(new_n402), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n674), .A2(new_n731), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT51), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n674), .A2(KEYINPUT51), .A3(new_n731), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n711), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(G85gat), .B1(new_n740), .B2(new_n655), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n735), .A2(new_n741), .ZN(G1336gat));
  NOR2_X1   g541(.A1(new_n423), .A2(G92gat), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n685), .A2(new_n442), .A3(new_n687), .A4(new_n733), .ZN(new_n744));
  AOI22_X1  g543(.A1(new_n740), .A2(new_n743), .B1(new_n744), .B2(G92gat), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n746), .B1(new_n744), .B2(G92gat), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n745), .A2(KEYINPUT52), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n744), .A2(G92gat), .ZN(new_n749));
  INV_X1    g548(.A(new_n739), .ZN(new_n750));
  AOI21_X1  g549(.A(KEYINPUT51), .B1(new_n674), .B2(new_n731), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n652), .B(new_n743), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n749), .B(new_n752), .C1(KEYINPUT113), .C2(KEYINPUT52), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n748), .A2(new_n754), .ZN(G1337gat));
  OAI21_X1  g554(.A(G99gat), .B1(new_n734), .B2(new_n466), .ZN(new_n756));
  INV_X1    g555(.A(G99gat), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n757), .A3(new_n432), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(G1338gat));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n685), .A2(new_n458), .A3(new_n687), .A4(new_n733), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n760), .B1(new_n761), .B2(G106gat), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n257), .A2(G106gat), .A3(new_n711), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT114), .Z(new_n764));
  OAI21_X1  g563(.A(new_n764), .B1(new_n750), .B2(new_n751), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n730), .A2(KEYINPUT115), .A3(new_n458), .A4(new_n733), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n761), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n767), .A2(new_n769), .A3(G106gat), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n763), .B1(new_n750), .B2(new_n751), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n766), .B1(new_n772), .B2(new_n760), .ZN(G1339gat));
  NAND2_X1  g572(.A1(new_n655), .A2(new_n423), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT54), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n647), .B1(new_n636), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n634), .A2(new_n629), .A3(new_n635), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n645), .A2(new_n777), .A3(KEYINPUT54), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n776), .A2(KEYINPUT55), .A3(new_n778), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(new_n648), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n783), .B1(new_n538), .B2(new_n541), .ZN(new_n784));
  OAI22_X1  g583(.A1(new_n529), .A2(new_n517), .B1(new_n525), .B2(new_n526), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n536), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n541), .A2(new_n652), .A3(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n576), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n541), .A2(new_n786), .ZN(new_n789));
  INV_X1    g588(.A(new_n783), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(new_n682), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n676), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n624), .A2(new_n686), .A3(new_n652), .ZN(new_n794));
  INV_X1    g593(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n774), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  AND3_X1   g595(.A1(new_n257), .A2(new_n350), .A3(new_n355), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n799), .A2(new_n262), .A3(new_n686), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n458), .A2(new_n723), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n796), .A2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(G113gat), .B1(new_n802), .B2(new_n544), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n800), .A2(new_n803), .ZN(G1340gat));
  OAI21_X1  g603(.A(G120gat), .B1(new_n802), .B2(new_n711), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n652), .A2(new_n260), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n805), .B1(new_n798), .B2(new_n806), .ZN(G1341gat));
  INV_X1    g606(.A(new_n676), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n802), .A2(new_n267), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n799), .A2(new_n676), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n809), .B1(new_n267), .B2(new_n810), .ZN(G1342gat));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n682), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(new_n269), .A3(new_n797), .ZN(new_n814));
  XOR2_X1   g613(.A(new_n814), .B(KEYINPUT56), .Z(new_n815));
  AOI21_X1  g614(.A(new_n269), .B1(new_n813), .B2(new_n801), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(KEYINPUT116), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(G1343gat));
  NOR2_X1   g617(.A1(new_n668), .A2(new_n774), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n458), .B1(new_n792), .B2(new_n794), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(G141gat), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n823), .A3(new_n545), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n790), .B1(new_n542), .B2(new_n543), .ZN(new_n828));
  INV_X1    g627(.A(new_n787), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n682), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n791), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n808), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n827), .B1(new_n832), .B2(new_n795), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n833), .A2(new_n458), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n821), .A2(new_n827), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n826), .B(new_n819), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  AOI22_X1  g635(.A1(new_n833), .A2(new_n458), .B1(new_n827), .B2(new_n821), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT117), .B1(new_n837), .B2(new_n820), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n686), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n825), .B1(new_n840), .B2(G141gat), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n837), .A2(new_n544), .A3(new_n820), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n842), .B1(new_n843), .B2(new_n823), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n824), .B(KEYINPUT118), .ZN(new_n845));
  OAI22_X1  g644(.A1(new_n841), .A2(new_n842), .B1(new_n844), .B2(new_n845), .ZN(G1344gat));
  NAND2_X1  g645(.A1(new_n653), .A2(new_n544), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n257), .A2(KEYINPUT57), .ZN(new_n849));
  AOI22_X1  g648(.A1(new_n848), .A2(new_n849), .B1(KEYINPUT57), .B2(new_n821), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n850), .A2(KEYINPUT59), .A3(new_n652), .A4(new_n819), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n711), .B1(new_n836), .B2(new_n838), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n852), .B2(KEYINPUT59), .ZN(new_n853));
  AOI21_X1  g652(.A(G148gat), .B1(new_n822), .B2(new_n652), .ZN(new_n854));
  AOI22_X1  g653(.A1(new_n853), .A2(G148gat), .B1(KEYINPUT59), .B2(new_n854), .ZN(G1345gat));
  AOI21_X1  g654(.A(G155gat), .B1(new_n822), .B2(new_n676), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n808), .B1(new_n836), .B2(new_n838), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n857), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g657(.A(G162gat), .B1(new_n822), .B2(new_n682), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n576), .B1(new_n836), .B2(new_n838), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n859), .B1(new_n860), .B2(G162gat), .ZN(G1347gat));
  OAI21_X1  g660(.A(new_n402), .B1(new_n792), .B2(new_n794), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(new_n801), .A3(new_n442), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(KEYINPUT120), .ZN(new_n865));
  OAI21_X1  g664(.A(G169gat), .B1(new_n865), .B2(new_n544), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n862), .A2(KEYINPUT119), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT119), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n868), .B(new_n402), .C1(new_n792), .C2(new_n794), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(new_n442), .A3(new_n797), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(new_n294), .A3(new_n686), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n866), .A2(new_n873), .ZN(G1348gat));
  XOR2_X1   g673(.A(new_n864), .B(KEYINPUT120), .Z(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(G176gat), .A3(new_n652), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n295), .B1(new_n871), .B2(new_n711), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(KEYINPUT121), .ZN(G1349gat));
  OAI21_X1  g678(.A(G183gat), .B1(new_n865), .B2(new_n808), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n676), .A2(new_n277), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n871), .B2(new_n881), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g682(.A1(new_n872), .A2(new_n278), .A3(new_n682), .ZN(new_n884));
  OAI21_X1  g683(.A(G190gat), .B1(new_n865), .B2(new_n576), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n885), .A2(KEYINPUT61), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n885), .A2(KEYINPUT61), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n884), .B1(new_n886), .B2(new_n887), .ZN(G1351gat));
  AND3_X1   g687(.A1(new_n466), .A2(new_n458), .A3(new_n442), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n870), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(G197gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n891), .A2(new_n892), .A3(new_n686), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n668), .A2(new_n655), .A3(new_n423), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n850), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G197gat), .B1(new_n895), .B2(new_n544), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n893), .A2(new_n896), .ZN(G1352gat));
  NOR2_X1   g696(.A1(new_n711), .A2(G204gat), .ZN(new_n898));
  AND4_X1   g697(.A1(new_n867), .A2(new_n869), .A3(new_n889), .A4(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT122), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n867), .A2(new_n889), .A3(new_n869), .A4(new_n898), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT122), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT123), .B1(new_n904), .B2(KEYINPUT62), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n907));
  AOI211_X1 g706(.A(new_n906), .B(new_n907), .C1(new_n901), .C2(new_n903), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n850), .A2(new_n652), .A3(new_n894), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT124), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n850), .A2(new_n912), .A3(new_n652), .A4(new_n894), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n911), .A2(G204gat), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n902), .B(new_n900), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n907), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT125), .B1(new_n909), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n906), .B1(new_n915), .B2(new_n907), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n904), .A2(KEYINPUT123), .A3(KEYINPUT62), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n921), .A2(new_n922), .A3(new_n916), .A4(new_n914), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n918), .A2(new_n923), .ZN(G1353gat));
  NOR2_X1   g723(.A1(new_n895), .A2(new_n808), .ZN(new_n925));
  NOR2_X1   g724(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n925), .A2(new_n230), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n891), .A2(new_n230), .A3(new_n676), .ZN(new_n930));
  OAI211_X1 g729(.A(KEYINPUT126), .B(KEYINPUT63), .C1(new_n925), .C2(new_n230), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(G1354gat));
  NOR3_X1   g731(.A1(new_n895), .A2(new_n231), .A3(new_n576), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n231), .B1(new_n890), .B2(new_n576), .ZN(new_n934));
  OR2_X1    g733(.A1(new_n934), .A2(KEYINPUT127), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(KEYINPUT127), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(G1355gat));
endmodule


