//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n806, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT28), .ZN(new_n205));
  NOR2_X1   g004(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(KEYINPUT66), .B(G183gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n206), .B1(new_n207), .B2(KEYINPUT27), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n205), .B1(new_n208), .B2(G190gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT27), .B(G183gat), .ZN(new_n210));
  INV_X1    g009(.A(G190gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(KEYINPUT28), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G169gat), .ZN(new_n214));
  INV_X1    g013(.A(G176gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n214), .A2(new_n215), .ZN(new_n218));
  NOR3_X1   g017(.A1(new_n217), .A2(new_n218), .A3(KEYINPUT26), .ZN(new_n219));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT26), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n220), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n213), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n216), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT64), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT24), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n220), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n229), .B(new_n230), .C1(G183gat), .C2(G190gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT64), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(new_n216), .B2(new_n225), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n216), .B1(new_n218), .B2(new_n225), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n227), .A2(new_n231), .A3(new_n233), .A4(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT25), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n226), .A2(new_n236), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n230), .B1(new_n207), .B2(G190gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n220), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n242));
  NOR3_X1   g041(.A1(new_n241), .A2(KEYINPUT24), .A3(new_n242), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n234), .B(new_n238), .C1(new_n239), .C2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n237), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n224), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n247));
  NAND2_X1  g046(.A1(G113gat), .A2(G120gat), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NOR2_X1   g048(.A1(G113gat), .A2(G120gat), .ZN(new_n250));
  NOR3_X1   g049(.A1(new_n249), .A2(new_n250), .A3(KEYINPUT1), .ZN(new_n251));
  XNOR2_X1  g050(.A(G127gat), .B(G134gat), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n247), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n250), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(KEYINPUT68), .A3(new_n248), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n256), .B1(new_n249), .B2(new_n250), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT1), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n255), .A2(new_n257), .A3(new_n258), .A4(new_n252), .ZN(new_n259));
  INV_X1    g058(.A(new_n252), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n254), .A2(new_n258), .A3(new_n248), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT67), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n253), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n263), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n213), .A2(new_n223), .B1(new_n237), .B2(new_n244), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n253), .A2(new_n259), .A3(new_n262), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(G227gat), .ZN(new_n268));
  INV_X1    g067(.A(G233gat), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n264), .A2(new_n267), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n204), .B1(new_n271), .B2(KEYINPUT32), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT33), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n204), .A2(KEYINPUT69), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n204), .A2(KEYINPUT69), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(KEYINPUT33), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n271), .A2(KEYINPUT32), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT34), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n267), .ZN(new_n282));
  INV_X1    g081(.A(new_n270), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AOI211_X1 g083(.A(KEYINPUT34), .B(new_n270), .C1(new_n264), .C2(new_n267), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n275), .A3(new_n279), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(KEYINPUT70), .B1(new_n275), .B2(new_n279), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(new_n286), .ZN(new_n292));
  MUX2_X1   g091(.A(new_n290), .B(new_n292), .S(KEYINPUT36), .Z(new_n293));
  INV_X1    g092(.A(KEYINPUT4), .ZN(new_n294));
  INV_X1    g093(.A(G141gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G148gat), .ZN(new_n296));
  INV_X1    g095(.A(G148gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G141gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n296), .A2(new_n298), .B1(KEYINPUT2), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(G155gat), .B(G162gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n299), .ZN(new_n303));
  INV_X1    g102(.A(G155gat), .ZN(new_n304));
  INV_X1    g103(.A(G162gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(new_n305), .A3(KEYINPUT74), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(G155gat), .B2(G162gat), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n303), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n299), .A2(KEYINPUT2), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n297), .A2(G141gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n295), .A2(G148gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  AND3_X1   g112(.A1(new_n309), .A2(new_n313), .A3(KEYINPUT75), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT75), .B1(new_n309), .B2(new_n313), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n302), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n294), .B1(new_n316), .B2(new_n266), .ZN(new_n317));
  INV_X1    g116(.A(new_n302), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT75), .ZN(new_n319));
  NOR3_X1   g118(.A1(new_n307), .A2(G155gat), .A3(G162gat), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT74), .B1(new_n304), .B2(new_n305), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n299), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n319), .B1(new_n322), .B2(new_n300), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n309), .A2(new_n313), .A3(KEYINPUT75), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n318), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n325), .A2(new_n263), .A3(KEYINPUT4), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n266), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  AOI211_X1 g127(.A(KEYINPUT3), .B(new_n318), .C1(new_n323), .C2(new_n324), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n317), .B(new_n326), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G225gat), .A2(G233gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT76), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n317), .A2(new_n326), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT76), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n316), .A2(KEYINPUT3), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n325), .A2(new_n327), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n337), .A3(new_n266), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n334), .A2(new_n335), .A3(new_n331), .A4(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n333), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n325), .A2(new_n263), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n316), .A2(new_n266), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n332), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT5), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n347));
  XNOR2_X1  g146(.A(G1gat), .B(G29gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(G57gat), .B(G85gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n338), .A2(new_n331), .A3(new_n317), .A4(new_n326), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n352), .B1(new_n353), .B2(KEYINPUT5), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n346), .A2(new_n347), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n352), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n344), .B1(new_n333), .B2(new_n339), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n353), .A2(KEYINPUT5), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT78), .B1(new_n358), .B2(new_n354), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT6), .ZN(new_n362));
  NAND4_X1  g161(.A1(new_n356), .A2(new_n360), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  OAI211_X1 g162(.A(KEYINPUT6), .B(new_n357), .C1(new_n358), .C2(new_n359), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(G226gat), .ZN(new_n366));
  OAI22_X1  g165(.A1(new_n265), .A2(KEYINPUT29), .B1(new_n366), .B2(new_n269), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n246), .A2(G226gat), .A3(G233gat), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT72), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT22), .ZN(new_n370));
  XOR2_X1   g169(.A(KEYINPUT71), .B(G211gat), .Z(new_n371));
  INV_X1    g170(.A(G218gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G197gat), .B(G204gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(G211gat), .B(G218gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n375), .B1(new_n373), .B2(new_n374), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n369), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n378), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(KEYINPUT72), .A3(new_n376), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n367), .A2(new_n368), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n382), .B1(new_n367), .B2(new_n368), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n384), .A2(KEYINPUT37), .A3(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G8gat), .B(G36gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(G64gat), .B(G92gat), .ZN(new_n388));
  XOR2_X1   g187(.A(new_n387), .B(new_n388), .Z(new_n389));
  OR2_X1    g188(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n384), .A2(new_n385), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT37), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(KEYINPUT38), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n389), .ZN(new_n395));
  NOR3_X1   g194(.A1(new_n384), .A2(new_n385), .A3(new_n395), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n385), .A2(KEYINPUT86), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n383), .A2(KEYINPUT85), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n385), .A2(KEYINPUT86), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n383), .A2(KEYINPUT85), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n397), .A2(new_n398), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT37), .ZN(new_n402));
  XOR2_X1   g201(.A(new_n389), .B(KEYINPUT73), .Z(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n386), .A2(KEYINPUT38), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n396), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n365), .A2(new_n394), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(G228gat), .A2(G233gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT29), .B1(new_n380), .B2(new_n376), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n316), .B1(new_n410), .B2(KEYINPUT3), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n379), .B(new_n381), .C1(new_n329), .C2(KEYINPUT29), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n409), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(G22gat), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n411), .A2(new_n412), .A3(new_n409), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT82), .ZN(new_n418));
  XOR2_X1   g217(.A(KEYINPUT31), .B(G50gat), .Z(new_n419));
  XNOR2_X1  g218(.A(new_n419), .B(KEYINPUT81), .ZN(new_n420));
  XOR2_X1   g219(.A(G78gat), .B(G106gat), .Z(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n416), .ZN(new_n423));
  OAI21_X1  g222(.A(G22gat), .B1(new_n423), .B2(new_n413), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n418), .A2(new_n422), .B1(new_n417), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT82), .ZN(new_n426));
  AND4_X1   g225(.A1(new_n426), .A2(new_n417), .A3(new_n424), .A4(new_n422), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n385), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n404), .B1(new_n429), .B2(new_n383), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT30), .B1(new_n430), .B2(new_n396), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n391), .A2(new_n389), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT30), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n341), .A2(new_n342), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT39), .B1(new_n436), .B2(new_n332), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n331), .B1(new_n334), .B2(new_n338), .ZN(new_n438));
  OR2_X1    g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT39), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n357), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT40), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT83), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n442), .A2(new_n443), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n435), .B(new_n360), .C1(new_n444), .C2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n439), .A2(KEYINPUT40), .A3(new_n441), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT84), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n428), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n293), .B1(new_n407), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n428), .ZN(new_n452));
  INV_X1    g251(.A(new_n364), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT79), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n453), .B1(new_n363), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n354), .B1(new_n340), .B2(new_n345), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT6), .B1(new_n456), .B2(new_n347), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n457), .A2(KEYINPUT79), .A3(new_n360), .A4(new_n361), .ZN(new_n458));
  AOI211_X1 g257(.A(KEYINPUT80), .B(new_n435), .C1(new_n455), .C2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT80), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n363), .A2(new_n454), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n461), .A2(new_n458), .A3(new_n364), .ZN(new_n462));
  INV_X1    g261(.A(new_n435), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n452), .B1(new_n459), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n451), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT35), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n459), .A2(new_n464), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT87), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n292), .A2(new_n428), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n469), .B1(new_n292), .B2(new_n428), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n467), .B1(new_n468), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n290), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n463), .A2(new_n474), .ZN(new_n475));
  NOR4_X1   g274(.A1(new_n452), .A2(new_n475), .A3(new_n365), .A4(KEYINPUT35), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n466), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G15gat), .B(G22gat), .ZN(new_n478));
  INV_X1    g277(.A(G1gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT16), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n481), .B1(G1gat), .B2(new_n478), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(G8gat), .ZN(new_n483));
  INV_X1    g282(.A(G8gat), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n481), .B(new_n484), .C1(G1gat), .C2(new_n478), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G43gat), .B(G50gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(KEYINPUT88), .B(G36gat), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n491), .A2(G29gat), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NOR3_X1   g293(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n490), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n491), .A2(G29gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n498), .A2(new_n499), .A3(new_n489), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n495), .A2(KEYINPUT89), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n495), .A2(KEYINPUT89), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n494), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n497), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n504), .A2(KEYINPUT17), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT17), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n497), .B(new_n506), .C1(new_n500), .C2(new_n503), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n487), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n504), .A2(new_n486), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT90), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT90), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n504), .A2(new_n486), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(G229gat), .A2(G233gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n509), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT18), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XOR2_X1   g317(.A(new_n515), .B(KEYINPUT13), .Z(new_n519));
  AND3_X1   g318(.A1(new_n504), .A2(new_n486), .A3(new_n512), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n512), .B1(new_n504), .B2(new_n486), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n504), .A2(new_n486), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n509), .A2(new_n514), .A3(KEYINPUT18), .A4(new_n515), .ZN(new_n525));
  XNOR2_X1  g324(.A(G113gat), .B(G141gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(G197gat), .ZN(new_n527));
  XOR2_X1   g326(.A(KEYINPUT11), .B(G169gat), .Z(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT12), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n518), .A2(new_n524), .A3(new_n525), .A4(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n530), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n525), .A2(new_n524), .A3(KEYINPUT91), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n518), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT91), .B1(new_n525), .B2(new_n524), .ZN(new_n535));
  OAI211_X1 g334(.A(KEYINPUT92), .B(new_n532), .C1(new_n534), .C2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n525), .A2(new_n524), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT91), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(new_n518), .A3(new_n533), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT92), .B1(new_n541), .B2(new_n532), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n531), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  XOR2_X1   g342(.A(G57gat), .B(G64gat), .Z(new_n544));
  INV_X1    g343(.A(KEYINPUT9), .ZN(new_n545));
  INV_X1    g344(.A(G71gat), .ZN(new_n546));
  INV_X1    g345(.A(G78gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G71gat), .B(G78gat), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT93), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n544), .A2(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n551), .B1(new_n550), .B2(new_n549), .ZN(new_n552));
  INV_X1    g351(.A(new_n549), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n553), .A2(new_n544), .A3(KEYINPUT93), .A4(new_n548), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n555), .A2(KEYINPUT21), .ZN(new_n556));
  NAND2_X1  g355(.A1(G231gat), .A2(G233gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G127gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n486), .B1(new_n555), .B2(KEYINPUT21), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(new_n304), .ZN(new_n564));
  XOR2_X1   g363(.A(G183gat), .B(G211gat), .Z(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  OR2_X1    g365(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n562), .A2(new_n566), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(KEYINPUT95), .A2(G85gat), .A3(G92gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(KEYINPUT7), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT7), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(KEYINPUT94), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n571), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(G99gat), .ZN(new_n575));
  INV_X1    g374(.A(G106gat), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT8), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(G85gat), .ZN(new_n578));
  INV_X1    g377(.A(G92gat), .ZN(new_n579));
  OAI21_X1  g378(.A(KEYINPUT94), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n578), .A2(new_n579), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n574), .A2(new_n577), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G99gat), .B(G106gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  AND2_X1   g383(.A1(G232gat), .A2(G233gat), .ZN(new_n585));
  AOI22_X1  g384(.A1(new_n584), .A2(new_n504), .B1(KEYINPUT41), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n505), .A2(new_n508), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n586), .B1(new_n587), .B2(new_n584), .ZN(new_n588));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n585), .A2(KEYINPUT41), .ZN(new_n591));
  XNOR2_X1  g390(.A(G134gat), .B(G162gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n590), .A2(new_n593), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n569), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G230gat), .A2(G233gat), .ZN(new_n598));
  XOR2_X1   g397(.A(KEYINPUT97), .B(KEYINPUT10), .Z(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  AND2_X1   g399(.A1(new_n552), .A2(new_n554), .ZN(new_n601));
  INV_X1    g400(.A(new_n582), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n602), .A2(new_n583), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n583), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n584), .A2(new_n555), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n605), .A2(KEYINPUT96), .A3(new_n606), .ZN(new_n607));
  OR3_X1    g406(.A1(new_n584), .A2(KEYINPUT96), .A3(new_n555), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n600), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n606), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT10), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n598), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n598), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n607), .A2(new_n614), .A3(new_n608), .ZN(new_n615));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(G176gat), .B(G204gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n616), .B(new_n617), .Z(new_n618));
  AND3_X1   g417(.A1(new_n613), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n618), .B1(new_n613), .B2(new_n615), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n597), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n623), .B(KEYINPUT98), .Z(new_n624));
  AND3_X1   g423(.A1(new_n477), .A2(new_n543), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n462), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(G1gat), .ZN(G1324gat));
  XNOR2_X1  g427(.A(KEYINPUT99), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(G8gat), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n625), .A2(new_n435), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n484), .B1(new_n625), .B2(new_n435), .ZN(new_n632));
  OAI21_X1  g431(.A(KEYINPUT42), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(KEYINPUT42), .B2(new_n631), .ZN(G1325gat));
  INV_X1    g433(.A(G15gat), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n625), .A2(new_n635), .A3(new_n474), .ZN(new_n636));
  INV_X1    g435(.A(new_n293), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n625), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n636), .B1(new_n639), .B2(new_n635), .ZN(G1326gat));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n452), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT43), .B(G22gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(G1327gat));
  INV_X1    g442(.A(new_n596), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n462), .A2(new_n463), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT80), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n462), .A2(new_n460), .A3(new_n463), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n646), .A2(new_n472), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n476), .B1(new_n648), .B2(KEYINPUT35), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n647), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n450), .B1(new_n650), .B2(new_n452), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n644), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n543), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n654), .A2(new_n569), .A3(new_n622), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n656), .A2(G29gat), .A3(new_n462), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT100), .B(KEYINPUT45), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n652), .A2(new_n660), .ZN(new_n661));
  OAI211_X1 g460(.A(KEYINPUT44), .B(new_n644), .C1(new_n649), .C2(new_n651), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n655), .B(KEYINPUT101), .Z(new_n663));
  NAND3_X1  g462(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(G29gat), .B1(new_n664), .B2(new_n462), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n659), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n659), .A2(new_n665), .A3(KEYINPUT102), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(G1328gat));
  NOR3_X1   g469(.A1(new_n656), .A2(new_n463), .A3(new_n491), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT46), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n491), .B1(new_n664), .B2(new_n463), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(G1329gat));
  OAI21_X1  g473(.A(G43gat), .B1(new_n664), .B2(new_n293), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n290), .A2(G43gat), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n675), .B1(new_n656), .B2(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g477(.A(G50gat), .B1(new_n664), .B2(new_n428), .ZN(new_n679));
  INV_X1    g478(.A(new_n656), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT103), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n428), .A2(G50gat), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT104), .Z(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n680), .A2(KEYINPUT103), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n679), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT48), .Z(G1331gat));
  NOR3_X1   g486(.A1(new_n597), .A2(new_n543), .A3(new_n621), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n477), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n626), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n435), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT49), .B(G64gat), .Z(new_n694));
  OAI21_X1  g493(.A(new_n693), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT105), .ZN(G1333gat));
  AOI21_X1  g495(.A(new_n546), .B1(new_n689), .B2(new_n637), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n290), .A2(G71gat), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n697), .B1(new_n689), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g499(.A1(new_n689), .A2(new_n452), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g501(.A1(new_n569), .A2(new_n543), .A3(new_n621), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n661), .A2(new_n662), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(KEYINPUT106), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n661), .A2(new_n706), .A3(new_n662), .A4(new_n703), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n705), .A2(new_n626), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n569), .A2(new_n543), .ZN(new_n709));
  OAI211_X1 g508(.A(new_n644), .B(new_n709), .C1(new_n649), .C2(new_n651), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT51), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n477), .A2(KEYINPUT51), .A3(new_n644), .A4(new_n709), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n622), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n626), .A2(new_n578), .ZN(new_n716));
  OAI22_X1  g515(.A1(new_n708), .A2(new_n578), .B1(new_n715), .B2(new_n716), .ZN(G1336gat));
  OAI21_X1  g516(.A(G92gat), .B1(new_n704), .B2(new_n463), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT52), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n463), .A2(G92gat), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n718), .B(new_n719), .C1(new_n715), .C2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n705), .A2(new_n435), .A3(new_n707), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G92gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n712), .A2(new_n713), .A3(KEYINPUT107), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n710), .A2(new_n727), .A3(new_n711), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n721), .A2(new_n621), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n726), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n725), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n723), .B1(new_n732), .B2(KEYINPUT52), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n730), .B1(new_n724), .B2(G92gat), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n734), .A2(KEYINPUT108), .A3(new_n719), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n722), .B1(new_n733), .B2(new_n735), .ZN(G1337gat));
  AND3_X1   g535(.A1(new_n705), .A2(new_n637), .A3(new_n707), .ZN(new_n737));
  INV_X1    g536(.A(new_n714), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n474), .A2(new_n622), .A3(new_n575), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT109), .ZN(new_n740));
  OAI22_X1  g539(.A1(new_n737), .A2(new_n575), .B1(new_n738), .B2(new_n740), .ZN(G1338gat));
  NOR3_X1   g540(.A1(new_n428), .A2(new_n621), .A3(G106gat), .ZN(new_n742));
  AND3_X1   g541(.A1(new_n726), .A2(new_n728), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n705), .A2(new_n452), .A3(new_n707), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n743), .B1(new_n744), .B2(G106gat), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT53), .ZN(new_n746));
  INV_X1    g545(.A(new_n704), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n576), .B1(new_n747), .B2(new_n452), .ZN(new_n748));
  INV_X1    g547(.A(new_n742), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n746), .B1(new_n738), .B2(new_n749), .ZN(new_n750));
  OAI22_X1  g549(.A1(new_n745), .A2(new_n746), .B1(new_n748), .B2(new_n750), .ZN(G1339gat));
  NAND2_X1  g550(.A1(new_n607), .A2(new_n608), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n599), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n753), .A2(new_n614), .A3(new_n611), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n754), .A2(KEYINPUT54), .A3(new_n613), .ZN(new_n755));
  XOR2_X1   g554(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n756));
  OAI211_X1 g555(.A(new_n598), .B(new_n756), .C1(new_n609), .C2(new_n612), .ZN(new_n757));
  INV_X1    g556(.A(new_n618), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n619), .B1(new_n760), .B2(KEYINPUT55), .ZN(new_n761));
  OR3_X1    g560(.A1(new_n522), .A2(new_n523), .A3(new_n519), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n515), .B1(new_n509), .B2(new_n514), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n529), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n531), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n596), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n755), .B2(new_n759), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n761), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n621), .A2(new_n766), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(KEYINPUT111), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n621), .B2(new_n766), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n543), .A2(new_n761), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n775), .B1(new_n776), .B2(new_n769), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n770), .B1(new_n777), .B2(new_n644), .ZN(new_n778));
  INV_X1    g577(.A(new_n569), .ZN(new_n779));
  AOI22_X1  g578(.A1(new_n778), .A2(new_n779), .B1(new_n654), .B2(new_n623), .ZN(new_n780));
  NOR4_X1   g579(.A1(new_n780), .A2(new_n462), .A3(new_n471), .A4(new_n470), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n781), .A2(new_n463), .ZN(new_n782));
  AOI21_X1  g581(.A(G113gat), .B1(new_n782), .B2(new_n543), .ZN(new_n783));
  INV_X1    g582(.A(new_n780), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n784), .A2(KEYINPUT112), .A3(new_n428), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT112), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n786), .B1(new_n780), .B2(new_n452), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n462), .A2(new_n475), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n788), .A2(KEYINPUT113), .A3(new_n789), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n543), .A2(G113gat), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n783), .B1(new_n794), .B2(new_n795), .ZN(G1340gat));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n792), .A2(new_n622), .A3(new_n793), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(G120gat), .ZN(new_n799));
  INV_X1    g598(.A(G120gat), .ZN(new_n800));
  AND3_X1   g599(.A1(new_n782), .A2(new_n800), .A3(new_n622), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n797), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  AOI211_X1 g602(.A(KEYINPUT114), .B(new_n801), .C1(new_n798), .C2(G120gat), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n803), .A2(new_n804), .ZN(G1341gat));
  NAND3_X1  g604(.A1(new_n782), .A2(new_n559), .A3(new_n569), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n794), .A2(new_n569), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n806), .B1(new_n807), .B2(new_n559), .ZN(G1342gat));
  NAND2_X1  g607(.A1(new_n794), .A2(new_n644), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G134gat), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n596), .A2(new_n435), .A3(G134gat), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n781), .A2(new_n811), .ZN(new_n812));
  XOR2_X1   g611(.A(KEYINPUT115), .B(KEYINPUT56), .Z(new_n813));
  XNOR2_X1  g612(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n810), .A2(new_n814), .ZN(G1343gat));
  NOR3_X1   g614(.A1(new_n637), .A2(new_n462), .A3(new_n435), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n623), .A2(new_n654), .ZN(new_n817));
  INV_X1    g616(.A(new_n770), .ZN(new_n818));
  OAI21_X1  g617(.A(KEYINPUT116), .B1(new_n755), .B2(new_n759), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n754), .A2(KEYINPUT54), .A3(new_n613), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n820), .A2(new_n821), .A3(new_n758), .A4(new_n757), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(new_n768), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n543), .A2(new_n823), .A3(new_n761), .ZN(new_n824));
  INV_X1    g623(.A(new_n771), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n644), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n824), .A2(KEYINPUT117), .A3(new_n825), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n818), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n817), .B1(new_n830), .B2(new_n569), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n428), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n831), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n780), .B2(new_n428), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n832), .B1(new_n831), .B2(new_n834), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n816), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OR3_X1    g638(.A1(new_n839), .A2(new_n295), .A3(new_n654), .ZN(new_n840));
  NOR4_X1   g639(.A1(new_n780), .A2(new_n462), .A3(new_n428), .A4(new_n637), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(new_n463), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n543), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n295), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT58), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n840), .A2(KEYINPUT58), .A3(new_n844), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(G1344gat));
  NAND3_X1  g648(.A1(new_n842), .A2(new_n297), .A3(new_n622), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT59), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n816), .A2(new_n622), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n624), .A2(new_n654), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n779), .B1(new_n830), .B2(KEYINPUT119), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n855));
  AOI211_X1 g654(.A(new_n855), .B(new_n818), .C1(new_n828), .C2(new_n829), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n853), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT57), .B1(new_n857), .B2(new_n452), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n780), .A2(new_n833), .A3(new_n428), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n852), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n851), .B1(new_n860), .B2(G148gat), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n622), .B(new_n816), .C1(new_n837), .C2(new_n838), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n297), .A2(KEYINPUT59), .ZN(new_n863));
  AND2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n850), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(KEYINPUT120), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n867), .B(new_n850), .C1(new_n861), .C2(new_n864), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n868), .ZN(G1345gat));
  NAND2_X1  g668(.A1(new_n569), .A2(G155gat), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT121), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n839), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(G155gat), .B1(new_n842), .B2(new_n569), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(G1346gat));
  OAI21_X1  g674(.A(G162gat), .B1(new_n839), .B2(new_n596), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n841), .A2(new_n305), .A3(new_n463), .A4(new_n644), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1347gat));
  NAND2_X1  g677(.A1(new_n784), .A2(new_n462), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n463), .B1(new_n879), .B2(KEYINPUT122), .ZN(new_n880));
  OR3_X1    g679(.A1(new_n780), .A2(KEYINPUT122), .A3(new_n626), .ZN(new_n881));
  AND3_X1   g680(.A1(new_n880), .A2(new_n472), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(G169gat), .B1(new_n882), .B2(new_n543), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n626), .A2(new_n463), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n474), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n885), .B1(new_n785), .B2(new_n787), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n654), .A2(new_n214), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n883), .B1(new_n886), .B2(new_n887), .ZN(G1348gat));
  INV_X1    g687(.A(new_n886), .ZN(new_n889));
  OAI21_X1  g688(.A(G176gat), .B1(new_n889), .B2(new_n621), .ZN(new_n890));
  INV_X1    g689(.A(new_n882), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n622), .A2(new_n215), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(G1349gat));
  NAND3_X1  g692(.A1(new_n882), .A2(new_n210), .A3(new_n569), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT123), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n207), .B1(new_n889), .B2(new_n779), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT60), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT60), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n894), .A2(new_n895), .A3(new_n899), .A4(new_n896), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(G1350gat));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n644), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(G190gat), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(KEYINPUT125), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT125), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n902), .A2(new_n905), .A3(G190gat), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n644), .A2(new_n211), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT124), .B1(new_n891), .B2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n882), .A2(new_n912), .A3(new_n211), .A4(new_n644), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n904), .A2(new_n906), .A3(KEYINPUT61), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n909), .A2(new_n914), .A3(new_n915), .ZN(G1351gat));
  AND2_X1   g715(.A1(new_n880), .A2(new_n881), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n637), .A2(new_n428), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(G197gat), .B1(new_n919), .B2(new_n543), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n858), .A2(new_n859), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n884), .A2(new_n293), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n543), .A2(G197gat), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n920), .B1(new_n923), .B2(new_n924), .ZN(G1352gat));
  NOR2_X1   g724(.A1(new_n621), .A2(G204gat), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n917), .A2(new_n918), .A3(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT62), .ZN(new_n928));
  XNOR2_X1  g727(.A(new_n927), .B(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n923), .A2(new_n622), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(G204gat), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1353gat));
  NAND3_X1  g731(.A1(new_n919), .A2(new_n371), .A3(new_n569), .ZN(new_n933));
  NAND2_X1  g732(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n934));
  OAI21_X1  g733(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n935));
  AOI211_X1 g734(.A(new_n934), .B(new_n935), .C1(new_n923), .C2(new_n569), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n858), .A2(new_n859), .ZN(new_n937));
  INV_X1    g736(.A(new_n922), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n937), .A2(new_n569), .A3(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(new_n935), .ZN(new_n940));
  AOI22_X1  g739(.A1(new_n939), .A2(new_n940), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n933), .B1(new_n936), .B2(new_n941), .ZN(G1354gat));
  AOI21_X1  g741(.A(new_n372), .B1(new_n923), .B2(new_n644), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n596), .A2(G218gat), .ZN(new_n944));
  AND3_X1   g743(.A1(new_n917), .A2(new_n918), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(KEYINPUT127), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n937), .A2(new_n644), .A3(new_n938), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(G218gat), .ZN(new_n948));
  INV_X1    g747(.A(new_n945), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT127), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n946), .A2(new_n951), .ZN(G1355gat));
endmodule


