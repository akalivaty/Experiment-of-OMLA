//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1296, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  OAI21_X1  g0011(.A(G50), .B1(G58), .B2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  INV_X1    g0021(.A(G97), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT64), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n217), .B(new_n218), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AND2_X1   g0026(.A1(new_n224), .A2(new_n225), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n208), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XOR2_X1   g0030(.A(G238), .B(G244), .Z(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(KEYINPUT3), .ZN(new_n247));
  INV_X1    g0047(.A(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G1698), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n251), .A2(G222), .A3(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G77), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n251), .A2(G1698), .ZN(new_n255));
  INV_X1    g0055(.A(G223), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n253), .B1(new_n254), .B2(new_n251), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n214), .B1(G33), .B2(G41), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  INV_X1    g0060(.A(new_n214), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G41), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  INV_X1    g0068(.A(G45), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n205), .A2(new_n270), .B1(new_n261), .B2(new_n262), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n267), .B1(G226), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n259), .A2(KEYINPUT66), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(KEYINPUT66), .B1(new_n259), .B2(new_n272), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G169), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n214), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G13), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G1), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G20), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n281), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(KEYINPUT68), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n282), .A2(new_n206), .A3(G1), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n280), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT68), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n286), .A2(new_n290), .B1(new_n205), .B2(G20), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G50), .ZN(new_n292));
  XNOR2_X1  g0092(.A(KEYINPUT8), .B(G58), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n206), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(G150), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI22_X1  g0097(.A1(new_n293), .A2(new_n294), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G50), .A2(G58), .ZN(new_n299));
  INV_X1    g0099(.A(G68), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n206), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n280), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT67), .ZN(new_n303));
  INV_X1    g0103(.A(G50), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n302), .A2(new_n303), .B1(new_n304), .B2(new_n287), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n292), .B(new_n305), .C1(new_n303), .C2(new_n302), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n259), .A2(new_n272), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT66), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n273), .ZN(new_n310));
  INV_X1    g0110(.A(G179), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n278), .A2(new_n306), .A3(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT9), .ZN(new_n315));
  OR2_X1    g0115(.A1(new_n306), .A2(new_n315), .ZN(new_n316));
  XOR2_X1   g0116(.A(new_n316), .B(KEYINPUT69), .Z(new_n317));
  INV_X1    g0117(.A(KEYINPUT10), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n306), .A2(new_n315), .ZN(new_n319));
  INV_X1    g0119(.A(G190), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n276), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G200), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n310), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n317), .A2(new_n318), .A3(new_n319), .A4(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n319), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n316), .B(KEYINPUT69), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT10), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n314), .B1(new_n325), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n300), .A2(G20), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n330), .B1(new_n294), .B2(new_n254), .C1(new_n297), .C2(new_n304), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n331), .A2(new_n280), .ZN(new_n332));
  OR2_X1    g0132(.A1(new_n332), .A2(KEYINPUT11), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n205), .A2(G20), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n288), .A2(G68), .A3(new_n334), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n335), .B(KEYINPUT71), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n287), .A2(new_n300), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT12), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n332), .A2(KEYINPUT11), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n333), .A2(new_n336), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  AND2_X1   g0141(.A1(KEYINPUT3), .A2(G33), .ZN(new_n342));
  NOR2_X1   g0142(.A1(KEYINPUT3), .A2(G33), .ZN(new_n343));
  OAI211_X1 g0143(.A(G226), .B(new_n252), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT70), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n342), .A2(new_n343), .ZN(new_n346));
  INV_X1    g0146(.A(G232), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n348), .A2(G1698), .B1(G33), .B2(G97), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n258), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT13), .ZN(new_n352));
  INV_X1    g0152(.A(new_n271), .ZN(new_n353));
  INV_X1    g0153(.A(G238), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n266), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n351), .A2(new_n352), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n261), .A2(new_n262), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n358), .B1(new_n345), .B2(new_n349), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT13), .B1(new_n359), .B2(new_n355), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n341), .B1(new_n361), .B2(new_n320), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n322), .B1(new_n357), .B2(new_n360), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n352), .B1(new_n351), .B2(new_n356), .ZN(new_n365));
  NOR3_X1   g0165(.A1(new_n359), .A2(KEYINPUT13), .A3(new_n355), .ZN(new_n366));
  OAI21_X1  g0166(.A(G169), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT14), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n357), .A2(G179), .A3(new_n360), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT14), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n370), .B(G169), .C1(new_n365), .C2(new_n366), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n368), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n364), .B1(new_n372), .B2(new_n340), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n271), .A2(G244), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n251), .A2(G232), .A3(new_n252), .ZN(new_n375));
  INV_X1    g0175(.A(G107), .ZN(new_n376));
  OAI221_X1 g0176(.A(new_n375), .B1(new_n376), .B2(new_n251), .C1(new_n255), .C2(new_n354), .ZN(new_n377));
  AOI211_X1 g0177(.A(new_n267), .B(new_n374), .C1(new_n377), .C2(new_n258), .ZN(new_n378));
  AND2_X1   g0178(.A1(new_n378), .A2(new_n311), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n288), .A2(G77), .A3(new_n334), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G20), .A2(G77), .ZN(new_n381));
  XNOR2_X1  g0181(.A(KEYINPUT15), .B(G87), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n381), .B1(new_n382), .B2(new_n294), .ZN(new_n383));
  INV_X1    g0183(.A(new_n293), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n383), .B1(new_n296), .B2(new_n384), .ZN(new_n385));
  OAI221_X1 g0185(.A(new_n380), .B1(G77), .B2(new_n284), .C1(new_n385), .C2(new_n281), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n386), .B1(new_n378), .B2(G169), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n379), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n386), .B1(new_n378), .B2(G190), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n322), .B2(new_n378), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g0192(.A(KEYINPUT73), .B(KEYINPUT16), .Z(new_n393));
  NAND2_X1  g0193(.A1(new_n296), .A2(G159), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT72), .ZN(new_n395));
  XNOR2_X1  g0195(.A(G58), .B(G68), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n395), .B1(new_n396), .B2(G20), .ZN(new_n397));
  AND2_X1   g0197(.A1(G58), .A2(G68), .ZN(new_n398));
  NOR2_X1   g0198(.A1(G58), .A2(G68), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n395), .B(G20), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n394), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n249), .A2(new_n206), .A3(new_n250), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT7), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n249), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n250), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n300), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n393), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT7), .B1(new_n346), .B2(new_n206), .ZN(new_n409));
  INV_X1    g0209(.A(new_n406), .ZN(new_n410));
  OAI21_X1  g0210(.A(G68), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(G20), .B1(new_n398), .B2(new_n399), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT72), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n400), .B1(G159), .B2(new_n296), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n411), .A2(new_n414), .A3(KEYINPUT16), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n408), .A2(new_n280), .A3(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n384), .A2(new_n284), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n291), .B2(new_n384), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n256), .A2(new_n252), .ZN(new_n420));
  INV_X1    g0220(.A(G226), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G1698), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n420), .B(new_n422), .C1(new_n342), .C2(new_n343), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G33), .A2(G87), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n358), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n271), .A2(G232), .B1(new_n263), .B2(new_n265), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(new_n311), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n358), .A2(G232), .A3(new_n264), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n266), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n277), .B1(new_n430), .B2(new_n425), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n419), .A2(new_n433), .ZN(new_n434));
  XOR2_X1   g0234(.A(KEYINPUT74), .B(KEYINPUT18), .Z(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OR2_X1    g0236(.A1(KEYINPUT74), .A2(KEYINPUT18), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n436), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n430), .A2(new_n425), .A3(new_n320), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n322), .B1(new_n426), .B2(new_n427), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n441), .A2(new_n416), .A3(new_n418), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT17), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n442), .B(new_n443), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n392), .A2(new_n438), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n329), .A2(new_n373), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G116), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n205), .A2(new_n447), .A3(G13), .A4(G20), .ZN(new_n448));
  XOR2_X1   g0248(.A(new_n448), .B(KEYINPUT78), .Z(new_n449));
  AOI22_X1  g0249(.A1(new_n279), .A2(new_n214), .B1(G20), .B2(new_n447), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G283), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n451), .B(new_n206), .C1(G33), .C2(new_n222), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT79), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n454), .A2(KEYINPUT20), .ZN(new_n455));
  INV_X1    g0255(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(KEYINPUT20), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n453), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n205), .A2(G33), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n288), .A2(G116), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n450), .A2(new_n455), .A3(new_n452), .ZN(new_n461));
  AND4_X1   g0261(.A1(new_n449), .A2(new_n458), .A3(new_n460), .A4(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT80), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n269), .A2(G1), .ZN(new_n464));
  NAND2_X1  g0264(.A1(KEYINPUT5), .A2(G41), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(KEYINPUT5), .A2(G41), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n468), .A2(G270), .A3(new_n358), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n205), .A2(G45), .ZN(new_n470));
  OR2_X1    g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n470), .B1(new_n471), .B2(new_n465), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n263), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(G264), .B(G1698), .C1(new_n342), .C2(new_n343), .ZN(new_n475));
  OAI211_X1 g0275(.A(G257), .B(new_n252), .C1(new_n342), .C2(new_n343), .ZN(new_n476));
  INV_X1    g0276(.A(G303), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n475), .B(new_n476), .C1(new_n477), .C2(new_n251), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n474), .B1(new_n258), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n462), .B(new_n463), .C1(new_n479), .C2(new_n322), .ZN(new_n480));
  AND2_X1   g0280(.A1(new_n469), .A2(new_n473), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n478), .A2(new_n258), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n322), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n449), .A2(new_n458), .A3(new_n460), .A4(new_n461), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT80), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n479), .A2(G190), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n480), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT21), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n481), .A2(new_n482), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n489), .A2(new_n484), .A3(G169), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n489), .A2(new_n311), .ZN(new_n491));
  AOI22_X1  g0291(.A1(new_n488), .A2(new_n490), .B1(new_n491), .B2(new_n484), .ZN(new_n492));
  OR2_X1    g0292(.A1(new_n490), .A2(new_n488), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n487), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT6), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n222), .A2(new_n376), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(new_n202), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n376), .A2(KEYINPUT6), .A3(G97), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n499), .A2(G20), .B1(G77), .B2(new_n296), .ZN(new_n500));
  OAI21_X1  g0300(.A(G107), .B1(new_n409), .B2(new_n410), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n280), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n287), .A2(new_n222), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n288), .A2(new_n459), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n504), .B1(new_n505), .B2(new_n222), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n468), .A2(G257), .A3(new_n358), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n473), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n221), .B1(new_n249), .B2(new_n250), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT4), .ZN(new_n512));
  OAI21_X1  g0312(.A(G1698), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(G244), .B1(new_n342), .B2(new_n343), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n514), .A2(new_n512), .B1(G33), .B2(G283), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n251), .A2(KEYINPUT4), .A3(G244), .A4(new_n252), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n510), .B1(new_n517), .B2(new_n258), .ZN(new_n518));
  AND2_X1   g0318(.A1(new_n518), .A2(G179), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(new_n277), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n508), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n506), .B1(new_n502), .B2(new_n280), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n518), .A2(G190), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n522), .B(new_n523), .C1(new_n322), .C2(new_n518), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n494), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT23), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(new_n206), .B2(G107), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n376), .A2(KEYINPUT23), .A3(G20), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G116), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n528), .A2(new_n529), .B1(new_n531), .B2(new_n206), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n206), .B(G87), .C1(new_n342), .C2(new_n343), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT81), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT81), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n251), .A2(new_n535), .A3(new_n206), .A4(G87), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT22), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n537), .B1(new_n534), .B2(new_n536), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n532), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT82), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT24), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT24), .B1(new_n540), .B2(new_n541), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n534), .A2(new_n536), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(KEYINPUT22), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT82), .B1(new_n548), .B2(new_n532), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n280), .B(new_n543), .C1(new_n544), .C2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n505), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT25), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n284), .B2(G107), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n287), .A2(KEYINPUT25), .A3(new_n376), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n551), .A2(G107), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(G257), .B(G1698), .C1(new_n342), .C2(new_n343), .ZN(new_n557));
  OAI211_X1 g0357(.A(G250), .B(new_n252), .C1(new_n342), .C2(new_n343), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G33), .A2(G294), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n258), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n468), .A2(G264), .A3(new_n358), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT83), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n563), .B1(new_n561), .B2(new_n562), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n473), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n561), .A2(new_n562), .ZN(new_n569));
  INV_X1    g0369(.A(new_n473), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI22_X1  g0371(.A1(new_n568), .A2(new_n311), .B1(new_n277), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n556), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n571), .A2(new_n320), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n565), .A2(new_n566), .A3(new_n570), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n575), .B2(G200), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n550), .A2(new_n576), .A3(new_n555), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n206), .B(G68), .C1(new_n342), .C2(new_n343), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n294), .A2(new_n222), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n578), .B1(KEYINPUT19), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n206), .A2(new_n581), .B1(new_n202), .B2(new_n220), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n280), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n382), .A2(new_n287), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n583), .B(new_n584), .C1(new_n220), .C2(new_n505), .ZN(new_n585));
  OAI211_X1 g0385(.A(G244), .B(G1698), .C1(new_n342), .C2(new_n343), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT75), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT75), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n251), .A2(new_n588), .A3(G244), .A4(G1698), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n251), .A2(G238), .A3(new_n252), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n587), .A2(new_n589), .A3(new_n530), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n258), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n464), .A2(new_n260), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n470), .A2(new_n221), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n358), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT77), .B1(new_n596), .B2(new_n320), .ZN(new_n597));
  INV_X1    g0397(.A(new_n595), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n591), .B2(new_n258), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT77), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n599), .A2(new_n600), .A3(G190), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n585), .B1(new_n597), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n596), .A2(G200), .ZN(new_n603));
  INV_X1    g0403(.A(new_n382), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n288), .A2(new_n459), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n583), .A2(new_n605), .A3(new_n584), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT76), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n599), .A2(new_n311), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT76), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n583), .A2(new_n605), .A3(new_n609), .A4(new_n584), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n596), .A2(new_n277), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n602), .A2(new_n603), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n526), .A2(new_n573), .A3(new_n577), .A4(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n446), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g0415(.A(new_n615), .B(KEYINPUT84), .ZN(G372));
  NAND2_X1  g0416(.A1(new_n325), .A2(new_n328), .ZN(new_n617));
  OR2_X1    g0417(.A1(new_n362), .A2(new_n363), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n388), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n371), .A2(new_n369), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n370), .B1(new_n361), .B2(G169), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n340), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n444), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT18), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT90), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(new_n419), .B2(new_n433), .ZN(new_n626));
  AOI211_X1 g0426(.A(KEYINPUT90), .B(new_n432), .C1(new_n416), .C2(new_n418), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n624), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n288), .A2(new_n289), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n287), .A2(new_n280), .A3(KEYINPUT68), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n334), .B(new_n384), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n417), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n411), .A2(new_n414), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n281), .B1(new_n634), .B2(new_n393), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n633), .B1(new_n635), .B2(new_n415), .ZN(new_n636));
  OAI21_X1  g0436(.A(KEYINPUT90), .B1(new_n636), .B2(new_n432), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n419), .A2(new_n625), .A3(new_n433), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n637), .A2(KEYINPUT18), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n628), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n617), .B1(new_n623), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n313), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT85), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n591), .A2(new_n645), .A3(new_n258), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n645), .B1(new_n591), .B2(new_n258), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n595), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n277), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n611), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT87), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT26), .ZN(new_n653));
  INV_X1    g0453(.A(new_n585), .ZN(new_n654));
  INV_X1    g0454(.A(new_n601), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n600), .B1(new_n599), .B2(G190), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n592), .A2(KEYINPUT85), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n598), .B1(new_n658), .B2(new_n646), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(new_n322), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(G169), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n607), .A2(new_n608), .A3(new_n610), .ZN(new_n662));
  OAI22_X1  g0462(.A1(new_n657), .A2(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n518), .A2(G179), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n277), .B2(new_n518), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT88), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n522), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n664), .B(KEYINPUT88), .C1(new_n277), .C2(new_n518), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI211_X1 g0469(.A(KEYINPUT89), .B(new_n653), .C1(new_n663), .C2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n521), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n613), .A2(KEYINPUT26), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n649), .A2(G200), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n602), .A2(new_n674), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n675), .A2(new_n651), .A3(new_n668), .A4(new_n667), .ZN(new_n676));
  AOI21_X1  g0476(.A(KEYINPUT89), .B1(new_n676), .B2(new_n653), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n652), .B1(new_n673), .B2(new_n677), .ZN(new_n678));
  AOI22_X1  g0478(.A1(new_n602), .A2(new_n674), .B1(new_n650), .B2(new_n611), .ZN(new_n679));
  INV_X1    g0479(.A(new_n525), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(new_n680), .A3(new_n577), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT86), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n679), .A2(new_n680), .A3(new_n577), .A4(KEYINPUT86), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n492), .A2(new_n493), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n685), .B1(new_n556), .B2(new_n572), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  AND3_X1   g0487(.A1(new_n683), .A2(new_n684), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n678), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n644), .B1(new_n446), .B2(new_n689), .ZN(new_n690));
  XNOR2_X1  g0490(.A(new_n690), .B(KEYINPUT91), .ZN(G369));
  AND2_X1   g0491(.A1(new_n556), .A2(new_n572), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n283), .A2(new_n206), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(KEYINPUT27), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(new_n695), .A3(G213), .ZN(new_n696));
  INV_X1    g0496(.A(G343), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n556), .A2(new_n698), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n573), .A2(new_n700), .A3(new_n577), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(G330), .ZN(new_n704));
  INV_X1    g0504(.A(new_n698), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n462), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n494), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n685), .A2(new_n706), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n704), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n703), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n692), .A2(new_n705), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n573), .A2(new_n577), .A3(new_n685), .A4(new_n705), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(G399));
  INV_X1    g0513(.A(new_n209), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G41), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(G1), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n212), .B2(new_n716), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n721), .B1(new_n689), .B2(new_n698), .ZN(new_n722));
  OAI21_X1  g0522(.A(KEYINPUT26), .B1(new_n663), .B2(new_n669), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n613), .A2(new_n653), .A3(new_n671), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(new_n652), .A3(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n681), .A2(new_n686), .ZN(new_n726));
  OAI211_X1 g0526(.A(KEYINPUT29), .B(new_n705), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT95), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n722), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n518), .A2(new_n599), .A3(new_n479), .A4(G179), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n569), .A2(KEYINPUT83), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n564), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT30), .ZN(new_n736));
  NOR3_X1   g0536(.A1(new_n518), .A2(new_n479), .A3(G179), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n568), .A2(new_n649), .A3(new_n737), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT94), .ZN(new_n740));
  XOR2_X1   g0540(.A(KEYINPUT93), .B(KEYINPUT30), .Z(new_n741));
  INV_X1    g0541(.A(KEYINPUT92), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n741), .B1(new_n735), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(KEYINPUT92), .B1(new_n732), .B2(new_n734), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n740), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n599), .A2(new_n479), .A3(G179), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n746), .A2(new_n567), .A3(new_n742), .A4(new_n518), .ZN(new_n747));
  INV_X1    g0547(.A(new_n741), .ZN(new_n748));
  AND4_X1   g0548(.A1(new_n740), .A2(new_n747), .A3(new_n744), .A4(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n739), .B1(new_n745), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT31), .B1(new_n750), .B2(new_n698), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n736), .A2(new_n738), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n752), .B1(new_n744), .B2(new_n743), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n698), .A2(KEYINPUT31), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n614), .A2(new_n698), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G330), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n731), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n720), .B1(new_n758), .B2(G1), .ZN(G364));
  NOR3_X1   g0559(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n707), .A2(new_n708), .A3(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n282), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n205), .B1(new_n762), .B2(G45), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n715), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n242), .A2(new_n269), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n714), .A2(new_n251), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(G45), .B2(new_n212), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT96), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n766), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(new_n769), .B2(new_n768), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n714), .A2(new_n346), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n772), .A2(G355), .B1(new_n447), .B2(new_n714), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n774), .A2(KEYINPUT97), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n214), .B1(G20), .B2(new_n277), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n760), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(new_n774), .B2(KEYINPUT97), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n765), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n322), .A2(G190), .ZN(new_n780));
  OAI21_X1  g0580(.A(G20), .B1(new_n780), .B2(G179), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT100), .ZN(new_n782));
  OR2_X1    g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n786), .A2(KEYINPUT101), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(KEYINPUT101), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G97), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n206), .A2(G179), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n792), .A2(G190), .A3(G200), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n792), .A2(new_n320), .A3(G200), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n220), .A2(new_n793), .B1(new_n794), .B2(new_n376), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n206), .A2(new_n311), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n780), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n346), .B1(new_n798), .B2(G58), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G190), .A2(G200), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n796), .A2(new_n800), .ZN(new_n801));
  NOR3_X1   g0601(.A1(new_n797), .A2(new_n320), .A3(new_n322), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n799), .B1(new_n254), .B2(new_n801), .C1(new_n803), .C2(new_n304), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n797), .A2(new_n322), .A3(G190), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n805), .A2(KEYINPUT99), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(KEYINPUT99), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n795), .B(new_n804), .C1(G68), .C2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n792), .A2(new_n800), .ZN(new_n810));
  OR2_X1    g0610(.A1(new_n810), .A2(KEYINPUT98), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(KEYINPUT98), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(G159), .ZN(new_n814));
  OAI21_X1  g0614(.A(KEYINPUT32), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OR3_X1    g0615(.A1(new_n813), .A2(KEYINPUT32), .A3(new_n814), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n791), .A2(new_n809), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G311), .ZN(new_n818));
  INV_X1    g0618(.A(new_n798), .ZN(new_n819));
  INV_X1    g0619(.A(G322), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n346), .B1(new_n818), .B2(new_n801), .C1(new_n819), .C2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n808), .ZN(new_n822));
  XOR2_X1   g0622(.A(KEYINPUT33), .B(G317), .Z(new_n823));
  XNOR2_X1  g0623(.A(new_n802), .B(KEYINPUT102), .ZN(new_n824));
  INV_X1    g0624(.A(G326), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n822), .A2(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n793), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n821), .B(new_n826), .C1(G303), .C2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(G294), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n829), .B2(new_n786), .ZN(new_n830));
  INV_X1    g0630(.A(new_n813), .ZN(new_n831));
  INV_X1    g0631(.A(new_n794), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n831), .A2(G329), .B1(G283), .B2(new_n832), .ZN(new_n833));
  XOR2_X1   g0633(.A(new_n833), .B(KEYINPUT103), .Z(new_n834));
  OAI21_X1  g0634(.A(new_n817), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n779), .B1(new_n835), .B2(new_n776), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n709), .A2(new_n765), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n707), .A2(new_n704), .A3(new_n708), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n761), .A2(new_n836), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(G396));
  NAND2_X1  g0640(.A1(new_n386), .A2(new_n698), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n391), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n389), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n388), .A2(new_n705), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n689), .B2(new_n698), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n392), .A2(new_n698), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n678), .B2(new_n688), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n765), .B1(new_n849), .B2(new_n757), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n757), .B2(new_n849), .ZN(new_n851));
  NOR2_X1   g0651(.A1(G13), .A2(G33), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n845), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n776), .A2(new_n852), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n765), .B1(G77), .B2(new_n855), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT104), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n808), .A2(KEYINPUT105), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n808), .A2(KEYINPUT105), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(G283), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n813), .A2(new_n818), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n251), .B1(new_n798), .B2(G294), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n864), .B1(new_n447), .B2(new_n801), .C1(new_n803), .C2(new_n477), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n220), .A2(new_n794), .B1(new_n793), .B2(new_n376), .ZN(new_n866));
  NOR4_X1   g0666(.A1(new_n862), .A2(new_n863), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(G132), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n251), .B1(new_n813), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n832), .A2(G68), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n304), .B2(new_n793), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT106), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n869), .B(new_n872), .C1(G58), .C2(new_n785), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n802), .A2(G137), .B1(new_n798), .B2(G143), .ZN(new_n874));
  OAI221_X1 g0674(.A(new_n874), .B1(new_n814), .B2(new_n801), .C1(new_n822), .C2(new_n295), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n875), .B(KEYINPUT34), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n867), .A2(new_n791), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n776), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n853), .B(new_n857), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n851), .A2(new_n879), .ZN(G384));
  NOR2_X1   g0680(.A1(new_n762), .A2(new_n205), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n340), .B(new_n698), .C1(new_n372), .C2(new_n364), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n340), .A2(new_n698), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n622), .A2(new_n618), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n845), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n743), .A2(new_n740), .A3(new_n744), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n747), .A2(new_n744), .A3(new_n748), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT94), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n752), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  OAI22_X1  g0689(.A1(new_n889), .A2(new_n754), .B1(new_n614), .B2(new_n698), .ZN(new_n890));
  OAI211_X1 g0690(.A(KEYINPUT40), .B(new_n885), .C1(new_n890), .C2(new_n751), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT108), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n442), .B(KEYINPUT17), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n626), .A2(new_n627), .A3(new_n624), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT18), .B1(new_n637), .B2(new_n638), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT107), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(new_n636), .B2(new_n696), .ZN(new_n899));
  INV_X1    g0699(.A(new_n696), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n419), .A2(KEYINPUT107), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n442), .B1(new_n626), .B2(new_n627), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT37), .B1(new_n903), .B2(new_n902), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n434), .A2(new_n442), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n905), .A2(KEYINPUT37), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT107), .B1(new_n419), .B2(new_n900), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n898), .B(new_n696), .C1(new_n416), .C2(new_n418), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n897), .A2(new_n902), .B1(new_n904), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n893), .B1(new_n911), .B2(KEYINPUT38), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n419), .A2(new_n900), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n434), .A2(new_n913), .A3(new_n442), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT37), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n419), .B(new_n900), .C1(new_n438), .C2(new_n444), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT38), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT38), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n909), .B(new_n442), .C1(new_n626), .C2(new_n627), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n920), .A2(KEYINPUT37), .B1(new_n909), .B2(new_n906), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n909), .B1(new_n640), .B2(new_n894), .ZN(new_n922));
  OAI211_X1 g0722(.A(KEYINPUT108), .B(new_n919), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n912), .A2(new_n918), .A3(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT109), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n892), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n925), .B1(new_n892), .B2(new_n924), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT40), .ZN(new_n930));
  OR2_X1    g0730(.A1(new_n890), .A2(new_n751), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n636), .A2(new_n432), .A3(new_n437), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n434), .B2(new_n435), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n913), .B1(new_n933), .B2(new_n894), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n906), .A2(new_n909), .B1(new_n914), .B2(KEYINPUT37), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n919), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n918), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n931), .A2(new_n937), .A3(new_n885), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n927), .A2(new_n929), .B1(new_n930), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n890), .A2(new_n751), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n446), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n704), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n939), .B2(new_n941), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n372), .A2(new_n340), .A3(new_n705), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT39), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n937), .A2(new_n945), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n944), .B(new_n946), .C1(new_n924), .C2(new_n945), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n683), .A2(new_n684), .A3(new_n687), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n948), .B(new_n652), .C1(new_n677), .C2(new_n673), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n949), .A2(new_n847), .B1(new_n388), .B2(new_n705), .ZN(new_n950));
  INV_X1    g0750(.A(new_n937), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n884), .A2(new_n882), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n950), .A2(new_n951), .A3(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n640), .A2(new_n900), .ZN(new_n955));
  NOR3_X1   g0755(.A1(new_n947), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  AND3_X1   g0756(.A1(new_n722), .A2(new_n729), .A3(new_n730), .ZN(new_n957));
  INV_X1    g0757(.A(new_n446), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n643), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n956), .B(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n881), .B1(new_n943), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n960), .B2(new_n943), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n499), .A2(KEYINPUT35), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n963), .A2(G116), .A3(new_n215), .A4(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT36), .ZN(new_n966));
  NOR3_X1   g0766(.A1(new_n212), .A2(new_n398), .A3(new_n254), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n300), .A2(G50), .ZN(new_n968));
  OAI211_X1 g0768(.A(G1), .B(new_n282), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n962), .A2(new_n966), .A3(new_n969), .ZN(G367));
  OAI21_X1  g0770(.A(new_n680), .B1(new_n522), .B2(new_n705), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n667), .A2(new_n668), .A3(new_n698), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(KEYINPUT42), .B1(new_n974), .B2(new_n712), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n711), .A2(new_n712), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n711), .A2(KEYINPUT42), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n976), .A2(new_n977), .A3(new_n973), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n975), .B(new_n978), .C1(new_n521), .C2(new_n698), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n585), .A2(new_n698), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n679), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n652), .A2(new_n980), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT110), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(new_n983), .B2(new_n982), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT43), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n979), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n985), .A2(new_n986), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n987), .B(new_n988), .Z(new_n989));
  NOR2_X1   g0789(.A1(new_n710), .A2(new_n974), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n715), .B(KEYINPUT41), .Z(new_n992));
  NAND2_X1  g0792(.A1(new_n685), .A2(new_n705), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n702), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT113), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n709), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n994), .A2(new_n712), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n709), .A2(new_n995), .ZN(new_n998));
  INV_X1    g0798(.A(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n997), .B(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n731), .A2(new_n1000), .A3(new_n757), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT111), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT44), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n973), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n976), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1006), .A2(KEYINPUT111), .A3(KEYINPUT44), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n973), .A2(new_n711), .A3(new_n712), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT45), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1005), .B(new_n976), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1007), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n710), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(KEYINPUT112), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT112), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1012), .A2(new_n1016), .A3(new_n1013), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1007), .A2(new_n1010), .A3(new_n710), .A4(new_n1011), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1002), .A2(new_n1015), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n992), .B1(new_n1019), .B2(new_n758), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n763), .B1(new_n1020), .B2(KEYINPUT114), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n758), .B1(new_n1022), .B2(new_n1001), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n992), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT114), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n991), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n767), .A2(new_n238), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1029), .B(new_n777), .C1(new_n209), .C2(new_n382), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n819), .A2(new_n295), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n789), .A2(new_n300), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n824), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n1031), .B(new_n1032), .C1(G143), .C2(new_n1033), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1034), .A2(KEYINPUT117), .ZN(new_n1035));
  INV_X1    g0835(.A(G137), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n813), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n801), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n346), .B1(new_n1038), .B2(G50), .ZN(new_n1039));
  INV_X1    g0839(.A(G58), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1039), .B1(new_n1040), .B2(new_n793), .C1(new_n254), .C2(new_n794), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n860), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1037), .B(new_n1041), .C1(new_n1042), .C2(G159), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1034), .A2(KEYINPUT117), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1035), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT118), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1042), .A2(G294), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n346), .B1(new_n222), .B2(new_n794), .C1(new_n819), .C2(new_n477), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(G317), .B2(new_n831), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT46), .ZN(new_n1050));
  NOR3_X1   g0850(.A1(new_n793), .A2(new_n1050), .A3(new_n447), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(new_n1033), .B2(G311), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1050), .B1(new_n793), .B2(new_n447), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT116), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1047), .A2(new_n1049), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n785), .A2(G107), .B1(G283), .B2(new_n1038), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT115), .Z(new_n1057));
  OAI21_X1  g0857(.A(new_n1046), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT47), .Z(new_n1059));
  OAI211_X1 g0859(.A(new_n765), .B(new_n1030), .C1(new_n1059), .C2(new_n878), .ZN(new_n1060));
  AND2_X1   g0860(.A1(new_n985), .A2(new_n760), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1028), .A2(new_n1063), .ZN(G387));
  INV_X1    g0864(.A(new_n772), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n1065), .A2(new_n717), .B1(G107), .B2(new_n209), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT119), .Z(new_n1067));
  NAND2_X1  g0867(.A1(new_n235), .A2(G45), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n293), .A2(G50), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT50), .ZN(new_n1070));
  AOI21_X1  g0870(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1070), .A2(new_n717), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1068), .A2(new_n767), .A3(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1067), .A2(KEYINPUT120), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n777), .ZN(new_n1075));
  AOI21_X1  g0875(.A(KEYINPUT120), .B1(new_n1067), .B2(new_n1073), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n765), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n790), .A2(new_n604), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n793), .A2(new_n254), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G50), .A2(new_n798), .B1(new_n1038), .B2(G68), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1080), .B(new_n251), .C1(new_n814), .C2(new_n803), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1079), .B(new_n1081), .C1(G97), .C2(new_n832), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n808), .A2(new_n384), .B1(G150), .B2(new_n831), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1078), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n786), .A2(new_n861), .B1(new_n829), .B2(new_n793), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G317), .A2(new_n798), .B1(new_n1038), .B2(G303), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1086), .B1(new_n820), .B2(new_n824), .C1(new_n860), .C2(new_n818), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT48), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1085), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n1088), .B2(new_n1087), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(KEYINPUT121), .B(KEYINPUT49), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1090), .B(new_n1091), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n346), .B1(new_n447), .B2(new_n794), .C1(new_n813), .C2(new_n825), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1084), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1077), .B1(new_n1094), .B2(new_n776), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n702), .A2(new_n760), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n764), .A2(new_n1000), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n758), .A2(new_n1000), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1001), .A2(new_n715), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(G393));
  NAND2_X1  g0900(.A1(new_n974), .A2(new_n760), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n802), .A2(G317), .B1(new_n798), .B2(G311), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT52), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(G322), .B2(new_n831), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n251), .B1(new_n1038), .B2(G294), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1105), .B1(new_n376), .B2(new_n794), .C1(new_n861), .C2(new_n793), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(G116), .B2(new_n785), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1104), .B(new_n1107), .C1(new_n477), .C2(new_n860), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n802), .A2(G150), .B1(new_n798), .B2(G159), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(KEYINPUT122), .B(KEYINPUT51), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1109), .B(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(G143), .B2(new_n831), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n794), .A2(new_n220), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n251), .B1(new_n801), .B2(new_n293), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1113), .B(new_n1114), .C1(G68), .C2(new_n827), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1112), .B(new_n1115), .C1(new_n304), .C2(new_n860), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n789), .A2(new_n254), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1108), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n776), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n767), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n777), .B1(new_n222), .B2(new_n209), .C1(new_n1120), .C2(new_n245), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1101), .A2(new_n765), .A3(new_n1119), .A4(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1122), .B1(new_n1123), .B2(new_n763), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n715), .B1(new_n1022), .B2(new_n1001), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1001), .A2(new_n1123), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT123), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1001), .A2(new_n1123), .A3(KEYINPUT123), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1127), .A2(KEYINPUT124), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(KEYINPUT124), .B1(new_n1127), .B2(new_n1132), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1125), .B1(new_n1134), .B2(new_n1135), .ZN(G390));
  NOR3_X1   g0936(.A1(new_n934), .A2(new_n935), .A3(new_n919), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1137), .B1(new_n1138), .B2(new_n893), .ZN(new_n1139));
  AOI21_X1  g0939(.A(KEYINPUT39), .B1(new_n1139), .B2(new_n923), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n953), .B1(new_n848), .B2(new_n844), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n944), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n1140), .A2(new_n946), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n705), .B(new_n843), .C1(new_n725), .C2(new_n726), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n844), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(KEYINPUT125), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT125), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1144), .A2(new_n1147), .A3(new_n844), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1146), .A2(new_n952), .A3(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1142), .B1(new_n1139), .B2(new_n923), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n845), .ZN(new_n1152));
  OAI211_X1 g0952(.A(G330), .B(new_n1152), .C1(new_n751), .C2(new_n755), .ZN(new_n1153));
  OR2_X1    g0953(.A1(new_n1153), .A2(new_n953), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1143), .A2(new_n1151), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n946), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n924), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1156), .B1(new_n1157), .B2(KEYINPUT39), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n944), .B1(new_n950), .B2(new_n953), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1158), .A2(new_n1159), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n940), .A2(new_n704), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n885), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1155), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n958), .A2(new_n1161), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n644), .B(new_n1164), .C1(new_n731), .C2(new_n446), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n931), .A2(G330), .A3(new_n1152), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1167), .A2(new_n953), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n1154), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n1161), .A2(new_n885), .B1(new_n953), .B2(new_n1153), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n1169), .A2(new_n1171), .B1(new_n950), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1166), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n716), .B1(new_n1163), .B2(new_n1174), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n1143), .A2(new_n1151), .A3(new_n1154), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1162), .B1(new_n1143), .B2(new_n1151), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  AND2_X1   g0978(.A1(new_n1168), .A2(new_n1154), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n1170), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1172), .A2(new_n950), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1165), .B1(new_n1180), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1178), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1175), .A2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1155), .B(new_n764), .C1(new_n1160), .C2(new_n1162), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1158), .A2(new_n852), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n765), .B1(new_n384), .B2(new_n855), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n827), .A2(G150), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(new_n1189), .B(KEYINPUT53), .ZN(new_n1190));
  INV_X1    g0990(.A(G128), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n251), .B1(new_n803), .B2(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(KEYINPUT54), .B(G143), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n819), .A2(new_n868), .B1(new_n801), .B2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n304), .B2(new_n794), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1190), .B(new_n1196), .C1(G125), .C2(new_n831), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1197), .B1(new_n1036), .B2(new_n860), .C1(new_n814), .C2(new_n789), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n870), .B1(new_n813), .B2(new_n829), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT126), .Z(new_n1200));
  OAI21_X1  g1000(.A(new_n346), .B1(new_n801), .B2(new_n222), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n803), .A2(new_n861), .B1(new_n819), .B2(new_n447), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(G87), .C2(new_n827), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n1200), .B(new_n1203), .C1(new_n860), .C2(new_n376), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1198), .B1(new_n1117), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1188), .B1(new_n1205), .B2(new_n776), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1187), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1186), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1185), .A2(new_n1209), .ZN(G378));
  AOI21_X1  g1010(.A(new_n704), .B1(new_n938), .B2(new_n930), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n926), .B2(new_n928), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n306), .A2(new_n900), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n329), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n329), .A2(new_n1215), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1214), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OR2_X1    g1019(.A1(new_n329), .A2(new_n1215), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1220), .A2(new_n1216), .A3(new_n1213), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1212), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1224), .B(new_n1211), .C1(new_n926), .C2(new_n928), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n1223), .A2(new_n956), .A3(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n956), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1227));
  OAI21_X1  g1027(.A(KEYINPUT57), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1165), .B1(new_n1178), .B2(new_n1183), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n715), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n956), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1223), .A2(new_n1225), .A3(new_n956), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1181), .B1(new_n1179), .B2(new_n1170), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1166), .B1(new_n1163), .B2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT57), .B1(new_n1235), .B2(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1230), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1222), .A2(new_n852), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n802), .A2(G125), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n1036), .B2(new_n801), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G128), .B2(new_n798), .ZN(new_n1243));
  OAI221_X1 g1043(.A(new_n1243), .B1(new_n793), .B2(new_n1193), .C1(new_n822), .C2(new_n868), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(G150), .B2(new_n790), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1246), .A2(KEYINPUT59), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(KEYINPUT59), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n831), .A2(G124), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n248), .B(new_n268), .C1(new_n794), .C2(new_n814), .ZN(new_n1250));
  NOR4_X1   g1050(.A1(new_n1247), .A2(new_n1248), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n803), .A2(new_n447), .B1(new_n819), .B2(new_n376), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n268), .B(new_n346), .C1(new_n801), .C2(new_n382), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n794), .A2(new_n1040), .ZN(new_n1254));
  NOR4_X1   g1054(.A1(new_n1252), .A2(new_n1253), .A3(new_n1079), .A4(new_n1254), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1255), .B1(new_n222), .B2(new_n822), .C1(new_n861), .C2(new_n813), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1256), .A2(new_n1032), .ZN(new_n1257));
  OR2_X1    g1057(.A1(new_n1257), .A2(KEYINPUT58), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(KEYINPUT58), .ZN(new_n1259));
  AOI21_X1  g1059(.A(G50), .B1(new_n248), .B2(new_n268), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n251), .B2(G41), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1258), .A2(new_n1259), .A3(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n776), .B1(new_n1251), .B2(new_n1262), .ZN(new_n1263));
  XOR2_X1   g1063(.A(new_n1263), .B(KEYINPUT127), .Z(new_n1264));
  OAI21_X1  g1064(.A(new_n765), .B1(G50), .B2(new_n855), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1235), .A2(new_n764), .B1(new_n1240), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1239), .A2(new_n1267), .ZN(G375));
  NAND2_X1  g1068(.A1(new_n953), .A2(new_n852), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n765), .B1(G68), .B2(new_n855), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n254), .A2(new_n794), .B1(new_n793), .B2(new_n222), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(G283), .A2(new_n798), .B1(new_n1038), .B2(G107), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1272), .B(new_n346), .C1(new_n829), .C2(new_n803), .ZN(new_n1273));
  AOI211_X1 g1073(.A(new_n1271), .B(new_n1273), .C1(G303), .C2(new_n831), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1078), .B(new_n1274), .C1(new_n447), .C2(new_n860), .ZN(new_n1275));
  OAI22_X1  g1075(.A1(new_n1040), .A2(new_n794), .B1(new_n793), .B2(new_n814), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(G137), .A2(new_n798), .B1(new_n1038), .B2(G150), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1277), .B(new_n251), .C1(new_n868), .C2(new_n803), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n1276), .B(new_n1278), .C1(G128), .C2(new_n831), .ZN(new_n1279));
  OAI221_X1 g1079(.A(new_n1279), .B1(new_n304), .B2(new_n789), .C1(new_n860), .C2(new_n1193), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1275), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1270), .B1(new_n1281), .B2(new_n776), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(new_n1173), .A2(new_n764), .B1(new_n1269), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1174), .A2(new_n1024), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1166), .A2(new_n1173), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1283), .B1(new_n1284), .B2(new_n1285), .ZN(G381));
  NOR4_X1   g1086(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1208), .B1(new_n1175), .B2(new_n1184), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT124), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1290), .B1(new_n1291), .B2(new_n1126), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1124), .B1(new_n1292), .B2(new_n1133), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1028), .A2(new_n1293), .A3(new_n1063), .ZN(new_n1294));
  OR3_X1    g1094(.A1(new_n1289), .A2(G375), .A3(new_n1294), .ZN(G407));
  NAND2_X1  g1095(.A1(new_n1288), .A2(new_n697), .ZN(new_n1296));
  OAI211_X1 g1096(.A(G407), .B(G213), .C1(G375), .C2(new_n1296), .ZN(G409));
  INV_X1    g1097(.A(KEYINPUT63), .ZN(new_n1298));
  OAI211_X1 g1098(.A(G378), .B(new_n1267), .C1(new_n1230), .C2(new_n1238), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1235), .A2(new_n1024), .A3(new_n1237), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n764), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1240), .A2(new_n1266), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1288), .B1(new_n1300), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1299), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(G213), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1306), .A2(G343), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1305), .A2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1174), .A2(new_n715), .ZN(new_n1310));
  OAI21_X1  g1110(.A(KEYINPUT60), .B1(new_n1166), .B2(new_n1173), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT60), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1236), .A2(new_n1312), .A3(new_n1165), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1310), .B1(new_n1311), .B2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(G384), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1283), .ZN(new_n1316));
  NOR3_X1   g1116(.A1(new_n1314), .A2(new_n1315), .A3(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1183), .A2(new_n716), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(G384), .B1(new_n1320), .B2(new_n1283), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1317), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1298), .B1(new_n1309), .B2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n991), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n764), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1020), .A2(KEYINPUT114), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1325), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(G390), .B1(new_n1328), .B2(new_n1062), .ZN(new_n1329));
  XNOR2_X1  g1129(.A(G393), .B(G396), .ZN(new_n1330));
  AND3_X1   g1130(.A1(new_n1329), .A2(new_n1294), .A3(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1330), .B1(new_n1329), .B2(new_n1294), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1307), .A2(G2897), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  NOR3_X1   g1135(.A1(new_n1317), .A2(new_n1321), .A3(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1315), .B1(new_n1314), .B2(new_n1316), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1320), .A2(G384), .A3(new_n1283), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1334), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1336), .A2(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(KEYINPUT61), .B1(new_n1309), .B2(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1307), .B1(new_n1299), .B2(new_n1304), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1342), .A2(KEYINPUT63), .A3(new_n1322), .ZN(new_n1343));
  NAND4_X1  g1143(.A1(new_n1324), .A2(new_n1333), .A3(new_n1341), .A4(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT62), .ZN(new_n1345));
  AND3_X1   g1145(.A1(new_n1342), .A2(new_n1345), .A3(new_n1322), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT61), .ZN(new_n1347));
  OAI21_X1  g1147(.A(new_n1335), .B1(new_n1317), .B2(new_n1321), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1337), .A2(new_n1338), .A3(new_n1334), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1348), .A2(new_n1349), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1347), .B1(new_n1342), .B2(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1345), .B1(new_n1342), .B2(new_n1322), .ZN(new_n1352));
  NOR3_X1   g1152(.A1(new_n1346), .A2(new_n1351), .A3(new_n1352), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1344), .B1(new_n1353), .B2(new_n1333), .ZN(G405));
  NAND2_X1  g1154(.A1(G375), .A2(new_n1288), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1355), .A2(new_n1323), .A3(new_n1299), .ZN(new_n1356));
  INV_X1    g1156(.A(new_n1356), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1323), .B1(new_n1355), .B2(new_n1299), .ZN(new_n1358));
  OAI22_X1  g1158(.A1(new_n1357), .A2(new_n1358), .B1(new_n1332), .B2(new_n1331), .ZN(new_n1359));
  INV_X1    g1159(.A(new_n1358), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1360), .A2(new_n1333), .A3(new_n1356), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1359), .A2(new_n1361), .ZN(G402));
endmodule


