//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 0 0 1 0 0 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n789, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT85), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT85), .A2(G107), .ZN(new_n193));
  AOI21_X1  g007(.A(G104), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n191), .A2(G104), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(G101), .B1(new_n194), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT86), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(KEYINPUT3), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(new_n192), .A3(new_n193), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n202), .B1(G104), .B2(new_n191), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(G101), .B1(new_n199), .B2(G107), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  AND3_X1   g020(.A1(new_n197), .A2(new_n198), .A3(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n198), .B1(new_n197), .B2(new_n206), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G143), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT1), .B1(new_n210), .B2(G146), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(G146), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G143), .ZN(new_n214));
  OAI211_X1 g028(.A(G128), .B(new_n211), .C1(new_n212), .C2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(G143), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n210), .A2(G146), .ZN(new_n217));
  INV_X1    g031(.A(G128), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n216), .B(new_n217), .C1(KEYINPUT1), .C2(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n209), .A2(new_n220), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n215), .A2(new_n219), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n222), .A2(new_n206), .A3(new_n197), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT71), .ZN(new_n225));
  INV_X1    g039(.A(G137), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT64), .B1(new_n226), .B2(G134), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT64), .ZN(new_n228));
  INV_X1    g042(.A(G134), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n229), .A3(G137), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT11), .B1(new_n229), .B2(G137), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT11), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(new_n226), .A3(G134), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(KEYINPUT65), .A2(G131), .ZN(new_n236));
  AND3_X1   g050(.A1(new_n231), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n236), .B1(new_n231), .B2(new_n235), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n225), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n235), .A2(new_n227), .A3(new_n230), .ZN(new_n240));
  INV_X1    g054(.A(new_n236), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n231), .A2(new_n235), .A3(new_n236), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(KEYINPUT71), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n239), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n224), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT12), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n248), .B1(new_n242), .B2(new_n243), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n224), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT87), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n253), .B1(new_n207), .B2(new_n208), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n201), .A2(new_n204), .A3(new_n205), .ZN(new_n255));
  INV_X1    g069(.A(G101), .ZN(new_n256));
  AND2_X1   g070(.A1(KEYINPUT85), .A2(G107), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT85), .A2(G107), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n199), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n256), .B1(new_n259), .B2(new_n195), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT86), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n197), .A2(new_n206), .A3(new_n198), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n261), .A2(KEYINPUT87), .A3(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT10), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT72), .B1(new_n215), .B2(new_n219), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n215), .A2(KEYINPUT72), .A3(new_n219), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n264), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n254), .A2(new_n263), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n199), .A2(G107), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n201), .A2(new_n204), .A3(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(KEYINPUT4), .A3(G101), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n257), .A2(new_n258), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n203), .B1(new_n273), .B2(new_n200), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n256), .B1(new_n274), .B2(new_n270), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT4), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n276), .B1(new_n274), .B2(new_n205), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n272), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT0), .A4(G128), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n212), .A2(new_n214), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT0), .B(G128), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT70), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n279), .B(new_n284), .C1(new_n280), .C2(new_n281), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n278), .A2(new_n286), .B1(new_n264), .B2(new_n223), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n269), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n288), .A2(new_n246), .ZN(new_n289));
  INV_X1    g103(.A(G953), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G227), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n291), .B(KEYINPUT84), .ZN(new_n292));
  XNOR2_X1  g106(.A(G110), .B(G140), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n252), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT88), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n288), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n269), .A2(KEYINPUT88), .A3(new_n287), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n246), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT89), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n245), .B1(new_n288), .B2(new_n298), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT89), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(new_n300), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n289), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n297), .B1(new_n306), .B2(new_n294), .ZN(new_n307));
  INV_X1    g121(.A(G469), .ZN(new_n308));
  INV_X1    g122(.A(G902), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n308), .A2(new_n309), .ZN(new_n311));
  INV_X1    g125(.A(new_n289), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n294), .B1(new_n252), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n302), .A2(new_n305), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n313), .B1(new_n314), .B2(new_n296), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n311), .B1(new_n315), .B2(G469), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n189), .B1(new_n310), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT92), .ZN(new_n318));
  INV_X1    g132(.A(G237), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(new_n290), .A3(G214), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n210), .ZN(new_n321));
  NOR2_X1   g135(.A1(G237), .A2(G953), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(G143), .A3(G214), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n318), .B1(new_n324), .B2(G131), .ZN(new_n325));
  INV_X1    g139(.A(G131), .ZN(new_n326));
  AOI211_X1 g140(.A(KEYINPUT92), .B(new_n326), .C1(new_n321), .C2(new_n323), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT17), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G140), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G125), .ZN(new_n330));
  INV_X1    g144(.A(G125), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G140), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n330), .A2(new_n332), .A3(KEYINPUT16), .ZN(new_n333));
  OR3_X1    g147(.A1(new_n331), .A2(KEYINPUT16), .A3(G140), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n334), .A3(G146), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(G146), .B1(new_n333), .B2(new_n334), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n320), .A2(new_n210), .ZN(new_n339));
  AOI21_X1  g153(.A(G143), .B1(new_n322), .B2(G214), .ZN(new_n340));
  OAI21_X1  g154(.A(G131), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT92), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n324), .A2(new_n318), .A3(G131), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n339), .A2(new_n340), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(new_n326), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n342), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n328), .B(new_n338), .C1(new_n346), .C2(KEYINPUT17), .ZN(new_n347));
  XNOR2_X1  g161(.A(G113), .B(G122), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(new_n199), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n330), .A2(new_n332), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(G125), .B(G140), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT81), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n354), .A3(new_n213), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(new_n213), .B2(new_n353), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT18), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n344), .B1(new_n357), .B2(new_n326), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n324), .A2(KEYINPUT18), .A3(G131), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n347), .A2(new_n349), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n349), .B1(new_n347), .B2(new_n360), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n309), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G475), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT20), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT19), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n351), .B1(new_n366), .B2(KEYINPUT93), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n353), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(KEYINPUT93), .B1(new_n350), .B2(new_n351), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n368), .B1(new_n369), .B2(KEYINPUT19), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n336), .B1(new_n370), .B2(new_n213), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n346), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n360), .ZN(new_n373));
  INV_X1    g187(.A(new_n349), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n347), .A2(new_n349), .A3(new_n360), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(G475), .A2(G902), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n365), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n378), .ZN(new_n380));
  AOI211_X1 g194(.A(KEYINPUT20), .B(new_n380), .C1(new_n375), .C2(new_n376), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n364), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT94), .ZN(new_n383));
  INV_X1    g197(.A(G122), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n383), .B1(new_n384), .B2(G116), .ZN(new_n385));
  INV_X1    g199(.A(G116), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(KEYINPUT94), .A3(G122), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT14), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n384), .A2(G116), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT14), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n385), .A2(new_n391), .A3(new_n387), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G107), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n388), .A2(new_n273), .A3(new_n390), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n210), .A2(G128), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n218), .A2(G143), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(new_n229), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n229), .B1(new_n396), .B2(new_n397), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n394), .B(new_n395), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n388), .A2(new_n390), .ZN(new_n402));
  INV_X1    g216(.A(new_n273), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n395), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT96), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n398), .A2(KEYINPUT95), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT95), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n396), .A2(new_n397), .A3(new_n408), .A4(new_n229), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n396), .A2(new_n397), .A3(KEYINPUT13), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n218), .A2(G143), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT13), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n229), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n407), .A2(new_n409), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n405), .A2(new_n406), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n406), .B1(new_n405), .B2(new_n414), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n401), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G217), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n187), .A2(new_n418), .A3(G953), .ZN(new_n419));
  XOR2_X1   g233(.A(new_n419), .B(KEYINPUT97), .Z(new_n420));
  NAND2_X1  g234(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n395), .B1(new_n399), .B2(new_n400), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(G107), .B2(new_n393), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n388), .A2(new_n273), .A3(new_n390), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n273), .B1(new_n388), .B2(new_n390), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n407), .A2(new_n409), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n413), .A2(new_n410), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(KEYINPUT96), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n405), .A2(new_n406), .A3(new_n414), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n423), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n420), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(G902), .B1(new_n421), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G478), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n435), .B1(KEYINPUT15), .B2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n417), .A2(new_n420), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n432), .A2(new_n433), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n309), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n436), .A2(KEYINPUT15), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G952), .ZN(new_n444));
  AOI211_X1 g258(.A(G953), .B(new_n444), .C1(G234), .C2(G237), .ZN(new_n445));
  NAND2_X1  g259(.A1(G234), .A2(G237), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(G902), .A3(G953), .ZN(new_n447));
  XOR2_X1   g261(.A(new_n447), .B(KEYINPUT98), .Z(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(G898), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n445), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n382), .A2(new_n443), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n317), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT66), .ZN(new_n453));
  OAI21_X1  g267(.A(G131), .B1(new_n226), .B2(G134), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n454), .B1(G134), .B2(new_n226), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(new_n240), .B2(new_n326), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n453), .B1(new_n456), .B2(new_n220), .ZN(new_n457));
  AOI21_X1  g271(.A(G131), .B1(new_n231), .B2(new_n235), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n222), .B(KEYINPUT66), .C1(new_n458), .C2(new_n455), .ZN(new_n459));
  INV_X1    g273(.A(new_n282), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n237), .B2(new_n238), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n457), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT2), .B(G113), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(G116), .B(G119), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT68), .ZN(new_n466));
  OAI21_X1  g280(.A(KEYINPUT69), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NOR3_X1   g282(.A1(new_n465), .A2(new_n466), .A3(KEYINPUT69), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n464), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n469), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(new_n463), .A3(new_n467), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n462), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n239), .A2(new_n244), .A3(new_n286), .ZN(new_n476));
  INV_X1    g290(.A(new_n267), .ZN(new_n477));
  OAI22_X1  g291(.A1(new_n477), .A2(new_n265), .B1(new_n458), .B2(new_n455), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n476), .A2(new_n478), .A3(new_n473), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  XOR2_X1   g294(.A(KEYINPUT74), .B(KEYINPUT28), .Z(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT75), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT28), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n479), .A2(KEYINPUT76), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT76), .B1(new_n479), .B2(new_n485), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT75), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n480), .A2(new_n489), .A3(new_n482), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n322), .A2(G210), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(KEYINPUT27), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT26), .B(G101), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n492), .B(new_n493), .ZN(new_n494));
  XOR2_X1   g308(.A(new_n494), .B(KEYINPUT73), .Z(new_n495));
  NAND4_X1  g309(.A1(new_n484), .A2(new_n488), .A3(new_n490), .A4(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT30), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n462), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT67), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n476), .A2(KEYINPUT30), .A3(new_n478), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n462), .A2(KEYINPUT67), .A3(new_n497), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n500), .A2(new_n474), .A3(new_n501), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n479), .ZN(new_n504));
  INV_X1    g318(.A(new_n494), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT29), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n496), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n476), .A2(new_n478), .A3(new_n473), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n473), .B1(new_n476), .B2(new_n478), .ZN(new_n510));
  OAI21_X1  g324(.A(KEYINPUT28), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT77), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g327(.A(KEYINPUT77), .B(KEYINPUT28), .C1(new_n509), .C2(new_n510), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n505), .A2(new_n507), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n488), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n309), .ZN(new_n518));
  OAI21_X1  g332(.A(G472), .B1(new_n508), .B2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT32), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n509), .A2(new_n505), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n503), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT31), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n503), .A2(KEYINPUT31), .A3(new_n521), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n484), .A2(new_n488), .A3(new_n490), .ZN(new_n526));
  INV_X1    g340(.A(new_n495), .ZN(new_n527));
  AOI22_X1  g341(.A1(new_n524), .A2(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(G472), .A2(G902), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n520), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT76), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n532), .B1(new_n509), .B2(KEYINPUT28), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n479), .A2(KEYINPUT76), .A3(new_n485), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n489), .B1(new_n480), .B2(new_n482), .ZN(new_n536));
  AOI211_X1 g350(.A(KEYINPUT75), .B(new_n481), .C1(new_n475), .C2(new_n479), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n503), .A2(KEYINPUT31), .A3(new_n521), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT31), .B1(new_n503), .B2(new_n521), .ZN(new_n540));
  OAI22_X1  g354(.A1(new_n538), .A2(new_n495), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n530), .A2(new_n520), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n519), .A2(new_n531), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n418), .B1(G234), .B2(new_n309), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT79), .ZN(new_n547));
  XOR2_X1   g361(.A(KEYINPUT24), .B(G110), .Z(new_n548));
  XNOR2_X1  g362(.A(G119), .B(G128), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n336), .B2(new_n337), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT23), .ZN(new_n552));
  INV_X1    g366(.A(G119), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n552), .B1(new_n553), .B2(G128), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n218), .A2(KEYINPUT23), .A3(G119), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(G128), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT78), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT78), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n554), .A2(new_n555), .A3(new_n559), .A4(new_n556), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n558), .A2(G110), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n547), .B1(new_n551), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n333), .A2(new_n334), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n213), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n335), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n566), .A2(KEYINPUT79), .A3(new_n561), .A4(new_n550), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n355), .A2(new_n335), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n557), .A2(G110), .ZN(new_n570));
  OR2_X1    g384(.A1(new_n570), .A2(KEYINPUT80), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n548), .A2(new_n549), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n572), .B1(new_n570), .B2(KEYINPUT80), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n569), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n568), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n290), .A2(G221), .A3(G234), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(KEYINPUT82), .ZN(new_n578));
  XOR2_X1   g392(.A(KEYINPUT22), .B(G137), .Z(new_n579));
  OR2_X1    g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n579), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n576), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n582), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n568), .A2(new_n575), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n583), .A2(new_n309), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT83), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(KEYINPUT25), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  AOI211_X1 g403(.A(new_n582), .B(new_n574), .C1(new_n563), .C2(new_n567), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n584), .B1(new_n568), .B2(new_n575), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n588), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n309), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n546), .B1(new_n589), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n545), .A2(G902), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(G214), .B1(G237), .B2(G902), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n465), .A2(KEYINPUT5), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n386), .A2(KEYINPUT5), .A3(G119), .ZN(new_n601));
  INV_X1    g415(.A(G113), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI22_X1  g417(.A1(new_n600), .A2(new_n603), .B1(new_n464), .B2(new_n465), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n254), .A2(new_n263), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n474), .A2(new_n278), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(G110), .B(G122), .ZN(new_n608));
  XOR2_X1   g422(.A(new_n608), .B(KEYINPUT90), .Z(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n605), .A2(new_n606), .A3(new_n609), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(KEYINPUT6), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT6), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n607), .A2(new_n614), .A3(new_n610), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n222), .A2(new_n331), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n616), .B1(new_n331), .B2(new_n282), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n290), .A2(G224), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(KEYINPUT91), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n617), .B(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n613), .A2(new_n615), .A3(new_n620), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n618), .A2(KEYINPUT7), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n617), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n209), .A2(new_n604), .ZN(new_n624));
  XOR2_X1   g438(.A(new_n609), .B(KEYINPUT8), .Z(new_n625));
  NOR3_X1   g439(.A1(new_n604), .A2(new_n255), .A3(new_n260), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n623), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(G902), .B1(new_n628), .B2(new_n612), .ZN(new_n629));
  OAI21_X1  g443(.A(G210), .B1(G237), .B2(G902), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n621), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n630), .B1(new_n621), .B2(new_n629), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n599), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n544), .A2(new_n598), .A3(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n452), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(new_n256), .ZN(G3));
  INV_X1    g451(.A(G472), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n541), .B2(new_n309), .ZN(new_n639));
  INV_X1    g453(.A(new_n598), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n524), .A2(new_n525), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n526), .A2(new_n527), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n530), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n639), .A2(new_n640), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT33), .B1(new_n421), .B2(new_n434), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n436), .A2(G902), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT33), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n417), .A2(KEYINPUT99), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n648), .B1(new_n649), .B2(new_n433), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n417), .A2(KEYINPUT99), .A3(new_n420), .ZN(new_n651));
  AOI21_X1  g465(.A(KEYINPUT100), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT99), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n433), .B1(new_n432), .B2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n654), .A2(new_n651), .A3(KEYINPUT100), .A4(KEYINPUT33), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  OAI211_X1 g470(.A(new_n646), .B(new_n647), .C1(new_n652), .C2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT101), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n440), .A2(new_n658), .A3(new_n436), .ZN(new_n659));
  OAI21_X1  g473(.A(KEYINPUT101), .B1(new_n435), .B2(G478), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n450), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n662), .A2(new_n663), .A3(new_n382), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n633), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n317), .A2(new_n644), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT34), .B(G104), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT103), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n668), .B(KEYINPUT102), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n666), .B(new_n669), .ZN(G6));
  NAND2_X1  g484(.A1(new_n377), .A2(new_n378), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT20), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n377), .A2(new_n365), .A3(new_n378), .ZN(new_n673));
  AOI22_X1  g487(.A1(new_n672), .A2(new_n673), .B1(G475), .B2(new_n363), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n674), .A2(new_n663), .A3(new_n443), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT104), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n317), .A2(new_n644), .A3(new_n634), .A4(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT35), .B(G107), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G9));
  NOR2_X1   g493(.A1(new_n639), .A2(new_n643), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n582), .A2(KEYINPUT36), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n576), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n568), .A2(new_n575), .A3(new_n681), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n596), .A3(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n683), .A2(KEYINPUT105), .A3(new_n596), .A4(new_n684), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(KEYINPUT106), .B1(new_n595), .B2(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n593), .B1(new_n592), .B2(new_n309), .ZN(new_n691));
  NOR4_X1   g505(.A1(new_n590), .A2(new_n591), .A3(G902), .A4(new_n588), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n545), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n687), .A2(new_n688), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n690), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n633), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n317), .A2(new_n451), .A3(new_n680), .A4(new_n698), .ZN(new_n699));
  XOR2_X1   g513(.A(KEYINPUT37), .B(G110), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G12));
  INV_X1    g515(.A(new_n443), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n382), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(G900), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n445), .B1(new_n448), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n317), .A2(new_n544), .A3(new_n698), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G128), .ZN(G30));
  XOR2_X1   g523(.A(new_n706), .B(KEYINPUT39), .Z(new_n710));
  NAND2_X1  g524(.A1(new_n317), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g525(.A1(new_n711), .A2(KEYINPUT40), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(KEYINPUT40), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n621), .A2(new_n629), .ZN(new_n714));
  INV_X1    g528(.A(new_n630), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n621), .A2(new_n629), .A3(new_n630), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(KEYINPUT38), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n527), .B1(new_n509), .B2(new_n510), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n522), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n638), .B1(new_n721), .B2(new_n309), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n541), .B2(new_n542), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n531), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n382), .A2(new_n443), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n595), .A2(new_n689), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n599), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AND4_X1   g543(.A1(new_n719), .A2(new_n724), .A3(new_n725), .A4(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n712), .A2(new_n713), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G143), .ZN(G45));
  NAND3_X1  g546(.A1(new_n654), .A2(new_n651), .A3(KEYINPUT33), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT100), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n645), .B1(new_n735), .B2(new_n655), .ZN(new_n736));
  AOI22_X1  g550(.A1(new_n736), .A2(new_n647), .B1(new_n660), .B2(new_n659), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT107), .ZN(new_n738));
  NOR4_X1   g552(.A1(new_n737), .A2(new_n738), .A3(new_n674), .A4(new_n706), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n674), .B1(new_n657), .B2(new_n661), .ZN(new_n740));
  INV_X1    g554(.A(new_n706), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT107), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(new_n317), .A3(new_n544), .A4(new_n698), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G146), .ZN(G48));
  INV_X1    g559(.A(KEYINPUT109), .ZN(new_n746));
  AND4_X1   g560(.A1(new_n304), .A2(new_n299), .A3(new_n246), .A4(new_n300), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n304), .B1(new_n303), .B2(new_n300), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n312), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n295), .ZN(new_n750));
  AOI21_X1  g564(.A(G902), .B1(new_n750), .B2(new_n297), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n189), .B1(new_n751), .B2(new_n308), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT108), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n307), .A2(new_n309), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n753), .B1(new_n754), .B2(G469), .ZN(new_n755));
  AOI211_X1 g569(.A(KEYINPUT108), .B(new_n308), .C1(new_n307), .C2(new_n309), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n752), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n544), .A2(new_n598), .A3(new_n665), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n746), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n544), .A2(new_n598), .A3(new_n665), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n310), .A2(new_n188), .ZN(new_n761));
  OAI21_X1  g575(.A(KEYINPUT108), .B1(new_n751), .B2(new_n308), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n754), .A2(new_n753), .A3(G469), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n760), .A2(new_n764), .A3(KEYINPUT109), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n759), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(KEYINPUT41), .B(G113), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n766), .B(new_n767), .ZN(G15));
  OAI211_X1 g582(.A(new_n634), .B(new_n752), .C1(new_n755), .C2(new_n756), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n544), .A2(new_n676), .A3(new_n598), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n386), .ZN(G18));
  INV_X1    g586(.A(new_n697), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n544), .A2(new_n451), .A3(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n553), .ZN(G21));
  NAND2_X1  g590(.A1(new_n762), .A2(new_n763), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n539), .A2(new_n540), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n495), .B1(new_n515), .B2(new_n488), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n529), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(G902), .B1(new_n641), .B2(new_n642), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n780), .B(new_n598), .C1(new_n781), .C2(new_n638), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n718), .A2(new_n663), .A3(new_n599), .A4(new_n725), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n777), .A2(new_n752), .A3(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G122), .ZN(G24));
  OAI211_X1 g600(.A(new_n727), .B(new_n780), .C1(new_n781), .C2(new_n638), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n787), .A2(new_n739), .A3(new_n742), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n764), .A2(new_n788), .A3(new_n634), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G125), .ZN(G27));
  INV_X1    g604(.A(new_n542), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT110), .B1(new_n528), .B2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT110), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n541), .A2(new_n793), .A3(new_n542), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n519), .A2(new_n531), .A3(new_n792), .A4(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n743), .A2(new_n795), .A3(new_n598), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n718), .A2(new_n728), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n317), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT42), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n310), .A2(new_n316), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n800), .A2(new_n188), .A3(new_n797), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n544), .A2(new_n598), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT42), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n801), .A2(new_n802), .A3(new_n803), .A4(new_n743), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n799), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(new_n326), .ZN(G33));
  NAND3_X1  g620(.A1(new_n801), .A2(new_n802), .A3(new_n707), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G134), .ZN(G36));
  INV_X1    g622(.A(KEYINPUT45), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n314), .A2(new_n296), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n809), .B1(new_n810), .B2(new_n313), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n315), .A2(KEYINPUT45), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(G469), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n811), .A2(KEYINPUT111), .A3(new_n812), .A4(G469), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n311), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n817), .A2(KEYINPUT46), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(KEYINPUT46), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n310), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n820), .A2(new_n188), .A3(new_n710), .ZN(new_n821));
  INV_X1    g635(.A(new_n821), .ZN(new_n822));
  AOI211_X1 g636(.A(KEYINPUT43), .B(new_n382), .C1(new_n662), .C2(KEYINPUT112), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n662), .A2(KEYINPUT112), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n674), .B(KEYINPUT113), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n662), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT43), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n680), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(KEYINPUT44), .A3(new_n830), .A4(new_n727), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT44), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n825), .A2(new_n828), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n830), .A2(new_n727), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n832), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n831), .A2(new_n797), .A3(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(KEYINPUT114), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n822), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(G137), .ZN(G39));
  INV_X1    g653(.A(new_n797), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n544), .A2(new_n840), .A3(new_n598), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT47), .B1(new_n820), .B2(new_n188), .ZN(new_n842));
  INV_X1    g656(.A(new_n819), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n310), .B1(new_n817), .B2(KEYINPUT46), .ZN(new_n844));
  OAI211_X1 g658(.A(KEYINPUT47), .B(new_n188), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n743), .B(new_n841), .C1(new_n842), .C2(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(G140), .ZN(G42));
  NAND2_X1  g662(.A1(new_n777), .A2(new_n310), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n849), .A2(KEYINPUT49), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(KEYINPUT49), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n598), .A2(new_n188), .A3(new_n599), .ZN(new_n852));
  NOR4_X1   g666(.A1(new_n719), .A2(new_n827), .A3(new_n724), .A4(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n850), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n795), .A2(new_n598), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n764), .A2(new_n797), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n825), .A2(new_n828), .A3(new_n445), .ZN(new_n857));
  OR3_X1    g671(.A1(new_n856), .A2(KEYINPUT122), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT122), .B1(new_n856), .B2(new_n857), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n855), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  XOR2_X1   g674(.A(new_n860), .B(KEYINPUT48), .Z(new_n861));
  INV_X1    g675(.A(new_n782), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n829), .A2(new_n445), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n769), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n864), .A2(new_n444), .A3(G953), .ZN(new_n865));
  INV_X1    g679(.A(new_n740), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n598), .A2(new_n445), .ZN(new_n867));
  OR3_X1    g681(.A1(new_n856), .A2(new_n724), .A3(new_n867), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n861), .B(new_n865), .C1(new_n866), .C2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT50), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n719), .A2(new_n599), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n764), .ZN(new_n872));
  OR3_X1    g686(.A1(new_n863), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n870), .B1(new_n863), .B2(new_n872), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n873), .A2(KEYINPUT121), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT121), .B1(new_n873), .B2(new_n874), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n787), .B1(new_n858), .B2(new_n859), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  OR3_X1    g693(.A1(new_n868), .A2(new_n382), .A3(new_n662), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n877), .A2(new_n881), .A3(KEYINPUT51), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n883), .B1(new_n842), .B2(new_n846), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n188), .B1(new_n843), .B2(new_n844), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT47), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n887), .A2(KEYINPUT119), .A3(new_n845), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n188), .B1(new_n849), .B2(KEYINPUT120), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(KEYINPUT120), .B2(new_n849), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n884), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n863), .A2(new_n840), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n882), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n879), .A2(new_n880), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n873), .A2(new_n874), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n868), .A2(new_n382), .A3(new_n662), .ZN(new_n898));
  OAI21_X1  g712(.A(KEYINPUT123), .B1(new_n898), .B2(new_n878), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n842), .A2(new_n846), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n893), .B1(new_n901), .B2(new_n890), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT51), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n869), .B1(new_n894), .B2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT53), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n789), .A2(new_n708), .A3(new_n744), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n726), .A2(new_n741), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n531), .B2(new_n723), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n725), .B(new_n599), .C1(new_n631), .C2(new_n632), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n317), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT52), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT116), .B1(new_n906), .B2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(new_n744), .ZN(new_n914));
  INV_X1    g728(.A(new_n708), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT116), .ZN(new_n917));
  INV_X1    g731(.A(new_n912), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n916), .A2(new_n917), .A3(new_n789), .A4(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT52), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n744), .A2(new_n708), .A3(new_n911), .ZN(new_n921));
  INV_X1    g735(.A(new_n787), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n743), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n769), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n920), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n913), .A2(new_n919), .A3(new_n925), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n382), .A2(new_n443), .A3(new_n706), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n927), .A2(new_n599), .A3(new_n716), .A4(new_n717), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT115), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n631), .A2(new_n632), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n931), .A2(KEYINPUT115), .A3(new_n599), .A4(new_n927), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n933), .A2(new_n317), .A3(new_n544), .A4(new_n773), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n743), .A2(new_n922), .A3(new_n317), .A4(new_n797), .ZN(new_n935));
  INV_X1    g749(.A(new_n707), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n317), .A2(new_n544), .A3(new_n598), .A4(new_n797), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n934), .B(new_n935), .C1(new_n936), .C2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n805), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n666), .B1(new_n452), .B2(new_n635), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n771), .A2(new_n775), .A3(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n633), .A2(new_n675), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n317), .A2(new_n644), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n785), .A2(new_n699), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n759), .B2(new_n765), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n939), .A2(new_n941), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n905), .B1(new_n926), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n771), .A2(new_n940), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n785), .A2(new_n699), .A3(new_n943), .ZN(new_n949));
  INV_X1    g763(.A(new_n775), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n948), .A2(new_n766), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n934), .A2(new_n935), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n952), .A2(new_n799), .A3(new_n807), .A4(new_n804), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n544), .A2(new_n698), .A3(new_n707), .ZN(new_n955));
  INV_X1    g769(.A(new_n907), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n724), .A2(new_n910), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n317), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n958), .A2(KEYINPUT52), .A3(new_n789), .A4(new_n744), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT117), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n925), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n925), .A2(new_n959), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(KEYINPUT117), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n954), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n947), .B1(new_n905), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(KEYINPUT54), .ZN(new_n966));
  AOI21_X1  g780(.A(KEYINPUT118), .B1(new_n964), .B2(new_n905), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT54), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n913), .A2(new_n919), .A3(new_n925), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n954), .A2(new_n970), .A3(KEYINPUT53), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n964), .A2(KEYINPUT118), .A3(new_n905), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n968), .A2(new_n969), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n904), .A2(new_n966), .A3(new_n973), .ZN(new_n974));
  NOR2_X1   g788(.A1(G952), .A2(G953), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n854), .B1(new_n974), .B2(new_n975), .ZN(G75));
  NAND2_X1  g790(.A1(new_n972), .A2(new_n971), .ZN(new_n977));
  OAI211_X1 g791(.A(G210), .B(G902), .C1(new_n977), .C2(new_n967), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT56), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n613), .A2(new_n615), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(new_n620), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT55), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n978), .A2(new_n979), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n982), .B1(new_n978), .B2(new_n979), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n290), .A2(G952), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(G51));
  XNOR2_X1  g800(.A(new_n311), .B(KEYINPUT57), .ZN(new_n987));
  INV_X1    g801(.A(new_n971), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n960), .B1(new_n925), .B2(new_n959), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n946), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(KEYINPUT53), .B1(new_n990), .B2(new_n961), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n988), .B1(new_n991), .B2(KEYINPUT118), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n969), .B1(new_n992), .B2(new_n968), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n977), .A2(KEYINPUT54), .A3(new_n967), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n987), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n307), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n992), .A2(new_n968), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n997), .A2(G902), .A3(new_n815), .A4(new_n816), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n985), .B1(new_n996), .B2(new_n998), .ZN(G54));
  AND2_X1   g813(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n997), .A2(G902), .A3(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n1001), .A2(new_n376), .A3(new_n375), .ZN(new_n1002));
  INV_X1    g816(.A(new_n985), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n997), .A2(G902), .A3(new_n377), .A4(new_n1000), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(G60));
  NAND2_X1  g819(.A1(new_n973), .A2(new_n966), .ZN(new_n1006));
  NAND2_X1  g820(.A1(G478), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT59), .Z(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n736), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n736), .A2(new_n1009), .ZN(new_n1011));
  OAI21_X1  g825(.A(KEYINPUT54), .B1(new_n977), .B2(new_n967), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1011), .B1(new_n1012), .B2(new_n973), .ZN(new_n1013));
  NOR3_X1   g827(.A1(new_n1010), .A2(new_n985), .A3(new_n1013), .ZN(G63));
  AND2_X1   g828(.A1(new_n683), .A2(new_n684), .ZN(new_n1015));
  NAND2_X1  g829(.A1(G217), .A2(G902), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1016), .B(KEYINPUT60), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n1015), .B(new_n1018), .C1(new_n977), .C2(new_n967), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1017), .B1(new_n992), .B2(new_n968), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n1003), .B(new_n1019), .C1(new_n1020), .C2(new_n592), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT61), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n977), .A2(new_n967), .ZN(new_n1024));
  OAI22_X1  g838(.A1(new_n1024), .A2(new_n1017), .B1(new_n590), .B2(new_n591), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n1025), .A2(KEYINPUT61), .A3(new_n1003), .A4(new_n1019), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1023), .A2(new_n1026), .ZN(G66));
  INV_X1    g841(.A(G224), .ZN(new_n1028));
  OAI21_X1  g842(.A(G953), .B1(new_n449), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g843(.A(new_n951), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1029), .B1(new_n1030), .B2(G953), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n980), .B1(G898), .B2(new_n290), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1031), .B(new_n1032), .ZN(G69));
  AOI21_X1  g847(.A(new_n290), .B1(G227), .B2(G900), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1035), .B(new_n370), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1036), .ZN(new_n1037));
  INV_X1    g851(.A(new_n906), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1038), .A2(new_n731), .ZN(new_n1039));
  XOR2_X1   g853(.A(new_n1039), .B(KEYINPUT62), .Z(new_n1040));
  AOI21_X1  g854(.A(new_n840), .B1(new_n866), .B2(new_n704), .ZN(new_n1041));
  NAND4_X1  g855(.A1(new_n1041), .A2(new_n802), .A3(new_n317), .A4(new_n710), .ZN(new_n1042));
  NAND4_X1  g856(.A1(new_n1040), .A2(new_n838), .A3(new_n847), .A4(new_n1042), .ZN(new_n1043));
  AOI21_X1  g857(.A(new_n1037), .B1(new_n1043), .B2(new_n290), .ZN(new_n1044));
  INV_X1    g858(.A(KEYINPUT124), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g860(.A(new_n1046), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1036), .B1(G900), .B2(G953), .ZN(new_n1048));
  NOR2_X1   g862(.A1(new_n855), .A2(new_n909), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n822), .B1(new_n837), .B2(new_n1049), .ZN(new_n1050));
  AND4_X1   g864(.A1(new_n799), .A2(new_n1038), .A3(new_n804), .A4(new_n807), .ZN(new_n1051));
  NAND3_X1  g865(.A1(new_n1050), .A2(new_n847), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1048), .B1(new_n1052), .B2(G953), .ZN(new_n1053));
  OAI21_X1  g867(.A(new_n1053), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1054));
  OAI21_X1  g868(.A(new_n1034), .B1(new_n1047), .B2(new_n1054), .ZN(new_n1055));
  OR2_X1    g869(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1056));
  INV_X1    g870(.A(new_n1034), .ZN(new_n1057));
  NAND4_X1  g871(.A1(new_n1056), .A2(new_n1057), .A3(new_n1046), .A4(new_n1053), .ZN(new_n1058));
  NAND2_X1  g872(.A1(new_n1055), .A2(new_n1058), .ZN(G72));
  NOR2_X1   g873(.A1(new_n504), .A2(new_n494), .ZN(new_n1060));
  AOI21_X1  g874(.A(new_n505), .B1(new_n503), .B2(new_n479), .ZN(new_n1061));
  XNOR2_X1  g875(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1062));
  NOR2_X1   g876(.A1(new_n638), .A2(new_n309), .ZN(new_n1063));
  XOR2_X1   g877(.A(new_n1062), .B(new_n1063), .Z(new_n1064));
  INV_X1    g878(.A(new_n1064), .ZN(new_n1065));
  NOR3_X1   g879(.A1(new_n1060), .A2(new_n1061), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g880(.A1(new_n965), .A2(new_n1066), .ZN(new_n1067));
  XNOR2_X1  g881(.A(new_n1067), .B(KEYINPUT127), .ZN(new_n1068));
  OAI21_X1  g882(.A(new_n1064), .B1(new_n1043), .B2(new_n951), .ZN(new_n1069));
  NAND2_X1  g883(.A1(new_n1069), .A2(new_n1061), .ZN(new_n1070));
  OAI21_X1  g884(.A(new_n1064), .B1(new_n1052), .B2(new_n951), .ZN(new_n1071));
  XOR2_X1   g885(.A(new_n1060), .B(KEYINPUT126), .Z(new_n1072));
  AOI21_X1  g886(.A(new_n985), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  AND3_X1   g887(.A1(new_n1068), .A2(new_n1070), .A3(new_n1073), .ZN(G57));
endmodule


