//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1258, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  INV_X1    g0015(.A(G58), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(new_n210), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n212), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n215), .B(new_n223), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G226), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT65), .ZN(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT66), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(new_n217), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT12), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n221), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(KEYINPUT69), .B1(new_n210), .B2(G1), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT69), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(new_n209), .A3(G20), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n254), .B1(new_n217), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT73), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n263), .B(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n210), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(G77), .ZN(new_n267));
  OAI22_X1  g0067(.A1(new_n266), .A2(new_n267), .B1(new_n210), .B2(G68), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n210), .A2(new_n269), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n270), .A2(new_n202), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n256), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n272), .B(KEYINPUT11), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n265), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G169), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n269), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n279), .A2(G232), .A3(G1698), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G97), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G226), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n280), .B(new_n281), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT67), .ZN(new_n288));
  INV_X1    g0088(.A(G45), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G41), .ZN(new_n291));
  NAND2_X1  g0091(.A1(KEYINPUT67), .A2(G45), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n209), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT68), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n293), .A2(KEYINPUT68), .A3(new_n209), .ZN(new_n297));
  INV_X1    g0097(.A(G274), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n286), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n296), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n286), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G238), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n287), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT13), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT13), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n287), .A2(new_n307), .A3(new_n300), .A4(new_n304), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n275), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT14), .ZN(new_n310));
  AND2_X1   g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n306), .A2(G179), .A3(new_n308), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(new_n309), .B2(new_n310), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n274), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n265), .A2(new_n273), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n306), .A2(new_n308), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G190), .ZN(new_n317));
  INV_X1    g0117(.A(G200), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n315), .B(new_n317), .C1(new_n316), .C2(new_n318), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  AND2_X1   g0120(.A1(G58), .A2(G68), .ZN(new_n321));
  OAI21_X1  g0121(.A(G20), .B1(new_n321), .B2(new_n201), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT74), .ZN(new_n323));
  NOR2_X1   g0123(.A1(G20), .A2(G33), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G159), .ZN(new_n325));
  AND3_X1   g0125(.A1(new_n322), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n323), .B1(new_n322), .B2(new_n325), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n277), .A2(new_n210), .A3(new_n278), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT7), .ZN(new_n330));
  AND2_X1   g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  NOR2_X1   g0131(.A1(KEYINPUT3), .A2(G33), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT7), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n333), .A2(new_n334), .A3(new_n210), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n330), .A2(new_n335), .A3(G68), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n328), .B(new_n336), .C1(KEYINPUT75), .C2(KEYINPUT16), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT16), .ZN(new_n338));
  NAND2_X1  g0138(.A1(G58), .A2(G68), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n210), .B1(new_n218), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G159), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n270), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(KEYINPUT74), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n322), .A2(new_n323), .A3(new_n325), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n343), .A2(KEYINPUT75), .A3(new_n344), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n330), .A2(new_n335), .A3(G68), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n344), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n338), .B(new_n345), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n337), .A2(new_n348), .A3(new_n256), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT8), .B(G58), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(new_n252), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(new_n262), .B2(new_n351), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n297), .A2(new_n299), .ZN(new_n356));
  AOI21_X1  g0156(.A(KEYINPUT68), .B1(new_n293), .B2(new_n209), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n301), .A2(G232), .A3(new_n302), .ZN(new_n359));
  NOR2_X1   g0159(.A1(G223), .A2(G1698), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n284), .B2(G1698), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n361), .A2(new_n279), .B1(G33), .B2(G87), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n359), .B1(new_n362), .B2(new_n301), .ZN(new_n363));
  OAI21_X1  g0163(.A(G169), .B1(new_n358), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n361), .A2(new_n279), .ZN(new_n365));
  NAND2_X1  g0165(.A1(G33), .A2(G87), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n286), .ZN(new_n368));
  XNOR2_X1  g0168(.A(KEYINPUT71), .B(G179), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n300), .A2(new_n368), .A3(new_n370), .A4(new_n359), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n364), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n355), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT18), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT18), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n355), .A2(new_n375), .A3(new_n372), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT17), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n318), .B1(new_n358), .B2(new_n363), .ZN(new_n379));
  INV_X1    g0179(.A(G190), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n300), .A2(new_n368), .A3(new_n380), .A4(new_n359), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n349), .A2(new_n382), .A3(new_n354), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(KEYINPUT76), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT76), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n349), .A2(new_n382), .A3(new_n385), .A4(new_n354), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n378), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n383), .A2(new_n378), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n377), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n279), .A2(G222), .A3(new_n282), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n279), .A2(G223), .A3(G1698), .ZN(new_n391));
  OAI211_X1 g0191(.A(new_n390), .B(new_n391), .C1(new_n267), .C2(new_n279), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n392), .A2(new_n286), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n303), .A2(G226), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n300), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(G200), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n324), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n397), .B1(new_n350), .B2(new_n266), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n398), .A2(new_n256), .B1(new_n202), .B2(new_n252), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n202), .B1(new_n258), .B2(new_n260), .ZN(new_n400));
  OR2_X1    g0200(.A1(new_n400), .A2(KEYINPUT70), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(KEYINPUT70), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n401), .A2(new_n257), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT9), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n392), .A2(new_n286), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n407), .A2(new_n300), .A3(G190), .A4(new_n394), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n399), .A2(new_n403), .A3(KEYINPUT9), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n396), .A2(new_n406), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT10), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n411), .B1(new_n396), .B2(KEYINPUT72), .ZN(new_n412));
  OR2_X1    g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n410), .A2(new_n412), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n303), .A2(G244), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n279), .A2(G238), .A3(G1698), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n279), .A2(G232), .A3(new_n282), .ZN(new_n418));
  OAI211_X1 g0218(.A(new_n417), .B(new_n418), .C1(new_n206), .C2(new_n279), .ZN(new_n419));
  AOI211_X1 g0219(.A(new_n416), .B(new_n358), .C1(new_n286), .C2(new_n419), .ZN(new_n420));
  OR2_X1    g0220(.A1(new_n420), .A2(G169), .ZN(new_n421));
  XNOR2_X1  g0221(.A(KEYINPUT15), .B(G87), .ZN(new_n422));
  OAI22_X1  g0222(.A1(new_n422), .A2(new_n266), .B1(new_n210), .B2(new_n267), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n350), .A2(new_n270), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n256), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n252), .A2(new_n267), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n425), .B(new_n426), .C1(new_n267), .C2(new_n262), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n420), .A2(new_n369), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n421), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n395), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(new_n369), .A3(new_n407), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n275), .B1(new_n395), .B2(new_n393), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(new_n404), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n427), .B1(new_n420), .B2(G190), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n318), .B2(new_n420), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n429), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n320), .A2(new_n389), .A3(new_n415), .A4(new_n436), .ZN(new_n437));
  XNOR2_X1  g0237(.A(new_n437), .B(KEYINPUT77), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT82), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT81), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n209), .B(G45), .C1(new_n291), .C2(KEYINPUT5), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT79), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n289), .A2(G1), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT5), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(G41), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(KEYINPUT79), .A3(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT80), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n445), .B2(G41), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n291), .A2(KEYINPUT80), .A3(KEYINPUT5), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n443), .A2(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G257), .ZN(new_n452));
  NOR3_X1   g0252(.A1(new_n451), .A2(new_n452), .A3(new_n286), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n443), .A2(new_n447), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n449), .A2(new_n450), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(new_n299), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n440), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n441), .A2(new_n442), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT79), .B1(new_n444), .B2(new_n446), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n455), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n461), .A2(G257), .A3(new_n301), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n462), .A2(KEYINPUT81), .A3(new_n456), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT4), .ZN(new_n464));
  INV_X1    g0264(.A(G244), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n464), .B1(new_n283), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n279), .A2(G250), .A3(G1698), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n279), .A2(KEYINPUT4), .A3(G244), .A4(new_n282), .ZN(new_n468));
  NAND2_X1  g0268(.A1(G33), .A2(G283), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n466), .A2(new_n467), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n286), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n458), .A2(G190), .A3(new_n463), .A4(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n269), .A2(G1), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n252), .A2(new_n256), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G97), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(G97), .B2(new_n251), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT6), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n477), .A2(new_n205), .A3(G107), .ZN(new_n478));
  XNOR2_X1  g0278(.A(G97), .B(G107), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n478), .B1(new_n477), .B2(new_n479), .ZN(new_n480));
  OAI221_X1 g0280(.A(KEYINPUT78), .B1(new_n267), .B2(new_n270), .C1(new_n480), .C2(new_n210), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT78), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(new_n477), .ZN(new_n483));
  INV_X1    g0283(.A(new_n478), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n210), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n270), .A2(new_n267), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n482), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n330), .A2(new_n335), .A3(G107), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n481), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n476), .B1(new_n489), .B2(new_n256), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n472), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n462), .A2(new_n456), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n492), .A2(new_n440), .B1(new_n286), .B2(new_n470), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n318), .B1(new_n493), .B2(new_n463), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n439), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n458), .A2(new_n463), .A3(new_n471), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(G200), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n497), .A2(KEYINPUT82), .A3(new_n490), .A4(new_n472), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n495), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n490), .B1(new_n275), .B2(new_n496), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n493), .A2(new_n369), .A3(new_n463), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AND2_X1   g0302(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n209), .A2(G45), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G250), .ZN(new_n505));
  OAI22_X1  g0305(.A1(new_n286), .A2(new_n505), .B1(new_n298), .B2(new_n504), .ZN(new_n506));
  OAI211_X1 g0306(.A(G244), .B(G1698), .C1(new_n331), .C2(new_n332), .ZN(new_n507));
  OAI211_X1 g0307(.A(G238), .B(new_n282), .C1(new_n331), .C2(new_n332), .ZN(new_n508));
  INV_X1    g0308(.A(G116), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n507), .B(new_n508), .C1(new_n269), .C2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n506), .B1(new_n510), .B2(new_n286), .ZN(new_n511));
  OR2_X1    g0311(.A1(new_n511), .A2(new_n318), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n279), .A2(new_n210), .A3(G68), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT19), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n210), .B1(new_n281), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(G87), .B2(new_n207), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n514), .B1(new_n266), .B2(new_n205), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n513), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n256), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n422), .A2(new_n252), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n474), .A2(G87), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT83), .ZN(new_n523));
  AND3_X1   g0323(.A1(new_n511), .A2(new_n523), .A3(G190), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n523), .B1(new_n511), .B2(G190), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n512), .B(new_n522), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n422), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n474), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n519), .A2(new_n520), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n511), .A2(new_n369), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n529), .B(new_n530), .C1(G169), .C2(new_n511), .ZN(new_n531));
  OAI211_X1 g0331(.A(G250), .B(new_n282), .C1(new_n331), .C2(new_n332), .ZN(new_n532));
  OAI211_X1 g0332(.A(G257), .B(G1698), .C1(new_n331), .C2(new_n332), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G294), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT85), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n532), .A2(new_n533), .A3(KEYINPUT85), .A4(new_n534), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n286), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n286), .B1(new_n454), .B2(new_n455), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(G264), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n539), .A2(new_n541), .A3(G190), .A4(new_n456), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT24), .ZN(new_n543));
  INV_X1    g0343(.A(G87), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n544), .A2(KEYINPUT84), .A3(G20), .ZN(new_n545));
  AOI21_X1  g0345(.A(KEYINPUT22), .B1(new_n279), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n210), .A2(G33), .A3(G116), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT23), .B1(new_n206), .B2(G20), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n279), .A2(KEYINPUT22), .A3(new_n545), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n543), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT22), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT84), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n555), .A2(new_n210), .A3(G87), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n554), .B1(new_n333), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT23), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n210), .B2(G107), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n269), .A2(new_n509), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n559), .A2(new_n560), .B1(new_n561), .B2(new_n210), .ZN(new_n562));
  AND4_X1   g0362(.A1(new_n543), .A2(new_n557), .A3(new_n552), .A4(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n256), .B1(new_n553), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n252), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT25), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n251), .B2(G107), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n474), .A2(G107), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n542), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n301), .B1(new_n535), .B2(new_n536), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n570), .A2(new_n538), .B1(new_n540), .B2(G264), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n318), .B1(new_n571), .B2(new_n456), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n526), .B(new_n531), .C1(new_n569), .C2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n469), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n509), .A2(G20), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n574), .A2(new_n256), .A3(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT20), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n574), .A2(KEYINPUT20), .A3(new_n256), .A4(new_n575), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n251), .A2(G116), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n474), .B2(G116), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n461), .A2(G270), .A3(new_n301), .ZN(new_n585));
  OAI211_X1 g0385(.A(G264), .B(G1698), .C1(new_n331), .C2(new_n332), .ZN(new_n586));
  OAI211_X1 g0386(.A(G257), .B(new_n282), .C1(new_n331), .C2(new_n332), .ZN(new_n587));
  INV_X1    g0387(.A(G303), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n586), .B(new_n587), .C1(new_n588), .C2(new_n279), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n286), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n585), .A2(G190), .A3(new_n590), .A4(new_n456), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n585), .A2(new_n456), .A3(new_n590), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n584), .B(new_n591), .C1(new_n592), .C2(new_n318), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n585), .A2(new_n456), .A3(new_n590), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n275), .B1(new_n580), .B2(new_n582), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT21), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n592), .A2(G179), .A3(new_n583), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n593), .A2(new_n598), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n564), .A2(new_n568), .ZN(new_n602));
  INV_X1    g0402(.A(G179), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n571), .A2(new_n603), .A3(new_n456), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n539), .A2(new_n541), .A3(new_n456), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n275), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n602), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n573), .A2(new_n601), .A3(new_n607), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n438), .A2(new_n503), .A3(new_n608), .ZN(G372));
  AND3_X1   g0409(.A1(new_n421), .A2(new_n427), .A3(new_n428), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n319), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n314), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n384), .A2(new_n386), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n388), .B1(new_n613), .B2(KEYINPUT17), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n377), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT86), .B1(new_n413), .B2(new_n414), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n413), .A2(KEYINPUT86), .A3(new_n414), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n433), .B1(new_n615), .B2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT87), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n621), .B(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n526), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n569), .A2(new_n572), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n602), .A2(new_n606), .A3(new_n604), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n499), .A2(new_n502), .A3(new_n628), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n502), .A2(KEYINPUT26), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n624), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(KEYINPUT26), .B1(new_n502), .B2(new_n624), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n531), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n438), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n623), .A2(new_n634), .ZN(G369));
  INV_X1    g0435(.A(new_n626), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n637));
  OR2_X1    g0437(.A1(new_n637), .A2(KEYINPUT27), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(KEYINPUT27), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(G213), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g0440(.A(new_n640), .B(KEYINPUT88), .Z(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(G343), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n645), .A2(new_n584), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n636), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n647), .B1(new_n601), .B2(new_n646), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n648), .A2(G330), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n627), .A2(new_n644), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n625), .B1(new_n602), .B2(new_n644), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n651), .B1(new_n652), .B2(new_n607), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n652), .A2(new_n627), .A3(new_n636), .A4(new_n645), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n651), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n657), .B(KEYINPUT89), .ZN(G399));
  INV_X1    g0458(.A(new_n213), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(G41), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NOR3_X1   g0461(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n661), .A2(G1), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n219), .B2(new_n661), .ZN(new_n664));
  XNOR2_X1  g0464(.A(new_n664), .B(KEYINPUT28), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n608), .A2(new_n499), .A3(new_n502), .A4(new_n645), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n539), .A2(new_n541), .A3(new_n511), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n667), .A2(new_n603), .A3(new_n594), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n668), .A2(KEYINPUT30), .A3(new_n463), .A4(new_n493), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT30), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n592), .A2(new_n571), .A3(G179), .A4(new_n511), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(new_n671), .B2(new_n496), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n592), .A2(new_n370), .A3(new_n511), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n673), .A2(new_n496), .A3(new_n605), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n669), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n644), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT31), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n675), .A2(KEYINPUT31), .A3(new_n644), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n666), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G330), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n645), .B1(new_n631), .B2(new_n633), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT90), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT29), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT29), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n683), .A2(new_n684), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n682), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n665), .B1(new_n689), .B2(G1), .ZN(G364));
  AND2_X1   g0490(.A1(new_n210), .A2(G13), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n209), .B1(new_n691), .B2(G45), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n660), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n648), .B2(G330), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(G330), .B2(new_n648), .ZN(new_n696));
  NOR2_X1   g0496(.A1(G13), .A2(G33), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G20), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n221), .B1(G20), .B2(new_n275), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g0501(.A(new_n701), .B(KEYINPUT92), .Z(new_n702));
  NOR2_X1   g0502(.A1(new_n659), .A2(new_n333), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n703), .A2(G355), .B1(new_n509), .B2(new_n659), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT91), .Z(new_n705));
  NOR2_X1   g0505(.A1(new_n659), .A2(new_n279), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n290), .A2(new_n292), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n706), .B1(new_n219), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n249), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n708), .B1(G45), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n702), .B1(new_n705), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n694), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n210), .A2(G190), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(new_n603), .A3(new_n318), .ZN(new_n714));
  INV_X1    g0514(.A(G329), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n318), .A2(G179), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n713), .ZN(new_n717));
  INV_X1    g0517(.A(G283), .ZN(new_n718));
  OAI22_X1  g0518(.A1(new_n714), .A2(new_n715), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n210), .A2(new_n380), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n716), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n279), .B1(new_n722), .B2(G303), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT98), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n369), .A2(new_n210), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n380), .A2(G200), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(G322), .ZN(new_n728));
  OAI22_X1  g0528(.A1(new_n723), .A2(new_n724), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n719), .B(new_n729), .C1(new_n724), .C2(new_n723), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n369), .A2(new_n210), .A3(G190), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n731), .A2(KEYINPUT93), .A3(new_n318), .ZN(new_n732));
  AOI21_X1  g0532(.A(KEYINPUT93), .B1(new_n731), .B2(new_n318), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G311), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n731), .A2(G200), .ZN(new_n736));
  XOR2_X1   g0536(.A(KEYINPUT33), .B(G317), .Z(new_n737));
  OAI221_X1 g0537(.A(new_n730), .B1(new_n734), .B2(new_n735), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n370), .A2(G200), .A3(new_n720), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n739), .A2(KEYINPUT94), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(KEYINPUT94), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n210), .B1(new_n726), .B2(new_n603), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n743), .A2(KEYINPUT95), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(KEYINPUT95), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI22_X1  g0546(.A1(new_n742), .A2(G326), .B1(G294), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT97), .ZN(new_n748));
  OAI221_X1 g0548(.A(new_n279), .B1(new_n717), .B2(new_n206), .C1(new_n544), .C2(new_n721), .ZN(new_n749));
  INV_X1    g0549(.A(new_n714), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G159), .ZN(new_n751));
  XNOR2_X1  g0551(.A(new_n751), .B(KEYINPUT32), .ZN(new_n752));
  INV_X1    g0552(.A(new_n727), .ZN(new_n753));
  AOI211_X1 g0553(.A(new_n749), .B(new_n752), .C1(G58), .C2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n736), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n742), .A2(G50), .B1(new_n755), .B2(G68), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n754), .B(new_n756), .C1(new_n267), .C2(new_n734), .ZN(new_n757));
  INV_X1    g0557(.A(new_n746), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n758), .A2(KEYINPUT96), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(KEYINPUT96), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n205), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n738), .A2(new_n748), .B1(new_n757), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n712), .B1(new_n763), .B2(new_n700), .ZN(new_n764));
  INV_X1    g0564(.A(new_n699), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n764), .B1(new_n648), .B2(new_n765), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n696), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(G396));
  NOR2_X1   g0568(.A1(new_n429), .A2(new_n644), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n644), .A2(new_n427), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n435), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n769), .B1(new_n429), .B2(new_n771), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n683), .B(new_n772), .Z(new_n773));
  OR2_X1    g0573(.A1(new_n773), .A2(new_n681), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n694), .B1(new_n773), .B2(new_n681), .ZN(new_n775));
  AND2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n700), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n698), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n333), .B1(new_n714), .B2(new_n735), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n721), .A2(new_n206), .B1(new_n717), .B2(new_n544), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n779), .B(new_n780), .C1(new_n753), .C2(G294), .ZN(new_n781));
  INV_X1    g0581(.A(new_n742), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n781), .B1(new_n718), .B2(new_n736), .C1(new_n782), .C2(new_n588), .ZN(new_n783));
  INV_X1    g0583(.A(new_n734), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n783), .B(new_n762), .C1(G116), .C2(new_n784), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n742), .A2(G137), .B1(new_n755), .B2(G150), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT99), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n784), .A2(G159), .B1(G143), .B2(new_n753), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT34), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n279), .B1(new_n721), .B2(new_n202), .ZN(new_n791));
  INV_X1    g0591(.A(G132), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n714), .A2(new_n792), .B1(new_n717), .B2(new_n217), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n791), .B(new_n793), .C1(new_n746), .C2(G58), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n785), .B1(new_n790), .B2(new_n794), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n694), .B1(G77), .B2(new_n778), .C1(new_n795), .C2(new_n777), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT100), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n772), .A2(new_n698), .ZN(new_n800));
  NOR3_X1   g0600(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n776), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G384));
  INV_X1    g0603(.A(new_n480), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n804), .A2(KEYINPUT35), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(KEYINPUT35), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n805), .A2(G116), .A3(new_n222), .A4(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT36), .Z(new_n808));
  NAND3_X1  g0608(.A1(new_n220), .A2(G77), .A3(new_n339), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n202), .A2(G68), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n209), .B(G13), .C1(new_n809), .C2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n686), .A2(new_n438), .A3(new_n688), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n623), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT38), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n355), .A2(new_n641), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n374), .A2(new_n376), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n816), .B1(new_n614), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT37), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n355), .B1(new_n372), .B2(new_n641), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n819), .B1(new_n820), .B2(new_n383), .ZN(new_n821));
  INV_X1    g0621(.A(new_n613), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n820), .A2(new_n819), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n815), .B1(new_n818), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n338), .B1(new_n346), .B2(new_n347), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n328), .A2(KEYINPUT16), .A3(new_n336), .ZN(new_n827));
  AND3_X1   g0627(.A1(new_n826), .A2(new_n827), .A3(new_n256), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n828), .A2(new_n353), .B1(new_n372), .B2(new_n641), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n384), .A2(new_n829), .A3(new_n386), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT37), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n820), .A2(new_n819), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n831), .B1(new_n613), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n641), .B1(new_n828), .B2(new_n353), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n833), .B(KEYINPUT38), .C1(new_n389), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n825), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT39), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n314), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(new_n645), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n834), .B1(new_n614), .B2(new_n817), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n822), .A2(new_n823), .B1(new_n830), .B2(KEYINPUT37), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n815), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n844), .A2(new_n835), .A3(KEYINPUT39), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n838), .A2(new_n841), .A3(new_n845), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n645), .B(new_n772), .C1(new_n631), .C2(new_n633), .ZN(new_n847));
  INV_X1    g0647(.A(new_n769), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n844), .A2(new_n835), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n274), .A2(new_n644), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n314), .A2(new_n319), .A3(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n274), .B(new_n644), .C1(new_n311), .C2(new_n313), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n849), .A2(new_n850), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n377), .A2(new_n642), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n846), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n814), .B(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(G330), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n438), .A2(new_n680), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT40), .B1(new_n844), .B2(new_n835), .ZN(new_n861));
  AND3_X1   g0661(.A1(new_n680), .A2(new_n772), .A3(new_n854), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n680), .A2(new_n772), .A3(new_n854), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(new_n835), .B2(new_n825), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT40), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n863), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n859), .B1(new_n860), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n860), .B2(new_n867), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n858), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n209), .B2(new_n691), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n858), .A2(new_n869), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n812), .B1(new_n871), .B2(new_n872), .ZN(G367));
  INV_X1    g0673(.A(new_n761), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(G68), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n784), .A2(G50), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n755), .A2(G159), .ZN(new_n877));
  AOI22_X1  g0677(.A1(G137), .A2(new_n750), .B1(new_n722), .B2(G58), .ZN(new_n878));
  INV_X1    g0678(.A(new_n717), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n333), .B1(new_n879), .B2(G77), .ZN(new_n880));
  INV_X1    g0680(.A(G150), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n878), .B(new_n880), .C1(new_n727), .C2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(G143), .B2(new_n742), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n875), .A2(new_n876), .A3(new_n877), .A4(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n721), .A2(new_n509), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT46), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n727), .A2(new_n588), .ZN(new_n887));
  INV_X1    g0687(.A(G317), .ZN(new_n888));
  OAI221_X1 g0688(.A(new_n333), .B1(new_n717), .B2(new_n205), .C1(new_n888), .C2(new_n714), .ZN(new_n889));
  NOR3_X1   g0689(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n742), .A2(G311), .B1(new_n755), .B2(G294), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n784), .A2(G283), .B1(G107), .B2(new_n746), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT109), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n890), .B(new_n891), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(new_n892), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n895), .A2(KEYINPUT109), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n884), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT47), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n777), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n898), .B2(new_n897), .ZN(new_n900));
  INV_X1    g0700(.A(new_n694), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n706), .A2(new_n240), .ZN(new_n902));
  AOI211_X1 g0702(.A(new_n699), .B(new_n700), .C1(new_n659), .C2(new_n527), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n901), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(KEYINPUT108), .Z(new_n905));
  OR2_X1    g0705(.A1(new_n645), .A2(new_n522), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n906), .A2(new_n531), .A3(new_n526), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n531), .B2(new_n906), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n900), .B(new_n905), .C1(new_n908), .C2(new_n765), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n626), .A2(new_n644), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n653), .B(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(new_n649), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n689), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT106), .ZN(new_n915));
  XNOR2_X1  g0715(.A(KEYINPUT105), .B(KEYINPUT44), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n645), .A2(new_n490), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n503), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n502), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT101), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n919), .A2(new_n920), .A3(new_n644), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT101), .B1(new_n502), .B2(new_n645), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n918), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n656), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n915), .B(new_n916), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  XOR2_X1   g0726(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n927));
  AOI22_X1  g0727(.A1(new_n503), .A2(new_n917), .B1(new_n921), .B2(new_n922), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n927), .B1(new_n928), .B2(new_n656), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n928), .A2(new_n656), .A3(new_n927), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n926), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n916), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n928), .A2(new_n656), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(KEYINPUT106), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n933), .B1(new_n928), .B2(new_n656), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n654), .B1(new_n932), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT107), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT107), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n940), .B(new_n654), .C1(new_n932), .C2(new_n937), .ZN(new_n941));
  INV_X1    g0741(.A(new_n936), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n942), .A2(KEYINPUT106), .A3(new_n934), .ZN(new_n943));
  INV_X1    g0743(.A(new_n654), .ZN(new_n944));
  OR3_X1    g0744(.A1(new_n928), .A2(new_n656), .A3(new_n927), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n929), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n943), .A2(new_n944), .A3(new_n946), .A4(new_n926), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n914), .A2(new_n939), .A3(new_n941), .A4(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n689), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n660), .B(KEYINPUT41), .Z(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n693), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT42), .ZN(new_n953));
  INV_X1    g0753(.A(new_n655), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n953), .B1(new_n924), .B2(new_n954), .ZN(new_n955));
  NOR3_X1   g0755(.A1(new_n928), .A2(KEYINPUT42), .A3(new_n655), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT102), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n924), .A2(new_n607), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n958), .B1(new_n959), .B2(new_n502), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n958), .B(new_n502), .C1(new_n928), .C2(new_n627), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n645), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n957), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n908), .B(KEYINPUT43), .Z(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n908), .A2(KEYINPUT43), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n957), .B(new_n966), .C1(new_n960), .C2(new_n962), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n967), .A2(KEYINPUT103), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(KEYINPUT103), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n965), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n970), .B1(new_n944), .B2(new_n928), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n944), .A2(new_n928), .ZN(new_n972));
  OAI211_X1 g0772(.A(new_n972), .B(new_n965), .C1(new_n968), .C2(new_n969), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n909), .B1(new_n952), .B2(new_n974), .ZN(G387));
  OR3_X1    g0775(.A1(new_n689), .A2(KEYINPUT110), .A3(new_n912), .ZN(new_n976));
  OAI21_X1  g0776(.A(KEYINPUT110), .B1(new_n689), .B2(new_n912), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n976), .A2(new_n660), .A3(new_n913), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n874), .A2(new_n527), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n784), .A2(G68), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n755), .A2(new_n351), .ZN(new_n981));
  AOI22_X1  g0781(.A1(G150), .A2(new_n750), .B1(new_n722), .B2(G77), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n333), .B1(new_n879), .B2(G97), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n982), .B(new_n983), .C1(new_n727), .C2(new_n202), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(G159), .B2(new_n742), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n979), .A2(new_n980), .A3(new_n981), .A4(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n279), .B1(new_n750), .B2(G326), .ZN(new_n987));
  INV_X1    g0787(.A(G294), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n758), .A2(new_n718), .B1(new_n988), .B2(new_n721), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n736), .A2(new_n735), .B1(new_n727), .B2(new_n888), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n734), .A2(new_n588), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n990), .B(new_n991), .C1(G322), .C2(new_n742), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n989), .B1(new_n992), .B2(KEYINPUT48), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(KEYINPUT48), .B2(new_n992), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT49), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n987), .B1(new_n509), .B2(new_n717), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  AND2_X1   g0796(.A1(new_n994), .A2(new_n995), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n986), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n700), .ZN(new_n999));
  INV_X1    g0799(.A(new_n662), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n703), .A2(new_n1000), .B1(new_n206), .B2(new_n659), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n237), .A2(new_n707), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n351), .A2(new_n202), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT50), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n662), .B(new_n289), .C1(new_n217), .C2(new_n267), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n706), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1001), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n901), .B1(new_n1007), .B2(new_n702), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n999), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(new_n653), .B2(new_n699), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n693), .B2(new_n912), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n978), .A2(new_n1011), .ZN(G393));
  OAI21_X1  g0812(.A(new_n701), .B1(new_n205), .B2(new_n213), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n245), .B2(new_n706), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1014), .A2(new_n901), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT111), .Z(new_n1016));
  AOI22_X1  g0816(.A1(new_n742), .A2(G317), .B1(G311), .B2(new_n753), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT52), .Z(new_n1018));
  AOI22_X1  g0818(.A1(G322), .A2(new_n750), .B1(new_n722), .B2(G283), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n279), .B1(new_n879), .B2(G107), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1019), .B(new_n1020), .C1(new_n736), .C2(new_n588), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(G116), .B2(new_n746), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1018), .B(new_n1022), .C1(new_n988), .C2(new_n734), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n742), .A2(G150), .B1(G159), .B2(new_n753), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT51), .Z(new_n1025));
  NAND2_X1  g0825(.A1(new_n874), .A2(G77), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G143), .A2(new_n750), .B1(new_n722), .B2(G68), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n333), .B1(new_n879), .B2(G87), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(new_n736), .C2(new_n202), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n784), .B2(new_n351), .ZN(new_n1030));
  NAND3_X1  g0830(.A1(new_n1025), .A2(new_n1026), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(KEYINPUT112), .B1(new_n1023), .B2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1032), .A2(new_n777), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1023), .A2(KEYINPUT112), .A3(new_n1031), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1016), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n924), .B2(new_n765), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n938), .A2(new_n947), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1036), .B1(new_n1037), .B2(new_n692), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n661), .B1(new_n1037), .B2(new_n913), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1038), .B1(new_n948), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(G390));
  OAI21_X1  g0841(.A(new_n694), .B1(new_n351), .B2(new_n778), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n742), .A2(G128), .B1(G132), .B2(new_n753), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n1043), .B(KEYINPUT116), .Z(new_n1044));
  NOR2_X1   g0844(.A1(new_n721), .A2(new_n881), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT53), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n333), .B1(new_n750), .B2(G125), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1046), .B(new_n1047), .C1(new_n202), .C2(new_n717), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n874), .B2(G159), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(KEYINPUT54), .B(G143), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT114), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n784), .A2(new_n1051), .B1(G137), .B2(new_n755), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(KEYINPUT115), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1052), .A2(KEYINPUT115), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1044), .A2(new_n1049), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n734), .A2(new_n205), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(G294), .A2(new_n750), .B1(new_n879), .B2(G68), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n279), .B1(new_n722), .B2(G87), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1057), .B(new_n1058), .C1(new_n509), .C2(new_n727), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G283), .B2(new_n742), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1026), .B(new_n1060), .C1(new_n206), .C2(new_n736), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1055), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1042), .B1(new_n1062), .B2(new_n700), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n838), .A2(new_n845), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1063), .B1(new_n1064), .B2(new_n698), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n849), .A2(new_n854), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n836), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1066), .A2(new_n840), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n854), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n847), .B2(new_n848), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n838), .B(new_n845), .C1(new_n1070), .C2(new_n841), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n680), .A2(new_n854), .A3(G330), .A4(new_n772), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT113), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1073), .B(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1072), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1073), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1068), .A2(new_n1071), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1065), .B1(new_n1079), .B2(new_n692), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n438), .A2(new_n682), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n623), .A2(new_n813), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n680), .A2(G330), .A3(new_n772), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n1069), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n1084), .A2(new_n848), .A3(new_n847), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1073), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n1085), .A2(new_n1075), .B1(new_n849), .B2(new_n1086), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1082), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n661), .B1(new_n1079), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1082), .A2(new_n1087), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1090), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1080), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(G378));
  INV_X1    g0893(.A(KEYINPUT57), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n862), .A2(new_n836), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n1095), .A2(KEYINPUT40), .B1(new_n862), .B2(new_n861), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n618), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n433), .B1(new_n1097), .B2(new_n616), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n641), .A2(new_n404), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n619), .A2(new_n433), .A3(new_n1099), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1103), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n1096), .A2(new_n1107), .A3(new_n859), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1103), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n1104), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(new_n867), .B2(G330), .ZN(new_n1113));
  OAI21_X1  g0913(.A(KEYINPUT118), .B1(new_n1108), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n857), .A2(KEYINPUT119), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT119), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n846), .A2(new_n855), .A3(new_n1116), .A4(new_n856), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1107), .B1(new_n1096), .B2(new_n859), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n863), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n866), .B1(new_n862), .B2(new_n836), .ZN(new_n1122));
  OAI211_X1 g0922(.A(G330), .B(new_n1112), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1124), .A2(KEYINPUT118), .A3(new_n1115), .A4(new_n1117), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1119), .A2(new_n1125), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n1068), .A2(new_n1071), .A3(new_n1077), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1075), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n1068), .B2(new_n1071), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1082), .B1(new_n1130), .B2(new_n1090), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1094), .B1(new_n1126), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT120), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g0934(.A(KEYINPUT120), .B(new_n1094), .C1(new_n1126), .C2(new_n1131), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n846), .A2(new_n855), .A3(new_n856), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1120), .A2(new_n1136), .A3(new_n1123), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1136), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1138));
  OAI21_X1  g0938(.A(KEYINPUT57), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n660), .B1(new_n1131), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1134), .A2(new_n1135), .A3(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1107), .A2(new_n697), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n694), .B1(G50), .B2(new_n778), .ZN(new_n1144));
  AOI21_X1  g0944(.A(G50), .B1(new_n278), .B2(new_n291), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n291), .B(new_n333), .C1(new_n721), .C2(new_n267), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n714), .A2(new_n718), .B1(new_n717), .B2(new_n216), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1146), .B(new_n1147), .C1(new_n753), .C2(G107), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n205), .B2(new_n736), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G116), .B2(new_n742), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n875), .B(new_n1150), .C1(new_n422), .C2(new_n734), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT58), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1145), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n753), .A2(G128), .B1(new_n1051), .B2(new_n722), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n792), .B2(new_n736), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1155), .B1(G125), .B2(new_n742), .ZN(new_n1156));
  INV_X1    g0956(.A(G137), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1156), .B1(new_n1157), .B2(new_n734), .C1(new_n881), .C2(new_n761), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1159));
  AOI211_X1 g0959(.A(G33), .B(G41), .C1(new_n750), .C2(G124), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n341), .B2(new_n717), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT117), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1158), .A2(KEYINPUT59), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1153), .B1(new_n1152), .B2(new_n1151), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1144), .B1(new_n1165), .B2(new_n700), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1143), .A2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1167), .B1(new_n1126), .B2(new_n692), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1142), .A2(new_n1169), .ZN(G375));
  OAI21_X1  g0970(.A(new_n694), .B1(G68), .B2(new_n778), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n784), .A2(G107), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n588), .A2(new_n714), .B1(new_n721), .B2(new_n205), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n279), .B1(new_n879), .B2(G77), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n1174), .A2(KEYINPUT121), .B1(new_n727), .B2(new_n718), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1173), .B(new_n1175), .C1(KEYINPUT121), .C2(new_n1174), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n742), .A2(G294), .B1(new_n755), .B2(G116), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n979), .A2(new_n1172), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n755), .A2(new_n1051), .ZN(new_n1179));
  OAI221_X1 g0979(.A(new_n1179), .B1(new_n1157), .B2(new_n727), .C1(new_n782), .C2(new_n792), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT122), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n721), .A2(new_n341), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n279), .B1(new_n717), .B2(new_n216), .ZN(new_n1183));
  AOI211_X1 g0983(.A(new_n1182), .B(new_n1183), .C1(G128), .C2(new_n750), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n734), .B2(new_n881), .C1(new_n761), .C2(new_n202), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1178), .B1(new_n1181), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1171), .B1(new_n1186), .B2(new_n700), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n854), .B2(new_n698), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n1087), .B2(new_n692), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1090), .A2(new_n950), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1082), .A2(new_n1087), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1189), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(G381));
  AOI21_X1  g0993(.A(new_n1140), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1168), .B1(new_n1194), .B2(new_n1135), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n1092), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(G393), .A2(G396), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1197), .A2(new_n802), .A3(new_n1040), .A4(new_n1192), .ZN(new_n1198));
  OR3_X1    g0998(.A1(new_n1196), .A2(G387), .A3(new_n1198), .ZN(G407));
  OAI211_X1 g0999(.A(G407), .B(G213), .C1(G343), .C2(new_n1196), .ZN(G409));
  INV_X1    g1000(.A(new_n1082), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1091), .A2(new_n1201), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1202), .A2(new_n951), .A3(new_n1125), .A4(new_n1119), .ZN(new_n1203));
  OAI21_X1  g1003(.A(KEYINPUT123), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1124), .A2(new_n857), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT123), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1120), .A2(new_n1136), .A3(new_n1123), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1204), .A2(new_n1208), .A3(new_n693), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1092), .A2(new_n1203), .A3(new_n1167), .A4(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n643), .A2(G213), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n1195), .B2(new_n1092), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1082), .A2(new_n1087), .A3(KEYINPUT60), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(new_n660), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1088), .A2(KEYINPUT60), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1215), .B1(new_n1216), .B2(new_n1191), .ZN(new_n1217));
  OR3_X1    g1017(.A1(new_n1217), .A2(new_n802), .A3(new_n1189), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n802), .B1(new_n1217), .B2(new_n1189), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n643), .A2(G213), .A3(G2897), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1220), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT61), .B1(new_n1213), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(G375), .A2(G378), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT62), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1219), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1217), .A2(new_n802), .A3(new_n1189), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1225), .A2(new_n1226), .A3(new_n1229), .A4(new_n1212), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1212), .B(new_n1229), .C1(new_n1195), .C2(new_n1092), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(KEYINPUT62), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1224), .A2(new_n1230), .A3(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(G387), .A2(KEYINPUT124), .A3(new_n1040), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT124), .B1(G387), .B2(new_n1040), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G390), .B(new_n909), .C1(new_n952), .C2(new_n974), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n767), .B1(new_n978), .B2(new_n1011), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1197), .A2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1235), .A2(new_n1236), .A3(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n950), .B1(new_n948), .B2(new_n689), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n971), .B(new_n973), .C1(new_n1242), .C2(new_n693), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT125), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1243), .A2(new_n1244), .A3(new_n909), .A4(G390), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1239), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1244), .B1(G387), .B2(new_n1040), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1247), .B1(new_n1237), .B2(new_n1248), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1241), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1233), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT63), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1231), .A2(new_n1253), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1225), .A2(KEYINPUT63), .A3(new_n1229), .A4(new_n1212), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1224), .A2(new_n1250), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1252), .A2(new_n1256), .ZN(G405));
  AND2_X1   g1057(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(G387), .A2(new_n1040), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1259), .A2(KEYINPUT125), .A3(new_n1237), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT124), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1259), .A2(new_n1262), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(new_n1264), .A3(new_n1234), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT126), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1229), .A2(new_n1266), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1261), .A2(new_n1265), .A3(new_n1267), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1225), .B(new_n1196), .C1(new_n1266), .C2(new_n1229), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1267), .B1(new_n1261), .B2(new_n1265), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1267), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1241), .B2(new_n1249), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1261), .A2(new_n1265), .A3(new_n1267), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1229), .A2(new_n1266), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(new_n1092), .B2(new_n1195), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n1273), .A2(new_n1274), .B1(new_n1225), .B2(new_n1276), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1271), .A2(new_n1277), .ZN(G402));
endmodule


