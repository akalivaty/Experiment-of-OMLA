//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:50 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1246, new_n1247, new_n1248, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n202), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n206), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n209), .B(new_n217), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(new_n219), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT66), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT65), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n234), .B(new_n236), .Z(new_n237));
  INV_X1    g0037(.A(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n232), .B(new_n238), .ZN(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  INV_X1    g0046(.A(G13), .ZN(new_n247));
  NOR3_X1   g0047(.A1(new_n247), .A2(new_n215), .A3(G1), .ZN(new_n248));
  NOR2_X1   g0048(.A1(new_n248), .A2(G50), .ZN(new_n249));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G20), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT69), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n214), .B1(new_n206), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(new_n248), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n249), .B1(new_n257), .B2(G50), .ZN(new_n258));
  INV_X1    g0058(.A(new_n255), .ZN(new_n259));
  XNOR2_X1  g0059(.A(KEYINPUT8), .B(G58), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n215), .A2(G33), .ZN(new_n261));
  OR2_X1    g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n259), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT9), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n266), .B(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(G1698), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n272), .A2(G222), .B1(G77), .B2(new_n271), .ZN(new_n273));
  INV_X1    g0073(.A(G223), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n273), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n214), .ZN(new_n279));
  NAND2_X1  g0079(.A1(G33), .A2(G41), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n250), .A2(G274), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT67), .B(G45), .ZN(new_n285));
  INV_X1    g0085(.A(G41), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G45), .ZN(new_n288));
  AOI21_X1  g0088(.A(G1), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT68), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n280), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(KEYINPUT68), .A2(G33), .A3(G41), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n289), .B1(new_n293), .B2(new_n279), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n287), .B1(new_n294), .B2(G226), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n283), .A2(new_n295), .A3(G190), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n283), .A2(new_n295), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G200), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n268), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT10), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n297), .A2(G169), .ZN(new_n301));
  INV_X1    g0101(.A(G179), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n301), .B1(new_n302), .B2(new_n297), .ZN(new_n303));
  INV_X1    g0103(.A(new_n266), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n260), .A2(G20), .A3(G33), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT15), .B(G87), .ZN(new_n307));
  OAI22_X1  g0107(.A1(new_n307), .A2(new_n261), .B1(new_n215), .B2(new_n220), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n255), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n248), .A2(new_n220), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(new_n257), .B2(new_n220), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n272), .A2(G232), .B1(G107), .B2(new_n271), .ZN(new_n315));
  INV_X1    g0115(.A(G238), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(new_n277), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n282), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n287), .B1(new_n294), .B2(G244), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G200), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G190), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n318), .A2(new_n319), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n314), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n320), .A2(G169), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n318), .A2(new_n319), .A3(G179), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n313), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n300), .A2(new_n305), .A3(new_n329), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n247), .A2(G1), .ZN(new_n331));
  INV_X1    g0131(.A(G68), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(G20), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT12), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT70), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(KEYINPUT12), .B2(new_n333), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n334), .A2(KEYINPUT70), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT11), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n263), .A2(G50), .B1(G20), .B2(new_n332), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(new_n220), .B2(new_n261), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n255), .ZN(new_n341));
  OAI22_X1  g0141(.A1(new_n336), .A2(new_n337), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n338), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(new_n332), .B2(new_n257), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n276), .A2(G232), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G33), .A2(G97), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT3), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n254), .ZN(new_n351));
  NAND2_X1  g0151(.A1(KEYINPUT3), .A2(G33), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n275), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n349), .B1(new_n354), .B2(new_n219), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n282), .B1(new_n348), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT13), .ZN(new_n357));
  INV_X1    g0157(.A(new_n287), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n294), .A2(G238), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n356), .A2(new_n357), .A3(new_n358), .A4(new_n359), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n272), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n281), .B1(new_n361), .B2(new_n347), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n359), .A2(new_n358), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT13), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n360), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT14), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n365), .A2(KEYINPUT71), .A3(new_n366), .A4(G169), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n360), .A2(new_n364), .A3(G179), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(G169), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT71), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n370), .B1(new_n371), .B2(KEYINPUT14), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n365), .A2(new_n372), .B1(KEYINPUT71), .B2(new_n366), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n346), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n365), .A2(new_n321), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n360), .A2(new_n364), .A3(new_n323), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n346), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n374), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n353), .A2(G223), .A3(new_n275), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G33), .A2(G87), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT73), .ZN(new_n382));
  XNOR2_X1  g0182(.A(new_n381), .B(new_n382), .ZN(new_n383));
  OAI211_X1 g0183(.A(G226), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n380), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n282), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n287), .B1(new_n294), .B2(G232), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n388), .A2(G190), .ZN(new_n389));
  AOI21_X1  g0189(.A(G200), .B1(new_n386), .B2(new_n387), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n351), .A2(new_n392), .A3(new_n215), .A4(new_n352), .ZN(new_n393));
  NOR3_X1   g0193(.A1(new_n269), .A2(new_n270), .A3(G20), .ZN(new_n394));
  XNOR2_X1  g0194(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n395));
  OAI211_X1 g0195(.A(G68), .B(new_n393), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  AND2_X1   g0196(.A1(G58), .A2(G68), .ZN(new_n397));
  OAI21_X1  g0197(.A(G20), .B1(new_n397), .B2(new_n201), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n263), .A2(G159), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n351), .A2(new_n215), .A3(new_n352), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n332), .B1(new_n405), .B2(KEYINPUT7), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n271), .A2(new_n395), .A3(new_n215), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n400), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT16), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n404), .A2(new_n409), .A3(new_n255), .ZN(new_n410));
  INV_X1    g0210(.A(new_n260), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n411), .A2(new_n248), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n257), .B2(new_n411), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n410), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n391), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT17), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n386), .A2(new_n302), .A3(new_n387), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n388), .A2(new_n370), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n415), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT18), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT18), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n415), .A2(new_n422), .A3(new_n418), .A4(new_n419), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n410), .B(new_n414), .C1(new_n389), .C2(new_n390), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT17), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n417), .A2(new_n421), .A3(new_n423), .A4(new_n426), .ZN(new_n427));
  NOR3_X1   g0227(.A1(new_n330), .A2(new_n379), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT6), .ZN(new_n429));
  AND2_X1   g0229(.A1(G97), .A2(G107), .ZN(new_n430));
  NOR2_X1   g0230(.A1(G97), .A2(G107), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(G107), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n433), .A2(KEYINPUT6), .A3(G97), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n435), .A2(G20), .B1(G77), .B2(new_n263), .ZN(new_n436));
  OAI211_X1 g0236(.A(G107), .B(new_n393), .C1(new_n394), .C2(new_n395), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n255), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n248), .A2(G97), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n250), .A2(G33), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n441), .B(KEYINPUT74), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n256), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n440), .B1(new_n443), .B2(G97), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT77), .B1(new_n439), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n259), .B1(new_n436), .B2(new_n437), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT77), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n447), .A2(new_n444), .A3(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT4), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(G1698), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n452), .B(G244), .C1(new_n270), .C2(new_n269), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G283), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n221), .B1(new_n351), .B2(new_n352), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n453), .B(new_n454), .C1(new_n455), .C2(KEYINPUT4), .ZN(new_n456));
  OAI21_X1  g0256(.A(G250), .B1(new_n269), .B2(new_n270), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n275), .B1(new_n457), .B2(KEYINPUT4), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n282), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g0259(.A(KEYINPUT5), .B(G41), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n288), .A2(G1), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n460), .A2(G274), .A3(new_n461), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n293), .A2(new_n279), .B1(new_n460), .B2(new_n461), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n462), .B1(new_n463), .B2(G257), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n459), .A2(new_n464), .A3(KEYINPUT76), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT76), .B1(new_n459), .B2(new_n464), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n370), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n459), .A2(new_n464), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G179), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n450), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT76), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n474), .A2(G190), .A3(new_n465), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n447), .A2(new_n444), .ZN(new_n476));
  AOI211_X1 g0276(.A(KEYINPUT75), .B(new_n321), .C1(new_n459), .C2(new_n464), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT75), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n478), .B1(new_n469), .B2(G200), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n475), .B(new_n476), .C1(new_n477), .C2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n215), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT79), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(KEYINPUT79), .A3(new_n215), .ZN(new_n485));
  NOR2_X1   g0285(.A1(G87), .A2(G97), .ZN(new_n486));
  AOI22_X1  g0286(.A1(new_n484), .A2(new_n485), .B1(new_n433), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n215), .B(G68), .C1(new_n269), .C2(new_n270), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n349), .A2(G20), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n488), .B1(KEYINPUT19), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n255), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n307), .A2(new_n248), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n442), .A2(G87), .A3(new_n256), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(G238), .B(new_n275), .C1(new_n269), .C2(new_n270), .ZN(new_n495));
  OAI211_X1 g0295(.A(G244), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G116), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n282), .ZN(new_n499));
  INV_X1    g0299(.A(new_n292), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT68), .B1(G33), .B2(G41), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n279), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G250), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n461), .A2(new_n503), .B1(new_n284), .B2(new_n288), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n499), .A2(G190), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n321), .B1(new_n499), .B2(new_n505), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n494), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT78), .ZN(new_n509));
  AOI221_X4 g0309(.A(G179), .B1(new_n502), .B2(new_n504), .C1(new_n498), .C2(new_n282), .ZN(new_n510));
  AOI21_X1  g0310(.A(G169), .B1(new_n499), .B2(new_n505), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n499), .A2(new_n302), .A3(new_n505), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n498), .A2(new_n282), .B1(new_n502), .B2(new_n504), .ZN(new_n514));
  OAI211_X1 g0314(.A(new_n513), .B(KEYINPUT78), .C1(G169), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n491), .B(new_n492), .C1(new_n307), .C2(new_n443), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n508), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n472), .A2(new_n480), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n254), .A2(G97), .ZN(new_n520));
  AOI21_X1  g0320(.A(G20), .B1(new_n520), .B2(new_n454), .ZN(new_n521));
  INV_X1    g0321(.A(G116), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n215), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n255), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT20), .ZN(new_n525));
  XNOR2_X1  g0325(.A(new_n524), .B(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n248), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n259), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT74), .ZN(new_n529));
  XNOR2_X1  g0329(.A(new_n441), .B(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(G116), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n527), .A2(new_n522), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n370), .B1(new_n526), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n353), .A2(G264), .A3(G1698), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n353), .A2(G257), .A3(new_n275), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n271), .A2(G303), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n282), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n462), .B1(new_n463), .B2(G270), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT80), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT80), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n539), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n534), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT21), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n534), .A2(new_n542), .A3(KEYINPUT21), .A4(new_n544), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n541), .A2(new_n302), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n526), .A2(new_n533), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n547), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n542), .A2(new_n544), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n323), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n542), .A2(new_n321), .A3(new_n544), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n550), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n497), .A2(G20), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT23), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n215), .B2(G107), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n433), .A2(KEYINPUT23), .A3(G20), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n558), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n353), .A2(new_n215), .A3(G87), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT22), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT22), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n353), .A2(new_n566), .A3(new_n215), .A4(G87), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n563), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  OR2_X1    g0368(.A1(new_n568), .A2(KEYINPUT24), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n259), .B1(new_n568), .B2(KEYINPUT24), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n443), .A2(new_n433), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n331), .A2(G20), .A3(new_n433), .ZN(new_n573));
  XNOR2_X1  g0373(.A(new_n573), .B(KEYINPUT25), .ZN(new_n574));
  NOR2_X1   g0374(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(G250), .B(new_n275), .C1(new_n269), .C2(new_n270), .ZN(new_n577));
  OAI211_X1 g0377(.A(G257), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n578));
  XOR2_X1   g0378(.A(KEYINPUT81), .B(G294), .Z(new_n579));
  OAI211_X1 g0379(.A(new_n577), .B(new_n578), .C1(new_n579), .C2(new_n254), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n282), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n463), .A2(G264), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT82), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n462), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n581), .A2(KEYINPUT82), .A3(new_n582), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n321), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n583), .A2(new_n462), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n323), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n576), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n575), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n570), .B2(new_n569), .ZN(new_n594));
  OAI21_X1  g0394(.A(G169), .B1(new_n583), .B2(new_n462), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n585), .A2(G179), .A3(new_n586), .A4(new_n587), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  AND4_X1   g0398(.A1(new_n428), .A2(new_n519), .A3(new_n557), .A4(new_n598), .ZN(G372));
  AND2_X1   g0399(.A1(new_n421), .A2(new_n423), .ZN(new_n600));
  AND2_X1   g0400(.A1(new_n417), .A2(new_n426), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n378), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n365), .A2(new_n372), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n366), .A2(KEYINPUT71), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(new_n367), .A3(new_n368), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n328), .B1(new_n606), .B2(new_n346), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n600), .B1(new_n602), .B2(new_n607), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n608), .A2(new_n300), .B1(new_n304), .B2(new_n303), .ZN(new_n609));
  INV_X1    g0409(.A(new_n428), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n474), .A2(new_n465), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n470), .B1(new_n611), .B2(new_n370), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n518), .A2(new_n612), .A3(KEYINPUT26), .A4(new_n450), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT85), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n450), .A2(new_n468), .A3(new_n471), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n616), .A2(KEYINPUT85), .A3(KEYINPUT26), .A4(new_n518), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT26), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n505), .A2(KEYINPUT83), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT83), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n620), .B1(new_n502), .B2(new_n504), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n499), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n506), .B1(new_n622), .B2(G200), .ZN(new_n623));
  INV_X1    g0423(.A(new_n494), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n510), .B1(new_n622), .B2(new_n370), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n517), .ZN(new_n627));
  INV_X1    g0427(.A(new_n476), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n625), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n468), .A2(new_n471), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n618), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n615), .A2(new_n617), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n596), .A2(new_n595), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n576), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT84), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT84), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n633), .A2(new_n636), .A3(new_n576), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n552), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n581), .A2(KEYINPUT82), .A3(new_n582), .ZN(new_n639));
  AOI21_X1  g0439(.A(KEYINPUT82), .B1(new_n581), .B2(new_n582), .ZN(new_n640));
  NOR3_X1   g0440(.A1(new_n639), .A2(new_n640), .A3(new_n462), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n591), .B1(new_n641), .B2(G200), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n594), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n625), .A2(new_n627), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n643), .A2(new_n644), .A3(new_n480), .A4(new_n472), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n627), .B1(new_n638), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n632), .A2(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n609), .B1(new_n610), .B2(new_n647), .ZN(G369));
  AND3_X1   g0448(.A1(new_n547), .A2(new_n548), .A3(new_n551), .ZN(new_n649));
  INV_X1    g0449(.A(new_n331), .ZN(new_n650));
  OR3_X1    g0450(.A1(new_n650), .A2(KEYINPUT27), .A3(G20), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT27), .B1(new_n650), .B2(G20), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(G213), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(G343), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n550), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n649), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n657), .B1(new_n557), .B2(new_n656), .ZN(new_n658));
  XNOR2_X1  g0458(.A(new_n658), .B(KEYINPUT86), .ZN(new_n659));
  INV_X1    g0459(.A(new_n655), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n643), .B(new_n634), .C1(new_n594), .C2(new_n660), .ZN(new_n661));
  XOR2_X1   g0461(.A(new_n661), .B(KEYINPUT87), .Z(new_n662));
  NAND2_X1  g0462(.A1(new_n597), .A2(new_n655), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n659), .A2(G330), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n635), .A2(new_n637), .A3(new_n660), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n552), .A2(new_n660), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n665), .A2(new_n666), .A3(new_n668), .ZN(G399));
  INV_X1    g0469(.A(new_n207), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(G41), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G1), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n486), .A2(new_n433), .A3(new_n522), .ZN(new_n674));
  INV_X1    g0474(.A(new_n213), .ZN(new_n675));
  OAI22_X1  g0475(.A1(new_n673), .A2(new_n674), .B1(new_n675), .B2(new_n672), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n676), .B(KEYINPUT28), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT29), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n678), .B1(new_n647), .B2(new_n655), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n472), .A2(new_n480), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n625), .A2(new_n627), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n592), .A2(new_n681), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n680), .B(new_n682), .C1(new_n552), .C2(new_n597), .ZN(new_n683));
  OAI21_X1  g0483(.A(KEYINPUT26), .B1(new_n629), .B2(new_n630), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n518), .A2(new_n612), .A3(new_n618), .A4(new_n450), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n684), .A2(new_n685), .A3(new_n627), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n687), .A2(KEYINPUT29), .A3(new_n660), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n679), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n519), .A2(new_n557), .A3(new_n598), .A4(new_n660), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT30), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n585), .A2(KEYINPUT88), .A3(new_n514), .A4(new_n587), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n692), .A2(new_n474), .A3(new_n465), .A4(new_n549), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n585), .A2(new_n514), .A3(new_n587), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT88), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n691), .B1(new_n693), .B2(new_n696), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n474), .A2(new_n549), .A3(new_n465), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n694), .A2(new_n695), .ZN(new_n699));
  NAND4_X1  g0499(.A1(new_n698), .A2(KEYINPUT30), .A3(new_n699), .A4(new_n692), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n469), .A2(new_n302), .A3(new_n622), .ZN(new_n701));
  OR3_X1    g0501(.A1(new_n641), .A2(new_n553), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n697), .A2(new_n700), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(KEYINPUT31), .A3(new_n655), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n690), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(KEYINPUT31), .B1(new_n703), .B2(new_n655), .ZN(new_n706));
  OAI21_X1  g0506(.A(G330), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n689), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g0508(.A(new_n708), .B(KEYINPUT89), .Z(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n677), .B1(new_n710), .B2(G1), .ZN(G364));
  NOR2_X1   g0511(.A1(new_n247), .A2(G20), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n673), .B1(G45), .B2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n670), .A2(new_n353), .ZN(new_n715));
  INV_X1    g0515(.A(new_n285), .ZN(new_n716));
  OAI221_X1 g0516(.A(new_n715), .B1(new_n675), .B2(new_n716), .C1(new_n242), .C2(new_n288), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n670), .A2(new_n271), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n718), .A2(G355), .B1(new_n522), .B2(new_n670), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n279), .B1(new_n215), .B2(G169), .ZN(new_n721));
  OR2_X1    g0521(.A1(new_n721), .A2(KEYINPUT90), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(KEYINPUT90), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G13), .A2(G33), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n714), .B1(new_n720), .B2(new_n728), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT91), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n321), .A2(G179), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n215), .A2(G190), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G179), .A2(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n734), .A2(G283), .B1(new_n737), .B2(G329), .ZN(new_n738));
  XOR2_X1   g0538(.A(new_n738), .B(KEYINPUT96), .Z(new_n739));
  NAND2_X1  g0539(.A1(G20), .A2(G179), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT92), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n323), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G200), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n739), .B1(G311), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n323), .A2(new_n321), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(G326), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n731), .A2(G20), .A3(G190), .ZN(new_n749));
  INV_X1    g0549(.A(G303), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n735), .A2(G190), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OAI221_X1 g0553(.A(new_n271), .B1(new_n749), .B2(new_n750), .C1(new_n753), .C2(new_n579), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n323), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n741), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n748), .B(new_n754), .C1(G322), .C2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n742), .A2(new_n321), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  XOR2_X1   g0560(.A(KEYINPUT33), .B(G317), .Z(new_n761));
  OAI211_X1 g0561(.A(new_n744), .B(new_n758), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n752), .A2(G97), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(new_n760), .B2(new_n332), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT94), .Z(new_n765));
  INV_X1    g0565(.A(G159), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n736), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g0567(.A(KEYINPUT93), .B(KEYINPUT32), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n767), .B(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n749), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G87), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n271), .B1(new_n734), .B2(G107), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n769), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n743), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n220), .ZN(new_n775));
  INV_X1    g0575(.A(G58), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n202), .A2(new_n746), .B1(new_n756), .B2(new_n776), .ZN(new_n777));
  NOR4_X1   g0577(.A1(new_n765), .A2(new_n773), .A3(new_n775), .A4(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n762), .B1(new_n779), .B2(KEYINPUT95), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT95), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n724), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n727), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n730), .B(new_n783), .C1(new_n659), .C2(new_n784), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT97), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n659), .A2(G330), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n659), .A2(G330), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(new_n714), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n786), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT98), .Z(G396));
  INV_X1    g0591(.A(new_n645), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n636), .B1(new_n633), .B2(new_n576), .ZN(new_n793));
  AND3_X1   g0593(.A1(new_n633), .A2(new_n636), .A3(new_n576), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n649), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n792), .A2(new_n795), .B1(new_n517), .B2(new_n626), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n615), .A2(new_n617), .A3(new_n631), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n655), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n328), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n313), .A2(new_n660), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n799), .B1(new_n325), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n328), .A2(new_n660), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n798), .B(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n707), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n713), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(new_n805), .B2(new_n804), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n724), .A2(new_n725), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n714), .B1(new_n808), .B2(new_n220), .ZN(new_n809));
  INV_X1    g0609(.A(new_n724), .ZN(new_n810));
  XNOR2_X1  g0610(.A(KEYINPUT99), .B(G283), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n522), .A2(new_n774), .B1(new_n760), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(G294), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n813), .A2(new_n756), .B1(new_n746), .B2(new_n750), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n353), .B1(new_n737), .B2(G311), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n770), .A2(G107), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n734), .A2(G87), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n815), .A2(new_n816), .A3(new_n763), .A4(new_n817), .ZN(new_n818));
  NOR3_X1   g0618(.A1(new_n812), .A2(new_n814), .A3(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n746), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G137), .A2(new_n820), .B1(new_n757), .B2(G143), .ZN(new_n821));
  INV_X1    g0621(.A(G150), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n821), .B1(new_n760), .B2(new_n822), .C1(new_n766), .C2(new_n774), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT34), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n353), .B1(new_n749), .B2(new_n202), .ZN(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n733), .A2(new_n332), .B1(new_n736), .B2(new_n826), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n825), .B(new_n827), .C1(G58), .C2(new_n752), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n819), .B1(new_n824), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n803), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n809), .B1(new_n810), .B2(new_n829), .C1(new_n830), .C2(new_n726), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n807), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G384));
  OAI211_X1 g0633(.A(G116), .B(new_n216), .C1(new_n435), .C2(KEYINPUT35), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(KEYINPUT35), .B2(new_n435), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT36), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n213), .B(G77), .C1(new_n776), .C2(new_n332), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n202), .A2(G68), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n250), .B(G13), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT40), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT100), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n842), .B(new_n255), .C1(new_n408), .C2(KEYINPUT16), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n843), .A2(new_n409), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n405), .A2(KEYINPUT7), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n407), .A2(new_n845), .A3(G68), .ZN(new_n846));
  AOI21_X1  g0646(.A(KEYINPUT16), .B1(new_n846), .B2(new_n401), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT100), .B1(new_n847), .B2(new_n259), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n413), .B1(new_n844), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n849), .A2(new_n653), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n427), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT37), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n419), .A2(new_n418), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n424), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n850), .B1(new_n854), .B2(KEYINPUT101), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT101), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n856), .B(new_n424), .C1(new_n849), .C2(new_n853), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n852), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(new_n653), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n415), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n420), .A2(new_n860), .A3(new_n852), .A4(new_n424), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(KEYINPUT38), .B(new_n851), .C1(new_n858), .C2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n848), .A2(new_n409), .A3(new_n843), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n853), .B1(new_n865), .B2(new_n414), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT101), .B1(new_n866), .B2(new_n416), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n865), .A2(new_n414), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n859), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n867), .A2(new_n857), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n862), .B1(new_n870), .B2(KEYINPUT37), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n427), .A2(new_n850), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n864), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n863), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n345), .A2(new_n660), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n374), .A2(new_n378), .A3(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n346), .B(new_n655), .C1(new_n606), .C2(new_n377), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n803), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n690), .B(new_n704), .C1(new_n706), .C2(KEYINPUT104), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n706), .A2(KEYINPUT104), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n841), .B1(new_n875), .B2(new_n883), .ZN(new_n884));
  OR2_X1    g0684(.A1(new_n706), .A2(KEYINPUT104), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n706), .A2(KEYINPUT104), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n885), .A2(new_n690), .A3(new_n704), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n862), .A2(KEYINPUT102), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT102), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n861), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n420), .A2(new_n424), .A3(new_n860), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT37), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n888), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n427), .A2(new_n415), .A3(new_n859), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT38), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n863), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n887), .A2(new_n897), .A3(KEYINPUT40), .A4(new_n880), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n884), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n887), .A2(new_n428), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n899), .B(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(G330), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI211_X1 g0703(.A(new_n660), .B(new_n830), .C1(new_n632), .C2(new_n646), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n802), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n878), .A2(new_n879), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(new_n874), .A3(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n600), .A2(new_n859), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n606), .A2(new_n346), .A3(new_n660), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n861), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT38), .B1(new_n913), .B2(new_n851), .ZN(new_n914));
  NOR3_X1   g0714(.A1(new_n871), .A2(new_n872), .A3(new_n864), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT39), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT39), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n896), .A2(new_n863), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n911), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n910), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n428), .B(new_n688), .C1(new_n798), .C2(KEYINPUT29), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT103), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n679), .A2(KEYINPUT103), .A3(new_n428), .A4(new_n688), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(new_n924), .A3(new_n609), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n920), .B(new_n925), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n903), .A2(new_n926), .B1(new_n250), .B2(new_n712), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n903), .A2(new_n926), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n840), .B1(new_n927), .B2(new_n928), .ZN(G367));
  NAND2_X1  g0729(.A1(new_n494), .A2(new_n655), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT105), .Z(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n627), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n644), .B2(new_n931), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n727), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n238), .A2(new_n715), .ZN(new_n935));
  INV_X1    g0735(.A(new_n307), .ZN(new_n936));
  AOI211_X1 g0736(.A(new_n727), .B(new_n724), .C1(new_n670), .C2(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n714), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n756), .A2(new_n822), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n733), .A2(new_n220), .ZN(new_n940));
  XOR2_X1   g0740(.A(KEYINPUT107), .B(G137), .Z(new_n941));
  AOI21_X1  g0741(.A(new_n940), .B1(new_n737), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n271), .B1(new_n770), .B2(G58), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n942), .B(new_n943), .C1(new_n332), .C2(new_n753), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n939), .B(new_n944), .C1(G143), .C2(new_n820), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n945), .B1(new_n202), .B2(new_n774), .C1(new_n766), .C2(new_n760), .ZN(new_n946));
  INV_X1    g0746(.A(G97), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n733), .A2(new_n947), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n353), .B(new_n948), .C1(G317), .C2(new_n737), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n750), .B2(new_n756), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(G311), .B2(new_n820), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n770), .A2(KEYINPUT46), .A3(G116), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT46), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n749), .B2(new_n522), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n952), .B(new_n954), .C1(new_n433), .C2(new_n753), .ZN(new_n955));
  INV_X1    g0755(.A(new_n579), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n955), .B1(new_n956), .B2(new_n759), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n951), .B(new_n957), .C1(new_n774), .C2(new_n811), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n946), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(KEYINPUT47), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n724), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n959), .A2(KEYINPUT47), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n934), .B(new_n938), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n250), .B1(new_n712), .B2(G45), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n680), .B1(new_n476), .B2(new_n660), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n612), .A2(new_n628), .A3(new_n655), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n668), .A2(new_n666), .A3(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT45), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n668), .A2(new_n666), .ZN(new_n972));
  INV_X1    g0772(.A(new_n968), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(KEYINPUT44), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT44), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n972), .A2(new_n976), .A3(new_n973), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n971), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n665), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n975), .A2(new_n977), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n981), .A2(new_n665), .A3(new_n971), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n664), .B1(new_n659), .B2(G330), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n985), .A2(new_n665), .B1(new_n552), .B2(new_n660), .ZN(new_n986));
  NOR3_X1   g0786(.A1(new_n979), .A2(new_n667), .A3(new_n984), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n710), .B1(new_n983), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n671), .B(new_n990), .Z(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n965), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n968), .A2(new_n597), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n655), .B1(new_n994), .B2(new_n472), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n662), .A2(new_n663), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n996), .A2(new_n667), .A3(new_n973), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT42), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n998), .B2(new_n997), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT43), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n933), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1003), .A2(new_n1001), .A3(new_n933), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n933), .A2(new_n1001), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1000), .A2(new_n1005), .A3(new_n1002), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n665), .B2(new_n973), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n665), .A2(new_n973), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1004), .A2(new_n1009), .A3(new_n1006), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n963), .B1(new_n993), .B2(new_n1011), .ZN(G387));
  NOR2_X1   g0812(.A1(new_n988), .A2(new_n709), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n988), .A2(new_n709), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1014), .A2(new_n671), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n988), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n965), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n715), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n232), .B2(new_n716), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(new_n674), .B2(new_n718), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n411), .A2(new_n202), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT50), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n288), .B1(new_n332), .B2(new_n220), .ZN(new_n1024));
  NOR3_X1   g0824(.A1(new_n1023), .A2(new_n674), .A3(new_n1024), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n1021), .A2(new_n1025), .B1(G107), .B2(new_n207), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n714), .B1(new_n1026), .B2(new_n728), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(G68), .A2(new_n743), .B1(new_n759), .B2(new_n411), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n753), .A2(new_n307), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n749), .A2(new_n220), .B1(new_n736), .B2(new_n822), .ZN(new_n1030));
  NOR4_X1   g0830(.A1(new_n1029), .A2(new_n1030), .A3(new_n271), .A4(new_n948), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G50), .A2(new_n757), .B1(new_n820), .B2(G159), .ZN(new_n1032));
  AND3_X1   g0832(.A1(new_n1028), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n820), .A2(G322), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n759), .A2(G311), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n757), .A2(G317), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n774), .B2(new_n750), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT108), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1034), .B(new_n1035), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1041), .A2(KEYINPUT48), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1041), .A2(KEYINPUT48), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n753), .A2(new_n811), .B1(new_n579), .B2(new_n749), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1045), .A2(KEYINPUT49), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n271), .B1(new_n736), .B2(new_n747), .C1(new_n522), .C2(new_n733), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n1045), .B2(KEYINPUT49), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1033), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1027), .B1(new_n1049), .B2(new_n810), .C1(new_n664), .C2(new_n784), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1016), .A2(new_n1018), .A3(new_n1050), .ZN(G393));
  AND2_X1   g0851(.A1(new_n980), .A2(new_n982), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n672), .B1(new_n1052), .B2(new_n1013), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT109), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n982), .A2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n981), .A2(KEYINPUT109), .A3(new_n665), .A4(new_n971), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1055), .A2(new_n980), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n1014), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1053), .A2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1055), .A2(new_n980), .A3(new_n1056), .A4(new_n965), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n728), .B1(new_n947), .B2(new_n207), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n245), .A2(new_n1019), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n713), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(G311), .A2(new_n757), .B1(new_n820), .B2(G317), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT52), .Z(new_n1065));
  AOI21_X1  g0865(.A(new_n353), .B1(new_n734), .B2(G107), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n737), .A2(G322), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1066), .B(new_n1067), .C1(new_n749), .C2(new_n811), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT112), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n760), .A2(new_n750), .B1(new_n522), .B2(new_n753), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(G294), .B2(new_n743), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1065), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n822), .A2(new_n746), .B1(new_n756), .B2(new_n766), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT110), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT51), .Z(new_n1075));
  AOI22_X1  g0875(.A1(new_n770), .A2(G68), .B1(new_n737), .B2(G143), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1076), .A2(new_n353), .A3(new_n817), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT111), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n759), .A2(G50), .B1(G77), .B2(new_n752), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(new_n260), .C2(new_n774), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1072), .B1(new_n1075), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1063), .B1(new_n1081), .B2(new_n724), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n968), .B2(new_n784), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1059), .A2(new_n1060), .A3(new_n1083), .ZN(G390));
  NOR2_X1   g0884(.A1(new_n803), .A2(new_n902), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n906), .B(new_n1085), .C1(new_n881), .C2(new_n882), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n906), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1087), .B1(new_n904), .B2(new_n802), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n911), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n916), .B(new_n918), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n655), .B1(new_n683), .B2(new_n686), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1091), .A2(new_n801), .B1(new_n328), .B2(new_n660), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n897), .B(new_n911), .C1(new_n1092), .C2(new_n1087), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1086), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n880), .B(G330), .C1(new_n705), .C2(new_n706), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1090), .A2(new_n1093), .A3(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  OAI211_X1 g0898(.A(G330), .B(new_n830), .C1(new_n705), .C2(new_n706), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n1087), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n1086), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1092), .A2(new_n1096), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1085), .B1(new_n881), .B2(new_n882), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n1087), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n905), .A2(new_n1101), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n887), .A2(G330), .A3(new_n428), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n923), .A2(new_n924), .A3(new_n1106), .A4(new_n609), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1098), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1108), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1110), .A2(new_n671), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1095), .A2(new_n965), .A3(new_n1097), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n916), .A2(new_n725), .A3(new_n918), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(G97), .A2(new_n743), .B1(new_n759), .B2(G107), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n734), .A2(G68), .B1(new_n737), .B2(G294), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n1116), .A2(new_n271), .A3(new_n771), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n752), .A2(G77), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(G116), .A2(new_n757), .B1(new_n820), .B2(G283), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1115), .A2(new_n1117), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT114), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n353), .B1(new_n733), .B2(new_n202), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G125), .B2(new_n737), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT113), .Z(new_n1124));
  NAND2_X1  g0924(.A1(new_n770), .A2(G150), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT53), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(G132), .B2(new_n757), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n820), .A2(G128), .B1(G159), .B2(new_n752), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT54), .B(G143), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n759), .A2(new_n941), .B1(new_n743), .B2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g0931(.A1(new_n1124), .A2(new_n1127), .A3(new_n1128), .A4(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n810), .B1(new_n1121), .B2(new_n1132), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n714), .B(new_n1133), .C1(new_n260), .C2(new_n808), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1114), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1113), .A2(new_n1135), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1136), .A2(KEYINPUT115), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(KEYINPUT115), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1112), .B1(new_n1137), .B2(new_n1138), .ZN(G378));
  INV_X1    g0939(.A(KEYINPUT57), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT119), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1107), .B(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1140), .B1(new_n1111), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n884), .A2(G330), .A3(new_n898), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n908), .B1(new_n1088), .B2(new_n874), .ZN(new_n1146));
  NOR3_X1   g0946(.A1(new_n915), .A2(new_n895), .A3(KEYINPUT39), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n917), .B1(new_n863), .B2(new_n873), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1089), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n300), .A2(new_n305), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n266), .A2(new_n653), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1153));
  XOR2_X1   g0953(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1152), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1155), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n1146), .A2(new_n1149), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1158), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1145), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1158), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n910), .B2(new_n919), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1146), .A2(new_n1149), .A3(new_n1158), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1163), .A2(new_n1144), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n672), .B1(new_n1143), .B2(new_n1166), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1163), .A2(new_n1144), .A3(new_n1164), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1144), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1169));
  OAI21_X1  g0969(.A(KEYINPUT117), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT117), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1161), .A2(new_n1171), .A3(new_n1165), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1170), .A2(new_n1172), .B1(new_n1111), .B2(new_n1142), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1167), .B1(new_n1173), .B2(KEYINPUT57), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n964), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1158), .A2(new_n725), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n808), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n713), .B1(new_n1177), .B2(G50), .ZN(new_n1178));
  INV_X1    g0978(.A(G283), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n286), .B(new_n271), .C1(new_n736), .C2(new_n1179), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n749), .A2(new_n220), .B1(new_n733), .B2(new_n776), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(G68), .C2(new_n752), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(G97), .A2(new_n759), .B1(new_n743), .B2(new_n936), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G107), .A2(new_n757), .B1(new_n820), .B2(G116), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n271), .A2(new_n286), .ZN(new_n1187));
  AOI21_X1  g0987(.A(G50), .B1(new_n254), .B2(new_n286), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1186), .A2(KEYINPUT58), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G132), .A2(new_n759), .B1(new_n743), .B2(G137), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n753), .A2(new_n822), .B1(new_n1129), .B2(new_n749), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G125), .B2(new_n820), .ZN(new_n1192));
  INV_X1    g0992(.A(G128), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1190), .B(new_n1192), .C1(new_n1193), .C2(new_n756), .ZN(new_n1194));
  XOR2_X1   g0994(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n254), .B(new_n286), .C1(new_n733), .C2(new_n766), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G124), .B2(new_n737), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1189), .B1(KEYINPUT58), .B2(new_n1186), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1178), .B1(new_n1201), .B2(new_n724), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1176), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(KEYINPUT118), .B1(new_n1175), .B2(new_n1204), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1174), .A2(new_n1205), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1161), .A2(new_n1171), .A3(new_n1165), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1171), .B1(new_n1161), .B2(new_n1165), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n965), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT118), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1209), .A2(new_n1210), .A3(new_n1203), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1206), .A2(new_n1211), .ZN(G375));
  NAND2_X1  g1012(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT121), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1213), .B(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n991), .B(KEYINPUT120), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n1108), .A2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1105), .A2(new_n964), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1087), .A2(new_n725), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n713), .B1(new_n1177), .B2(G68), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G107), .A2(new_n743), .B1(new_n759), .B2(G116), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n749), .A2(new_n947), .B1(new_n736), .B2(new_n750), .ZN(new_n1223));
  NOR4_X1   g1023(.A1(new_n1029), .A2(new_n1223), .A3(new_n353), .A4(new_n940), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(G283), .A2(new_n757), .B1(new_n820), .B2(G294), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1222), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n743), .A2(G150), .B1(G50), .B2(new_n752), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT122), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n749), .A2(new_n766), .B1(new_n736), .B2(new_n1193), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n271), .B(new_n1229), .C1(G58), .C2(new_n734), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n759), .A2(new_n1130), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n757), .A2(new_n941), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n820), .A2(G132), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1226), .B1(new_n1228), .B2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1221), .B1(new_n1235), .B2(new_n724), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1236), .B(KEYINPUT123), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1219), .B1(new_n1220), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1218), .A2(new_n1238), .ZN(G381));
  NOR2_X1   g1039(.A1(G387), .A2(G390), .ZN(new_n1240));
  NOR4_X1   g1040(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1112), .A2(new_n1113), .A3(new_n1135), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1206), .A2(new_n1211), .A3(new_n1243), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1242), .A2(new_n1244), .ZN(G407));
  NAND2_X1  g1045(.A1(new_n654), .A2(G213), .ZN(new_n1246));
  OR2_X1    g1046(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(G407), .A2(G213), .A3(new_n1247), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT124), .ZN(G409));
  NAND4_X1  g1049(.A1(new_n1174), .A2(new_n1205), .A3(G378), .A4(new_n1211), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1204), .B1(new_n1166), .B2(new_n965), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1111), .A2(new_n1142), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1251), .B1(new_n1253), .B2(new_n1216), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n1243), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1250), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1109), .A2(KEYINPUT60), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1215), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1105), .A2(new_n1107), .A3(KEYINPUT60), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(new_n671), .A3(new_n1259), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1260), .A2(G384), .A3(new_n1238), .ZN(new_n1261));
  AOI21_X1  g1061(.A(G384), .B1(new_n1260), .B2(new_n1238), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1256), .A2(new_n1246), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(KEYINPUT62), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1256), .A2(new_n1246), .ZN(new_n1266));
  INV_X1    g1066(.A(G2897), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n1261), .A2(new_n1262), .B1(new_n1267), .B2(new_n1246), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1260), .A2(new_n1238), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n832), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1260), .A2(G384), .A3(new_n1238), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1246), .A2(new_n1267), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1271), .A3(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1268), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1266), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT61), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT62), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1256), .A2(new_n1277), .A3(new_n1246), .A4(new_n1263), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1265), .A2(new_n1275), .A3(new_n1276), .A4(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(KEYINPUT126), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT61), .B1(new_n1266), .B2(new_n1274), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT126), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1281), .A2(new_n1265), .A3(new_n1282), .A4(new_n1278), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G387), .A2(G390), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1013), .A2(new_n982), .A3(new_n980), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n991), .B1(new_n1285), .B2(new_n710), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1010), .B(new_n1008), .C1(new_n1286), .C2(new_n965), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1060), .A2(new_n1083), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1287), .A2(new_n963), .A3(new_n1059), .A4(new_n1288), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(G393), .B(G396), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1284), .A2(new_n1289), .A3(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1290), .B1(new_n1284), .B2(new_n1289), .ZN(new_n1292));
  OAI21_X1  g1092(.A(KEYINPUT127), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1284), .A2(new_n1289), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1290), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT127), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1284), .A2(new_n1289), .A3(new_n1290), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1296), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1293), .A2(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1280), .A2(new_n1283), .A3(new_n1300), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1264), .ZN(new_n1302));
  OR2_X1    g1102(.A1(new_n1302), .A2(KEYINPUT63), .ZN(new_n1303));
  NOR3_X1   g1103(.A1(new_n1291), .A2(new_n1292), .A3(KEYINPUT61), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1302), .A2(KEYINPUT63), .ZN(new_n1305));
  AND3_X1   g1105(.A1(new_n1268), .A2(KEYINPUT125), .A3(new_n1273), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT125), .B1(new_n1268), .B2(new_n1273), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1266), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1303), .A2(new_n1304), .A3(new_n1305), .A4(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1301), .A2(new_n1309), .ZN(G405));
  INV_X1    g1110(.A(new_n1263), .ZN(new_n1311));
  NOR3_X1   g1111(.A1(new_n1291), .A2(new_n1292), .A3(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1263), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(G375), .A2(new_n1243), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1250), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(new_n1316), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n1250), .B(new_n1315), .C1(new_n1312), .C2(new_n1313), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(G402));
endmodule


