//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 0 0 0 1 0 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1139,
    new_n1140, new_n1141, new_n1142, new_n1143, new_n1144, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1162, new_n1163, new_n1164, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n206));
  INV_X1    g0006(.A(G116), .ZN(new_n207));
  INV_X1    g0007(.A(G270), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(G226), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n210), .B1(new_n202), .B2(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n209), .B(new_n214), .C1(G97), .C2(G257), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G1), .B2(G20), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT1), .Z(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR3_X1   g0020(.A1(new_n218), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G1), .ZN(new_n222));
  NOR3_X1   g0022(.A1(new_n222), .A2(new_n219), .A3(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT0), .Z(new_n225));
  NOR3_X1   g0025(.A1(new_n217), .A2(new_n221), .A3(new_n225), .ZN(G361));
  XNOR2_X1  g0026(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G226), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G250), .B(G257), .Z(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G87), .B(G97), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT65), .ZN(new_n237));
  XOR2_X1   g0037(.A(G107), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(new_n220), .ZN(new_n244));
  NAND2_X1  g0044(.A1(G33), .A2(G41), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g0046(.A(new_n222), .B1(G41), .B2(G45), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT70), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT70), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n250), .A2(G238), .A3(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G274), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n247), .A2(new_n254), .ZN(new_n255));
  XOR2_X1   g0055(.A(new_n255), .B(KEYINPUT69), .Z(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G97), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  OR2_X1    g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  AOI21_X1  g0060(.A(G1698), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AND2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  OAI211_X1 g0063(.A(G232), .B(G1698), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT68), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n259), .A2(new_n260), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT68), .ZN(new_n267));
  NAND4_X1  g0067(.A1(new_n266), .A2(new_n267), .A3(G232), .A4(G1698), .ZN(new_n268));
  AOI221_X4 g0068(.A(new_n258), .B1(G226), .B2(new_n261), .C1(new_n265), .C2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n246), .A2(KEYINPUT66), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT66), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n244), .A2(new_n271), .A3(new_n245), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n253), .B(new_n256), .C1(new_n269), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(KEYINPUT13), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT71), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n265), .A2(new_n268), .B1(G226), .B2(new_n261), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n257), .ZN(new_n278));
  AND2_X1   g0078(.A1(new_n270), .A2(new_n272), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT13), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n280), .A2(new_n281), .A3(new_n253), .A4(new_n256), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n275), .A2(new_n276), .A3(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n250), .A2(new_n252), .ZN(new_n284));
  AOI22_X1  g0084(.A1(G238), .A2(new_n284), .B1(new_n278), .B2(new_n279), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n285), .A2(KEYINPUT71), .A3(new_n281), .A4(new_n256), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n283), .A2(G169), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT73), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(KEYINPUT14), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n275), .A2(new_n282), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n292), .A2(G179), .B1(new_n288), .B2(KEYINPUT14), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n283), .A2(G169), .A3(new_n289), .A4(new_n286), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n220), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G20), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n219), .A2(G33), .ZN(new_n300));
  INV_X1    g0100(.A(G77), .ZN(new_n301));
  OAI22_X1  g0101(.A1(new_n299), .A2(new_n202), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n219), .A2(G68), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n297), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n304), .B(KEYINPUT11), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n297), .B1(new_n222), .B2(G20), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G68), .ZN(new_n307));
  INV_X1    g0107(.A(G13), .ZN(new_n308));
  NOR3_X1   g0108(.A1(new_n308), .A2(new_n219), .A3(G1), .ZN(new_n309));
  AOI21_X1  g0109(.A(KEYINPUT72), .B1(new_n309), .B2(new_n212), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT12), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n305), .A2(new_n307), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n295), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n292), .A2(G190), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n283), .A2(G200), .A3(new_n286), .ZN(new_n315));
  INV_X1    g0115(.A(new_n312), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G20), .A2(G77), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT15), .B(G87), .ZN(new_n319));
  XNOR2_X1  g0119(.A(KEYINPUT8), .B(G58), .ZN(new_n320));
  OAI221_X1 g0120(.A(new_n318), .B1(new_n319), .B2(new_n300), .C1(new_n299), .C2(new_n320), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n321), .A2(new_n297), .B1(new_n301), .B2(new_n309), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n306), .A2(G77), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G1698), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G232), .ZN(new_n326));
  OAI221_X1 g0126(.A(new_n326), .B1(new_n213), .B2(new_n325), .C1(new_n262), .C2(new_n263), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n262), .A2(new_n263), .ZN(new_n328));
  INV_X1    g0128(.A(G107), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n327), .A2(new_n270), .A3(new_n330), .A4(new_n272), .ZN(new_n331));
  INV_X1    g0131(.A(new_n255), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n246), .A2(G244), .A3(new_n247), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G169), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n331), .A2(new_n337), .A3(new_n332), .A4(new_n333), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT67), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n338), .A2(new_n339), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n324), .B(new_n336), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n322), .A2(new_n323), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n334), .A2(G200), .ZN(new_n345));
  INV_X1    g0145(.A(G190), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n344), .B(new_n345), .C1(new_n346), .C2(new_n334), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n313), .A2(new_n317), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n325), .A2(G222), .ZN(new_n350));
  INV_X1    g0150(.A(G223), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n266), .B(new_n350), .C1(new_n351), .C2(new_n325), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n279), .B(new_n352), .C1(G77), .C2(new_n266), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n249), .A2(G226), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n353), .A2(new_n332), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n203), .A2(G20), .ZN(new_n357));
  INV_X1    g0157(.A(G150), .ZN(new_n358));
  OAI221_X1 g0158(.A(new_n357), .B1(new_n358), .B2(new_n299), .C1(new_n320), .C2(new_n300), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n359), .A2(new_n297), .B1(new_n202), .B2(new_n309), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n306), .A2(G50), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n356), .A2(G190), .B1(new_n362), .B2(KEYINPUT9), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n355), .A2(G200), .ZN(new_n364));
  OR2_X1    g0164(.A1(new_n362), .A2(KEYINPUT9), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  XOR2_X1   g0166(.A(new_n366), .B(KEYINPUT10), .Z(new_n367));
  NAND2_X1  g0167(.A1(new_n351), .A2(new_n325), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n211), .A2(G1698), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n368), .B(new_n369), .C1(new_n262), .C2(new_n263), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G87), .ZN(new_n371));
  AND3_X1   g0171(.A1(new_n370), .A2(KEYINPUT75), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT75), .B1(new_n370), .B2(new_n371), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n279), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT76), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n279), .B(KEYINPUT76), .C1(new_n372), .C2(new_n373), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n255), .B1(new_n249), .B2(G232), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n380), .A2(G190), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(G200), .B1(new_n374), .B2(new_n379), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n320), .A2(new_n309), .ZN(new_n386));
  INV_X1    g0186(.A(new_n306), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n386), .B1(new_n387), .B2(new_n320), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n259), .A2(new_n219), .A3(new_n260), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT7), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n259), .A2(KEYINPUT7), .A3(new_n219), .A4(new_n260), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n212), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G58), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n394), .A2(new_n212), .ZN(new_n395));
  OAI21_X1  g0195(.A(G20), .B1(new_n395), .B2(new_n201), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n298), .A2(G159), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT16), .B1(new_n393), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT7), .B1(new_n328), .B2(new_n219), .ZN(new_n400));
  NOR4_X1   g0200(.A1(new_n262), .A2(new_n263), .A3(new_n390), .A4(G20), .ZN(new_n401));
  OAI21_X1  g0201(.A(G68), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  INV_X1    g0203(.A(new_n398), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n403), .A2(KEYINPUT74), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n399), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n297), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n393), .A2(new_n398), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n409), .B1(new_n410), .B2(new_n406), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n388), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n385), .A2(KEYINPUT17), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT17), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n408), .A2(new_n411), .ZN(new_n415));
  INV_X1    g0215(.A(new_n388), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n383), .B1(new_n378), .B2(new_n381), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n414), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n413), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(G169), .B1(new_n374), .B2(new_n379), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n380), .A2(G179), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n421), .B1(new_n378), .B2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT18), .B1(new_n417), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT77), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n417), .A2(new_n423), .A3(KEYINPUT18), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI211_X1 g0227(.A(KEYINPUT77), .B(KEYINPUT18), .C1(new_n417), .C2(new_n423), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n420), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n356), .A2(new_n337), .ZN(new_n430));
  INV_X1    g0230(.A(new_n362), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n355), .A2(new_n335), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n367), .A2(new_n429), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n349), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n219), .B(G87), .C1(new_n262), .C2(new_n263), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(KEYINPUT22), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT22), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n266), .A2(new_n440), .A3(new_n219), .A4(G87), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(KEYINPUT82), .B1(new_n219), .B2(G107), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n443), .A2(KEYINPUT23), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(KEYINPUT23), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n219), .A2(G33), .A3(G116), .ZN(new_n447));
  XNOR2_X1  g0247(.A(new_n447), .B(KEYINPUT81), .ZN(new_n448));
  NAND2_X1  g0248(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n442), .A2(new_n446), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(KEYINPUT83), .A2(KEYINPUT24), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n439), .A2(new_n441), .B1(new_n444), .B2(new_n445), .ZN(new_n453));
  INV_X1    g0253(.A(new_n451), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n453), .A2(new_n448), .A3(new_n449), .A4(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n452), .A2(new_n297), .A3(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n309), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G107), .ZN(new_n458));
  OR2_X1    g0258(.A1(new_n458), .A2(KEYINPUT25), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n459), .A2(KEYINPUT84), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT84), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n461), .B1(new_n458), .B2(KEYINPUT25), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n222), .A2(G33), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n457), .A2(new_n409), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n459), .A2(new_n462), .B1(G107), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n456), .A2(new_n460), .A3(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n266), .B1(G257), .B2(new_n325), .ZN(new_n468));
  NOR2_X1   g0268(.A1(G250), .A2(G1698), .ZN(new_n469));
  INV_X1    g0269(.A(G33), .ZN(new_n470));
  INV_X1    g0270(.A(G294), .ZN(new_n471));
  OAI22_X1  g0271(.A1(new_n468), .A2(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n279), .ZN(new_n473));
  XNOR2_X1  g0273(.A(KEYINPUT5), .B(G41), .ZN(new_n474));
  INV_X1    g0274(.A(G45), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(G1), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n477), .A2(new_n246), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G264), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n474), .A2(G274), .A3(new_n476), .ZN(new_n481));
  XNOR2_X1  g0281(.A(new_n481), .B(KEYINPUT78), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n335), .B1(new_n480), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n480), .A2(new_n483), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n337), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n467), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n325), .A2(G257), .ZN(new_n488));
  NAND2_X1  g0288(.A1(G264), .A2(G1698), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n266), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G303), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n328), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n490), .A2(new_n492), .A3(new_n270), .A4(new_n272), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n477), .A2(G270), .A3(new_n246), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n481), .A2(KEYINPUT78), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n481), .A2(KEYINPUT78), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n493), .B(new_n494), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G200), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n457), .A2(G116), .A3(new_n409), .A4(new_n463), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n309), .A2(new_n207), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n296), .A2(new_n220), .B1(G20), .B2(new_n207), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G283), .ZN(new_n502));
  INV_X1    g0302(.A(G97), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n502), .B(new_n219), .C1(G33), .C2(new_n503), .ZN(new_n504));
  AND3_X1   g0304(.A1(new_n501), .A2(KEYINPUT20), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(KEYINPUT20), .B1(new_n501), .B2(new_n504), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n499), .B(new_n500), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n498), .B(new_n508), .C1(new_n346), .C2(new_n497), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT21), .ZN(new_n510));
  INV_X1    g0310(.A(new_n497), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n507), .A2(G169), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(G179), .A3(new_n507), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n497), .A2(new_n507), .A3(KEYINPUT21), .A4(G169), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n509), .A2(new_n513), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  XNOR2_X1  g0316(.A(new_n516), .B(KEYINPUT80), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n266), .A2(KEYINPUT4), .A3(G244), .A4(new_n325), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT4), .ZN(new_n519));
  INV_X1    g0319(.A(G244), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n519), .B1(new_n328), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n518), .A2(new_n521), .A3(new_n502), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n266), .A2(G250), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n325), .B1(new_n523), .B2(KEYINPUT4), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n279), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n478), .A2(G257), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(new_n482), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G200), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n457), .A2(G97), .ZN(new_n529));
  OAI21_X1  g0329(.A(G107), .B1(new_n400), .B2(new_n401), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT6), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n503), .A2(new_n329), .ZN(new_n532));
  NOR2_X1   g0332(.A1(G97), .A2(G107), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n329), .A2(KEYINPUT6), .A3(G97), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G20), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n298), .A2(G77), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n530), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n529), .B1(new_n539), .B2(new_n297), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n465), .A2(G97), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n525), .A2(G190), .A3(new_n482), .A4(new_n526), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n528), .A2(new_n540), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n527), .A2(new_n335), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n539), .A2(new_n297), .ZN(new_n545));
  INV_X1    g0345(.A(new_n529), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(new_n541), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n525), .A2(new_n337), .A3(new_n482), .A4(new_n526), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n544), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT19), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n219), .B1(new_n257), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(G87), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n553), .A2(new_n503), .A3(new_n329), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT79), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n266), .A2(new_n219), .A3(G68), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n552), .A2(KEYINPUT79), .A3(new_n554), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n551), .B1(new_n300), .B2(new_n503), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n557), .A2(new_n558), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n297), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n319), .A2(new_n309), .ZN(new_n563));
  OR2_X1    g0363(.A1(new_n464), .A2(new_n319), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n476), .A2(G274), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n246), .B(G250), .C1(G1), .C2(new_n475), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n259), .A2(new_n260), .B1(new_n520), .B2(G1698), .ZN(new_n568));
  NOR2_X1   g0368(.A1(G238), .A2(G1698), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n568), .A2(new_n570), .B1(G33), .B2(G116), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n566), .B(new_n567), .C1(new_n571), .C2(new_n273), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n335), .ZN(new_n573));
  OAI22_X1  g0373(.A1(new_n262), .A2(new_n263), .B1(G244), .B2(new_n325), .ZN(new_n574));
  OAI22_X1  g0374(.A1(new_n574), .A2(new_n569), .B1(new_n470), .B2(new_n207), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n279), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n576), .A2(new_n337), .A3(new_n566), .A4(new_n567), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n565), .A2(new_n573), .A3(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n576), .A2(G190), .A3(new_n566), .A4(new_n567), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n572), .A2(G200), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n561), .A2(new_n297), .B1(new_n309), .B2(new_n319), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n465), .A2(G87), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n579), .A2(new_n580), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n456), .A2(new_n460), .A3(new_n466), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n485), .A2(G190), .ZN(new_n586));
  INV_X1    g0386(.A(new_n485), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G200), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n550), .A2(new_n584), .A3(new_n589), .ZN(new_n590));
  AND4_X1   g0390(.A1(new_n437), .A2(new_n487), .A3(new_n517), .A4(new_n590), .ZN(G372));
  NAND3_X1  g0391(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n487), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n594), .A2(new_n550), .A3(new_n584), .A4(new_n589), .ZN(new_n595));
  INV_X1    g0395(.A(new_n578), .ZN(new_n596));
  AND3_X1   g0396(.A1(new_n544), .A2(new_n547), .A3(new_n548), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n597), .A2(new_n584), .A3(KEYINPUT26), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT26), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n578), .A2(new_n583), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n599), .B1(new_n549), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n596), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n595), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n437), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g0404(.A(new_n366), .B(KEYINPUT10), .ZN(new_n605));
  OR2_X1    g0405(.A1(new_n338), .A2(new_n339), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n344), .B1(new_n340), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n607), .A2(KEYINPUT85), .A3(new_n336), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT85), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n343), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(new_n295), .B2(new_n312), .ZN(new_n612));
  INV_X1    g0412(.A(new_n317), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n413), .A2(new_n419), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n417), .A2(new_n423), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT18), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n426), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n605), .B1(new_n615), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n604), .A2(new_n433), .A3(new_n621), .ZN(G369));
  NOR2_X1   g0422(.A1(new_n308), .A2(G20), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n222), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n624), .A2(KEYINPUT27), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(KEYINPUT27), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(G213), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(G343), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n630), .A2(new_n508), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n592), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT80), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n516), .B(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n632), .B1(new_n634), .B2(new_n631), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n635), .B(KEYINPUT86), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n487), .A2(new_n629), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n589), .B1(new_n585), .B2(new_n630), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n637), .B1(new_n638), .B2(new_n487), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n636), .A2(G330), .A3(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n637), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n593), .A2(new_n629), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n487), .ZN(new_n644));
  INV_X1    g0444(.A(new_n589), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OR2_X1    g0446(.A1(new_n641), .A2(new_n646), .ZN(G399));
  INV_X1    g0447(.A(new_n223), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT87), .ZN(new_n649));
  OR3_X1    g0449(.A1(new_n648), .A2(new_n649), .A3(G41), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n649), .B1(new_n648), .B2(G41), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n554), .A2(G116), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n652), .A2(G1), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(new_n218), .B2(new_n652), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT28), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n629), .B1(new_n595), .B2(new_n602), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(KEYINPUT89), .A2(KEYINPUT29), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n659), .ZN(new_n661));
  NAND2_X1  g0461(.A1(KEYINPUT89), .A2(KEYINPUT29), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n661), .B1(new_n657), .B2(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n590), .A2(new_n487), .A3(new_n517), .A4(new_n630), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT88), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n497), .A2(new_n337), .ZN(new_n667));
  INV_X1    g0467(.A(new_n572), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n667), .A2(new_n473), .A3(new_n479), .A4(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n666), .B1(new_n669), .B2(new_n527), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(KEYINPUT30), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n668), .A2(G179), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n587), .A2(new_n672), .A3(new_n497), .A4(new_n527), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT30), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n666), .B(new_n674), .C1(new_n669), .C2(new_n527), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n671), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n629), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT31), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n676), .A2(KEYINPUT31), .A3(new_n629), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n665), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  AOI22_X1  g0481(.A1(new_n660), .A2(new_n664), .B1(new_n681), .B2(G330), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n656), .B1(new_n682), .B2(G1), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n683), .B(KEYINPUT90), .Z(G364));
  AOI21_X1  g0484(.A(new_n222), .B1(new_n623), .B2(G45), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n652), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g0486(.A(new_n686), .B(KEYINPUT91), .Z(new_n687));
  AOI21_X1  g0487(.A(new_n687), .B1(new_n636), .B2(G330), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(G330), .B2(new_n636), .ZN(new_n689));
  XOR2_X1   g0489(.A(new_n687), .B(KEYINPUT92), .Z(new_n690));
  NAND2_X1  g0490(.A1(new_n346), .A2(G20), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n691), .A2(new_n337), .A3(G200), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n266), .B1(new_n692), .B2(G311), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n219), .A2(new_n346), .ZN(new_n694));
  AND2_X1   g0494(.A1(G179), .A2(G200), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(G326), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n693), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n691), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n695), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(G317), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT33), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n703), .A2(KEYINPUT33), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n702), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(G179), .A2(G200), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n700), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(G329), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n694), .A2(new_n337), .A3(G200), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n706), .B(new_n710), .C1(new_n491), .C2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n219), .B1(new_n707), .B2(G190), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AOI211_X1 g0514(.A(new_n699), .B(new_n712), .C1(G294), .C2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n337), .A2(G200), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n694), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(G322), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n700), .A2(new_n337), .A3(G200), .ZN(new_n720));
  OR2_X1    g0520(.A1(new_n720), .A2(KEYINPUT95), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(KEYINPUT95), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT96), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(G283), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n715), .B(new_n719), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n713), .A2(new_n503), .ZN(new_n728));
  INV_X1    g0528(.A(new_n711), .ZN(new_n729));
  AOI22_X1  g0529(.A1(G68), .A2(new_n702), .B1(new_n729), .B2(G87), .ZN(new_n730));
  OAI221_X1 g0530(.A(new_n730), .B1(new_n202), .B2(new_n697), .C1(new_n394), .C2(new_n717), .ZN(new_n731));
  AOI211_X1 g0531(.A(new_n728), .B(new_n731), .C1(G77), .C2(new_n692), .ZN(new_n732));
  XNOR2_X1  g0532(.A(KEYINPUT93), .B(G159), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n709), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g0534(.A(new_n734), .B(KEYINPUT94), .Z(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(KEYINPUT32), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n735), .A2(KEYINPUT32), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n732), .A2(new_n266), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n725), .A2(new_n329), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n727), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n220), .B1(G20), .B2(new_n335), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n690), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n648), .A2(new_n266), .ZN(new_n743));
  OR2_X1    g0543(.A1(new_n218), .A2(G45), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n743), .B(new_n744), .C1(new_n242), .C2(new_n475), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n266), .A2(new_n223), .A3(G355), .ZN(new_n746));
  OAI211_X1 g0546(.A(new_n745), .B(new_n746), .C1(G116), .C2(new_n223), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G13), .A2(G33), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G20), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n741), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n747), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n750), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n742), .B(new_n752), .C1(new_n635), .C2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n689), .A2(new_n754), .ZN(G396));
  NOR2_X1   g0555(.A1(new_n344), .A2(new_n630), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n611), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT98), .ZN(new_n758));
  INV_X1    g0558(.A(new_n756), .ZN(new_n759));
  AND3_X1   g0559(.A1(new_n759), .A2(new_n343), .A3(new_n347), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n757), .A2(new_n758), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n759), .B1(new_n608), .B2(new_n610), .ZN(new_n763));
  OAI21_X1  g0563(.A(KEYINPUT98), .B1(new_n763), .B2(new_n760), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n658), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n603), .A2(new_n762), .A3(new_n630), .A4(new_n764), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n681), .A2(G330), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT99), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n687), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n768), .A2(new_n769), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n772), .B(new_n773), .C1(new_n771), .C2(new_n770), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n724), .A2(G87), .ZN(new_n775));
  AOI22_X1  g0575(.A1(G283), .A2(new_n702), .B1(new_n709), .B2(G311), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(new_n471), .B2(new_n717), .ZN(new_n777));
  INV_X1    g0577(.A(new_n692), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n328), .B1(new_n778), .B2(new_n207), .C1(new_n697), .C2(new_n491), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n777), .A2(new_n728), .A3(new_n779), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n775), .B(new_n780), .C1(new_n329), .C2(new_n711), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n724), .A2(G68), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n266), .B1(new_n713), .B2(new_n394), .C1(new_n711), .C2(new_n202), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n702), .A2(G150), .B1(new_n718), .B2(G143), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n692), .A2(new_n733), .ZN(new_n785));
  INV_X1    g0585(.A(G137), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n784), .B(new_n785), .C1(new_n786), .C2(new_n697), .ZN(new_n787));
  XNOR2_X1  g0587(.A(KEYINPUT97), .B(KEYINPUT34), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n783), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n782), .B(new_n789), .C1(new_n788), .C2(new_n787), .ZN(new_n790));
  INV_X1    g0590(.A(G132), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n708), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n781), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n690), .B1(new_n793), .B2(new_n741), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n741), .A2(new_n748), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n765), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n794), .B1(G77), .B2(new_n796), .C1(new_n797), .C2(new_n749), .ZN(new_n798));
  AND2_X1   g0598(.A1(new_n774), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(G384));
  INV_X1    g0600(.A(KEYINPUT40), .ZN(new_n801));
  INV_X1    g0601(.A(new_n627), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n399), .A2(new_n405), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n416), .B1(new_n803), .B2(new_n409), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n429), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n385), .A2(new_n412), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n417), .A2(new_n802), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n806), .A2(new_n616), .A3(new_n807), .ZN(new_n808));
  OR2_X1    g0608(.A1(new_n808), .A2(KEYINPUT37), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n804), .B1(new_n423), .B2(new_n802), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n806), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(KEYINPUT37), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n809), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AND3_X1   g0613(.A1(new_n805), .A2(KEYINPUT38), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(KEYINPUT38), .B1(new_n805), .B2(new_n813), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n312), .A2(new_n629), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n313), .A2(new_n317), .A3(new_n817), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n312), .B(new_n629), .C1(new_n295), .C2(new_n613), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n820), .A2(new_n681), .A3(new_n797), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n801), .B1(new_n816), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n807), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n619), .B1(new_n614), .B2(KEYINPUT102), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n614), .A2(KEYINPUT102), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n808), .B(KEYINPUT37), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT38), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n805), .A2(KEYINPUT38), .A3(new_n813), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n681), .A2(new_n797), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n832), .A2(KEYINPUT40), .A3(new_n820), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n822), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n437), .A2(new_n681), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n835), .B(new_n836), .Z(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(G330), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n620), .A2(new_n627), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n607), .A2(new_n336), .A3(new_n630), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n767), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n820), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n839), .B1(new_n816), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT101), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT39), .ZN(new_n846));
  AOI21_X1  g0646(.A(KEYINPUT38), .B1(new_n826), .B2(new_n827), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n814), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n426), .A2(new_n425), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n618), .ZN(new_n850));
  INV_X1    g0650(.A(new_n428), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n614), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n804), .ZN(new_n853));
  NOR3_X1   g0653(.A1(new_n852), .A2(new_n627), .A3(new_n853), .ZN(new_n854));
  MUX2_X1   g0654(.A(new_n808), .B(new_n811), .S(KEYINPUT37), .Z(new_n855));
  OAI21_X1  g0655(.A(new_n829), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n856), .A2(KEYINPUT39), .A3(new_n831), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n295), .A2(new_n312), .A3(new_n630), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n848), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(KEYINPUT101), .B(new_n839), .C1(new_n816), .C2(new_n842), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n845), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n349), .A2(new_n660), .A3(new_n664), .A4(new_n435), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n621), .A2(new_n433), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n862), .B(new_n864), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n838), .B(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n222), .B2(new_n623), .ZN(new_n867));
  OAI211_X1 g0667(.A(G20), .B(new_n244), .C1(new_n536), .C2(KEYINPUT35), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n207), .B(new_n868), .C1(KEYINPUT35), .C2(new_n536), .ZN(new_n869));
  XOR2_X1   g0669(.A(new_n869), .B(KEYINPUT36), .Z(new_n870));
  OAI21_X1  g0670(.A(G77), .B1(new_n394), .B2(new_n212), .ZN(new_n871));
  OAI22_X1  g0671(.A1(new_n871), .A2(new_n218), .B1(G50), .B2(new_n212), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(G1), .A3(new_n308), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n873), .B(KEYINPUT100), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n867), .A2(new_n870), .A3(new_n874), .ZN(G367));
  NOR2_X1   g0675(.A1(new_n713), .A2(new_n212), .ZN(new_n876));
  INV_X1    g0676(.A(G143), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n266), .B1(new_n394), .B2(new_n711), .C1(new_n697), .C2(new_n877), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n876), .B(new_n878), .C1(G150), .C2(new_n718), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n709), .A2(G137), .ZN(new_n880));
  INV_X1    g0680(.A(new_n723), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(G77), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n702), .A2(new_n733), .B1(G50), .B2(new_n692), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n879), .A2(new_n880), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n328), .B1(new_n713), .B2(new_n329), .ZN(new_n885));
  AOI22_X1  g0685(.A1(new_n718), .A2(G303), .B1(new_n692), .B2(G283), .ZN(new_n886));
  XNOR2_X1  g0686(.A(KEYINPUT105), .B(G311), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n886), .B1(new_n697), .B2(new_n887), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n885), .B(new_n888), .C1(G97), .C2(new_n881), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n729), .A2(KEYINPUT46), .A3(G116), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT46), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n711), .B2(new_n207), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n890), .B(new_n892), .C1(new_n471), .C2(new_n701), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT106), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n894), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n889), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n708), .A2(new_n703), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n884), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT107), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n900), .B(KEYINPUT47), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n741), .ZN(new_n902));
  INV_X1    g0702(.A(new_n690), .ZN(new_n903));
  INV_X1    g0703(.A(new_n743), .ZN(new_n904));
  OAI221_X1 g0704(.A(new_n751), .B1(new_n223), .B2(new_n319), .C1(new_n234), .C2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n581), .A2(new_n582), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n629), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n584), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(new_n578), .B2(new_n907), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n909), .A2(new_n753), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n902), .A2(new_n903), .A3(new_n905), .A4(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n685), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n636), .A2(G330), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n639), .A2(new_n643), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n644), .A2(new_n645), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n913), .B(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n547), .A2(new_n629), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n550), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n597), .A2(new_n629), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n646), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT45), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n646), .A2(new_n921), .B1(KEYINPUT104), .B2(KEYINPUT44), .ZN(new_n924));
  OR2_X1    g0724(.A1(KEYINPUT104), .A2(KEYINPUT44), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n923), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n641), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n640), .A2(new_n923), .A3(new_n927), .A4(new_n926), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n917), .A2(new_n929), .A3(new_n682), .A4(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n682), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n652), .B(KEYINPUT41), .Z(new_n933));
  AOI21_X1  g0733(.A(new_n912), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n915), .A2(new_n550), .A3(new_n918), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT103), .ZN(new_n936));
  OR3_X1    g0736(.A1(new_n935), .A2(new_n936), .A3(KEYINPUT42), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(KEYINPUT42), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n936), .B1(new_n935), .B2(KEYINPUT42), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n549), .B1(new_n919), .B2(new_n487), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n630), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n937), .A2(new_n938), .A3(new_n939), .A4(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n921), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n636), .A2(G330), .A3(new_n639), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n909), .A2(KEYINPUT43), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n942), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n909), .A2(KEYINPUT43), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n944), .B1(new_n942), .B2(new_n945), .ZN(new_n950));
  OR3_X1    g0750(.A1(new_n947), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n949), .B1(new_n947), .B2(new_n950), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n911), .B1(new_n934), .B2(new_n953), .ZN(G387));
  AOI22_X1  g0754(.A1(new_n696), .A2(G322), .B1(new_n692), .B2(G303), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n955), .B1(new_n703), .B2(new_n717), .C1(new_n701), .C2(new_n887), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT48), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n711), .A2(new_n471), .B1(new_n713), .B2(new_n726), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT108), .Z(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(KEYINPUT49), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n266), .B1(new_n881), .B2(G116), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n961), .B(new_n962), .C1(new_n698), .C2(new_n708), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n729), .A2(G77), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n964), .B1(new_n778), .B2(new_n212), .C1(new_n202), .C2(new_n717), .ZN(new_n965));
  INV_X1    g0765(.A(G159), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n266), .B1(new_n708), .B2(new_n358), .C1(new_n697), .C2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n713), .A2(new_n319), .ZN(new_n968));
  NOR3_X1   g0768(.A1(new_n965), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n969), .B1(new_n320), .B2(new_n701), .C1(new_n725), .C2(new_n503), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n963), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n690), .B1(new_n971), .B2(new_n741), .ZN(new_n972));
  OR3_X1    g0772(.A1(new_n320), .A2(KEYINPUT50), .A3(G50), .ZN(new_n973));
  OAI21_X1  g0773(.A(KEYINPUT50), .B1(new_n320), .B2(G50), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n973), .A2(new_n974), .A3(new_n475), .A4(new_n653), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G68), .B2(G77), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n743), .B1(new_n231), .B2(new_n475), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n266), .B(new_n223), .C1(G116), .C2(new_n554), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n223), .A2(G107), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n751), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n972), .B(new_n981), .C1(new_n639), .C2(new_n753), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(new_n917), .B2(new_n912), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n917), .A2(new_n682), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n652), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n917), .B2(new_n682), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n984), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(KEYINPUT109), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT109), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n991), .B(new_n984), .C1(new_n986), .C2(new_n988), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n990), .A2(new_n992), .ZN(G393));
  NAND2_X1  g0793(.A1(new_n929), .A2(new_n930), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n985), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n995), .A2(new_n987), .A3(new_n931), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n929), .A2(new_n912), .A3(new_n930), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n751), .B1(new_n503), .B2(new_n223), .C1(new_n239), .C2(new_n904), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n877), .A2(new_n708), .B1(new_n711), .B2(new_n212), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT110), .Z(new_n1000));
  OAI22_X1  g0800(.A1(new_n778), .A2(new_n320), .B1(new_n713), .B2(new_n301), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n328), .B(new_n1001), .C1(G50), .C2(new_n702), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n697), .A2(new_n358), .B1(new_n717), .B2(new_n966), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT51), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n775), .A2(new_n1000), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n328), .B1(new_n713), .B2(new_n207), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n729), .A2(G283), .B1(G294), .B2(new_n692), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n491), .B2(new_n701), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1006), .B(new_n1008), .C1(G322), .C2(new_n709), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n725), .B2(new_n329), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n718), .A2(G311), .B1(new_n696), .B2(G317), .ZN(new_n1011));
  XOR2_X1   g0811(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n1012));
  XNOR2_X1  g0812(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1005), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n690), .B1(new_n1014), .B2(new_n741), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n998), .B(new_n1015), .C1(new_n943), .C2(new_n753), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n997), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n996), .A2(new_n1017), .ZN(G390));
  NAND4_X1  g0818(.A1(new_n818), .A2(new_n767), .A3(new_n819), .A4(new_n840), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n818), .A2(new_n819), .B1(new_n767), .B2(new_n840), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n1020), .A2(new_n1021), .B1(new_n769), .B2(new_n765), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n769), .A2(new_n765), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1023), .A2(new_n842), .A3(new_n1019), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n349), .A2(new_n435), .A3(new_n681), .A4(G330), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n621), .A2(new_n863), .A3(new_n433), .A4(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n842), .A2(new_n858), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1029), .A2(new_n848), .A3(new_n857), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n842), .A2(new_n858), .A3(new_n831), .A4(new_n830), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1023), .A2(new_n820), .ZN(new_n1032));
  AND3_X1   g0832(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1032), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1028), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(KEYINPUT112), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT112), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1037), .B(new_n1028), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n652), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1032), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1030), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n864), .A2(new_n1024), .A3(new_n1022), .A4(new_n1026), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n749), .B1(new_n848), .B2(new_n857), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n718), .A2(G132), .B1(new_n696), .B2(G128), .ZN(new_n1047));
  XOR2_X1   g0847(.A(KEYINPUT54), .B(G143), .Z(new_n1048));
  NAND2_X1  g0848(.A1(new_n692), .A2(new_n1048), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1047), .B(new_n1049), .C1(new_n786), .C2(new_n701), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n328), .B(new_n1050), .C1(G159), .C2(new_n714), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n881), .A2(G50), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n709), .A2(G125), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n711), .A2(new_n358), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1054), .B(new_n1055), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .A4(new_n1056), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n697), .A2(new_n726), .B1(new_n778), .B2(new_n503), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G107), .B2(new_n702), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT115), .Z(new_n1060));
  NAND2_X1  g0860(.A1(new_n729), .A2(G87), .ZN(new_n1061));
  AND3_X1   g0861(.A1(new_n1061), .A2(KEYINPUT116), .A3(new_n328), .ZN(new_n1062));
  AOI21_X1  g0862(.A(KEYINPUT116), .B1(new_n1061), .B2(new_n328), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n717), .A2(new_n207), .B1(new_n713), .B2(new_n301), .ZN(new_n1064));
  NOR3_X1   g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1060), .A2(new_n782), .A3(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n708), .A2(new_n471), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1057), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1046), .B1(new_n741), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n690), .B1(new_n320), .B2(new_n795), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT113), .Z(new_n1071));
  AOI22_X1  g0871(.A1(new_n1039), .A2(new_n1045), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(new_n912), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1074), .ZN(G378));
  INV_X1    g0875(.A(new_n1027), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1037), .B1(new_n1073), .B2(new_n1028), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1038), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(G330), .ZN(new_n1080));
  OAI21_X1  g0880(.A(KEYINPUT55), .B1(new_n367), .B2(new_n434), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT55), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n605), .A2(new_n1082), .A3(new_n433), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n431), .A2(new_n802), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT56), .Z(new_n1085));
  NAND3_X1  g0885(.A1(new_n1081), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1085), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n835), .A2(new_n1080), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT118), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1088), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1092), .A2(KEYINPUT118), .A3(new_n1086), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1094), .A2(G330), .A3(new_n822), .A4(new_n834), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n1089), .A2(new_n862), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n862), .B1(new_n1089), .B2(new_n1095), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1079), .A2(new_n1098), .A3(KEYINPUT57), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT57), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1027), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1100), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1099), .A2(new_n1103), .A3(new_n987), .ZN(new_n1104));
  INV_X1    g0904(.A(G128), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n717), .A2(new_n1105), .B1(new_n713), .B2(new_n358), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n729), .A2(new_n1048), .B1(G137), .B2(new_n692), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n791), .B2(new_n701), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1106), .B(new_n1108), .C1(G125), .C2(new_n696), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT59), .ZN(new_n1110));
  AOI21_X1  g0910(.A(G41), .B1(new_n881), .B2(new_n733), .ZN(new_n1111));
  AOI21_X1  g0911(.A(G33), .B1(new_n709), .B2(G124), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n964), .B1(new_n717), .B2(new_n329), .C1(new_n503), .C2(new_n701), .ZN(new_n1114));
  NOR4_X1   g0914(.A1(new_n1114), .A2(G41), .A3(new_n266), .A4(new_n876), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n778), .A2(new_n319), .B1(new_n708), .B2(new_n726), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n881), .B2(G58), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1115), .B(new_n1117), .C1(new_n207), .C2(new_n697), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT58), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n202), .B1(new_n262), .B2(G41), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1113), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n741), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(KEYINPUT117), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n687), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1122), .A2(KEYINPUT117), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1094), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1126), .B1(G50), .B2(new_n796), .C1(new_n1127), .C2(new_n749), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1128), .B1(new_n1102), .B2(new_n685), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1104), .A2(new_n1130), .ZN(G375));
  NAND2_X1  g0931(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1132), .A2(new_n1044), .A3(new_n933), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1022), .A2(new_n1024), .A3(new_n912), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n696), .A2(G294), .B1(new_n692), .B2(G107), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1135), .B1(new_n207), .B2(new_n701), .C1(new_n726), .C2(new_n717), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n708), .A2(new_n491), .B1(new_n319), .B2(new_n713), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n266), .B1(new_n724), .B2(G77), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1136), .B(new_n1137), .C1(new_n1138), .C2(KEYINPUT119), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n1139), .B1(KEYINPUT119), .B2(new_n1138), .C1(new_n503), .C2(new_n711), .ZN(new_n1140));
  NOR2_X1   g0940(.A1(new_n697), .A2(new_n791), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT120), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n1141), .A2(new_n1142), .B1(new_n202), .B2(new_n713), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1141), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n266), .B1(new_n1144), .B2(KEYINPUT120), .ZN(new_n1145));
  AOI211_X1 g0945(.A(new_n1143), .B(new_n1145), .C1(new_n702), .C2(new_n1048), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G128), .A2(new_n709), .B1(new_n729), .B2(G159), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n786), .B2(new_n717), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(G58), .B2(new_n881), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1146), .B(new_n1149), .C1(new_n358), .C2(new_n778), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1140), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n690), .B1(new_n1151), .B2(new_n741), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1152), .B1(G68), .B2(new_n796), .C1(new_n820), .C2(new_n749), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1134), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1133), .A2(new_n1155), .ZN(G381));
  XOR2_X1   g0956(.A(G375), .B(KEYINPUT121), .Z(new_n1157));
  INV_X1    g0957(.A(G378), .ZN(new_n1158));
  NOR4_X1   g0958(.A1(G387), .A2(G393), .A3(G396), .A4(G390), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(G384), .A2(G381), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .A4(new_n1160), .ZN(G407));
  NAND2_X1  g0961(.A1(new_n628), .A2(G213), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n1162), .B(KEYINPUT122), .Z(new_n1163));
  NAND3_X1  g0963(.A1(new_n1157), .A2(new_n1158), .A3(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(G407), .A2(G213), .A3(new_n1164), .ZN(G409));
  XNOR2_X1  g0965(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1104), .A2(G378), .A3(new_n1130), .ZN(new_n1167));
  AND3_X1   g0967(.A1(new_n1079), .A2(new_n1098), .A3(new_n933), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1074), .B(new_n1072), .C1(new_n1168), .C2(new_n1129), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1163), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1132), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1028), .B1(new_n1171), .B2(KEYINPUT60), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT60), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n652), .B1(new_n1132), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT123), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1172), .A2(KEYINPUT123), .A3(new_n1174), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(G384), .B1(new_n1179), .B2(new_n1155), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n799), .B(new_n1154), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1181));
  OAI211_X1 g0981(.A(G2897), .B(new_n1163), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1178), .ZN(new_n1183));
  AOI21_X1  g0983(.A(KEYINPUT123), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1155), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n799), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1179), .A2(G384), .A3(new_n1155), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1162), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(G2897), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1186), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1182), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1166), .B1(new_n1170), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1162), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT62), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1170), .A2(KEYINPUT62), .A3(new_n1195), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1192), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(G390), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(G387), .A2(new_n1201), .ZN(new_n1202));
  OAI211_X1 g1002(.A(G390), .B(new_n911), .C1(new_n934), .C2(new_n953), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1202), .A2(KEYINPUT124), .A3(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(G396), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n990), .A2(new_n1205), .A3(new_n992), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1205), .B1(new_n990), .B2(new_n992), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n934), .A2(new_n953), .ZN(new_n1209));
  INV_X1    g1009(.A(KEYINPUT124), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1209), .A2(new_n1210), .A3(new_n911), .A4(G390), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1204), .A2(new_n1208), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(KEYINPUT125), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT125), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1204), .A2(new_n1214), .A3(new_n1208), .A4(new_n1211), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1202), .B(new_n1203), .C1(new_n1206), .C2(new_n1207), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(KEYINPUT127), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT127), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1216), .A2(new_n1220), .A3(new_n1217), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1170), .A2(KEYINPUT63), .A3(new_n1195), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1188), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1223), .B(new_n1218), .C1(new_n1224), .C2(new_n1191), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT61), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1188), .B(new_n1194), .C1(new_n1167), .C2(new_n1169), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1226), .B1(new_n1227), .B2(KEYINPUT63), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n1200), .A2(new_n1222), .B1(new_n1225), .B2(new_n1228), .ZN(G405));
  NAND2_X1  g1029(.A1(G375), .A2(new_n1158), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(new_n1167), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1195), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1230), .A2(new_n1167), .A3(new_n1194), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1218), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1234), .B(new_n1235), .ZN(G402));
endmodule


