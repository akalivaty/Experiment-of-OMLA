

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732;

  AND2_X1 U371 ( .A1(n709), .A2(n366), .ZN(n598) );
  XNOR2_X1 U372 ( .A(n596), .B(n595), .ZN(n597) );
  OR2_X1 U373 ( .A1(n514), .A2(KEYINPUT34), .ZN(n370) );
  INV_X1 U374 ( .A(G953), .ZN(n719) );
  OR2_X2 U375 ( .A1(n467), .A2(n468), .ZN(n470) );
  XNOR2_X2 U376 ( .A(n457), .B(KEYINPUT4), .ZN(n467) );
  NOR2_X1 U377 ( .A1(G953), .A2(G237), .ZN(n471) );
  XNOR2_X1 U378 ( .A(n430), .B(n429), .ZN(n480) );
  INV_X1 U379 ( .A(KEYINPUT88), .ZN(n349) );
  NOR2_X1 U380 ( .A1(n362), .A2(n702), .ZN(n682) );
  NOR2_X1 U381 ( .A1(n696), .A2(n702), .ZN(n697) );
  AND2_X2 U382 ( .A1(n412), .A2(n653), .ZN(n698) );
  NAND2_X1 U383 ( .A1(n530), .A2(n503), .ZN(n504) );
  AND2_X1 U384 ( .A1(n574), .A2(n408), .ZN(n668) );
  XNOR2_X1 U385 ( .A(n418), .B(n480), .ZN(n703) );
  XNOR2_X1 U386 ( .A(n365), .B(G110), .ZN(n488) );
  XNOR2_X1 U387 ( .A(n360), .B(G107), .ZN(n456) );
  XNOR2_X1 U388 ( .A(G134), .B(G131), .ZN(n468) );
  XNOR2_X1 U389 ( .A(n349), .B(n350), .ZN(n519) );
  NAND2_X1 U390 ( .A1(n522), .A2(n355), .ZN(n350) );
  XNOR2_X1 U391 ( .A(n351), .B(KEYINPUT22), .ZN(n507) );
  NAND2_X1 U392 ( .A1(n522), .A2(n413), .ZN(n351) );
  XNOR2_X1 U393 ( .A(n456), .B(KEYINPUT16), .ZN(n419) );
  XNOR2_X1 U394 ( .A(n383), .B(G137), .ZN(n498) );
  INV_X1 U395 ( .A(KEYINPUT67), .ZN(n383) );
  XOR2_X1 U396 ( .A(G125), .B(G146), .Z(n449) );
  OR2_X1 U397 ( .A1(n679), .A2(n648), .ZN(n435) );
  NOR2_X1 U398 ( .A1(n527), .A2(n526), .ZN(n539) );
  NOR2_X1 U399 ( .A1(n685), .A2(G902), .ZN(n495) );
  XNOR2_X1 U400 ( .A(n449), .B(n392), .ZN(n715) );
  XNOR2_X1 U401 ( .A(n393), .B(G140), .ZN(n392) );
  INV_X1 U402 ( .A(KEYINPUT10), .ZN(n393) );
  NOR2_X1 U403 ( .A1(G902), .A2(G237), .ZN(n434) );
  NOR2_X1 U404 ( .A1(n585), .A2(n676), .ZN(n586) );
  INV_X1 U405 ( .A(KEYINPUT48), .ZN(n407) );
  XNOR2_X1 U406 ( .A(n462), .B(n401), .ZN(n499) );
  INV_X1 U407 ( .A(KEYINPUT8), .ZN(n401) );
  NAND2_X1 U408 ( .A1(G234), .A2(n719), .ZN(n462) );
  INV_X1 U409 ( .A(KEYINPUT103), .ZN(n414) );
  XNOR2_X1 U410 ( .A(n618), .B(KEYINPUT6), .ZN(n511) );
  INV_X1 U411 ( .A(G116), .ZN(n360) );
  XOR2_X1 U412 ( .A(KEYINPUT23), .B(G119), .Z(n497) );
  XNOR2_X1 U413 ( .A(G128), .B(G110), .ZN(n496) );
  AND2_X1 U414 ( .A1(n499), .A2(G221), .ZN(n400) );
  XNOR2_X1 U415 ( .A(n498), .B(KEYINPUT24), .ZN(n403) );
  XOR2_X1 U416 ( .A(G134), .B(KEYINPUT97), .Z(n459) );
  XNOR2_X1 U417 ( .A(KEYINPUT9), .B(KEYINPUT7), .ZN(n458) );
  XNOR2_X1 U418 ( .A(n457), .B(n381), .ZN(n461) );
  XNOR2_X1 U419 ( .A(n382), .B(KEYINPUT98), .ZN(n381) );
  INV_X1 U420 ( .A(G122), .ZN(n382) );
  XNOR2_X1 U421 ( .A(n390), .B(n453), .ZN(n689) );
  XNOR2_X1 U422 ( .A(n452), .B(n391), .ZN(n390) );
  XNOR2_X1 U423 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U424 ( .A(G146), .B(G101), .Z(n492) );
  INV_X1 U425 ( .A(G140), .ZN(n490) );
  NAND2_X1 U426 ( .A1(n486), .A2(n487), .ZN(n716) );
  INV_X1 U427 ( .A(KEYINPUT74), .ZN(n365) );
  XNOR2_X1 U428 ( .A(n703), .B(n415), .ZN(n679) );
  INV_X1 U429 ( .A(KEYINPUT41), .ZN(n542) );
  NOR2_X1 U430 ( .A1(n605), .A2(n607), .ZN(n543) );
  XNOR2_X1 U431 ( .A(n399), .B(n398), .ZN(n592) );
  INV_X1 U432 ( .A(KEYINPUT39), .ZN(n398) );
  NOR2_X1 U433 ( .A1(n578), .A2(n563), .ZN(n399) );
  NOR2_X2 U434 ( .A1(n553), .A2(n554), .ZN(n574) );
  XNOR2_X1 U435 ( .A(n369), .B(n552), .ZN(n553) );
  XNOR2_X1 U436 ( .A(n551), .B(KEYINPUT107), .ZN(n552) );
  XNOR2_X1 U437 ( .A(n502), .B(KEYINPUT25), .ZN(n409) );
  OR2_X1 U438 ( .A1(n700), .A2(G902), .ZN(n410) );
  AND2_X1 U439 ( .A1(n539), .A2(n404), .ZN(n413) );
  NAND2_X1 U440 ( .A1(n698), .A2(G210), .ZN(n411) );
  NOR2_X1 U441 ( .A1(G952), .A2(n719), .ZN(n702) );
  NAND2_X1 U442 ( .A1(n668), .A2(n606), .ZN(n577) );
  NOR2_X1 U443 ( .A1(n577), .A2(KEYINPUT47), .ZN(n576) );
  NAND2_X1 U444 ( .A1(G237), .A2(G234), .ZN(n437) );
  XOR2_X1 U445 ( .A(KEYINPUT73), .B(KEYINPUT5), .Z(n473) );
  XNOR2_X1 U446 ( .A(G116), .B(G146), .ZN(n474) );
  XOR2_X1 U447 ( .A(KEYINPUT89), .B(G137), .Z(n475) );
  INV_X1 U448 ( .A(KEYINPUT44), .ZN(n386) );
  XNOR2_X1 U449 ( .A(G902), .B(KEYINPUT15), .ZN(n647) );
  XOR2_X1 U450 ( .A(KEYINPUT11), .B(G131), .Z(n444) );
  INV_X1 U451 ( .A(n715), .ZN(n391) );
  XNOR2_X1 U452 ( .A(KEYINPUT93), .B(KEYINPUT12), .ZN(n445) );
  XOR2_X1 U453 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n446) );
  XNOR2_X1 U454 ( .A(n433), .B(KEYINPUT18), .ZN(n417) );
  INV_X1 U455 ( .A(KEYINPUT2), .ZN(n366) );
  XNOR2_X1 U456 ( .A(n540), .B(n541), .ZN(n603) );
  INV_X1 U457 ( .A(KEYINPUT38), .ZN(n541) );
  OR2_X1 U458 ( .A1(n556), .A2(n367), .ZN(n557) );
  AND2_X2 U459 ( .A1(n394), .A2(n594), .ZN(n717) );
  XNOR2_X1 U460 ( .A(n395), .B(n407), .ZN(n394) );
  INV_X1 U461 ( .A(G113), .ZN(n429) );
  AND2_X1 U462 ( .A1(n717), .A2(n648), .ZN(n649) );
  NOR2_X1 U463 ( .A1(n376), .A2(n572), .ZN(n513) );
  NOR2_X1 U464 ( .A1(n571), .A2(n572), .ZN(n587) );
  NOR2_X1 U465 ( .A1(n670), .A2(n568), .ZN(n569) );
  AND2_X1 U466 ( .A1(n522), .A2(n638), .ZN(n514) );
  BUF_X1 U467 ( .A(n540), .Z(n363) );
  XNOR2_X1 U468 ( .A(n379), .B(n378), .ZN(n575) );
  INV_X1 U469 ( .A(KEYINPUT19), .ZN(n378) );
  XNOR2_X1 U470 ( .A(n454), .B(n387), .ZN(n527) );
  XNOR2_X1 U471 ( .A(n455), .B(G475), .ZN(n387) );
  BUF_X1 U472 ( .A(n505), .Z(n618) );
  XNOR2_X1 U473 ( .A(n371), .B(n402), .ZN(n700) );
  XNOR2_X1 U474 ( .A(n500), .B(n403), .ZN(n402) );
  XNOR2_X1 U475 ( .A(n400), .B(n715), .ZN(n371) );
  XNOR2_X1 U476 ( .A(n464), .B(n380), .ZN(n695) );
  XNOR2_X1 U477 ( .A(n463), .B(n465), .ZN(n380) );
  XNOR2_X1 U478 ( .A(n421), .B(n489), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n488), .B(n352), .ZN(n489) );
  XNOR2_X1 U480 ( .A(n493), .B(n490), .ZN(n421) );
  XNOR2_X1 U481 ( .A(n555), .B(n364), .ZN(n732) );
  XNOR2_X1 U482 ( .A(KEYINPUT42), .B(KEYINPUT109), .ZN(n364) );
  XNOR2_X1 U483 ( .A(n565), .B(n564), .ZN(n731) );
  NOR2_X1 U484 ( .A1(n588), .A2(n573), .ZN(n676) );
  XNOR2_X1 U485 ( .A(n389), .B(n388), .ZN(n573) );
  XNOR2_X1 U486 ( .A(KEYINPUT36), .B(KEYINPUT110), .ZN(n388) );
  NAND2_X1 U487 ( .A1(n587), .A2(n363), .ZN(n389) );
  INV_X1 U488 ( .A(n575), .ZN(n408) );
  NAND2_X1 U489 ( .A1(n528), .A2(n527), .ZN(n670) );
  NAND2_X1 U490 ( .A1(n374), .A2(n373), .ZN(n372) );
  INV_X1 U491 ( .A(n702), .ZN(n373) );
  XNOR2_X1 U492 ( .A(n654), .B(n358), .ZN(n374) );
  XNOR2_X1 U493 ( .A(n690), .B(n356), .ZN(n691) );
  XNOR2_X1 U494 ( .A(n411), .B(n357), .ZN(n362) );
  XOR2_X1 U495 ( .A(G107), .B(G104), .Z(n352) );
  XOR2_X1 U496 ( .A(KEYINPUT3), .B(G119), .Z(n353) );
  AND2_X1 U497 ( .A1(n544), .A2(n404), .ZN(n354) );
  AND2_X1 U498 ( .A1(n550), .A2(n354), .ZN(n355) );
  XNOR2_X1 U499 ( .A(n520), .B(KEYINPUT90), .ZN(n657) );
  XNOR2_X1 U500 ( .A(n716), .B(n420), .ZN(n685) );
  XOR2_X1 U501 ( .A(n689), .B(n688), .Z(n356) );
  XOR2_X1 U502 ( .A(n681), .B(n680), .Z(n357) );
  XOR2_X1 U503 ( .A(n645), .B(KEYINPUT62), .Z(n358) );
  XOR2_X1 U504 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n359) );
  INV_X1 U505 ( .A(n602), .ZN(n367) );
  NAND2_X1 U506 ( .A1(n540), .A2(n602), .ZN(n379) );
  INV_X1 U507 ( .A(n615), .ZN(n404) );
  NOR2_X1 U508 ( .A1(n559), .A2(n615), .ZN(n406) );
  NAND2_X2 U509 ( .A1(n470), .A2(n469), .ZN(n484) );
  XNOR2_X1 U510 ( .A(n505), .B(KEYINPUT102), .ZN(n556) );
  XNOR2_X1 U511 ( .A(n361), .B(n386), .ZN(n536) );
  NAND2_X1 U512 ( .A1(n518), .A2(n517), .ZN(n361) );
  INV_X1 U513 ( .A(n709), .ZN(n650) );
  XNOR2_X1 U514 ( .A(n372), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U515 ( .A(n508), .B(KEYINPUT64), .ZN(n509) );
  NAND2_X1 U516 ( .A1(n562), .A2(n561), .ZN(n578) );
  XNOR2_X2 U517 ( .A(n442), .B(KEYINPUT0), .ZN(n522) );
  XNOR2_X1 U518 ( .A(n368), .B(KEYINPUT76), .ZN(n601) );
  NOR2_X2 U519 ( .A1(n598), .A2(n597), .ZN(n368) );
  NAND2_X1 U520 ( .A1(n384), .A2(n570), .ZN(n369) );
  NAND2_X1 U521 ( .A1(n515), .A2(n370), .ZN(n375) );
  NOR2_X1 U522 ( .A1(n570), .A2(n615), .ZN(n620) );
  NAND2_X1 U523 ( .A1(n651), .A2(n652), .ZN(n412) );
  XNOR2_X1 U524 ( .A(n416), .B(n432), .ZN(n415) );
  NAND2_X1 U525 ( .A1(n375), .A2(n581), .ZN(n516) );
  XNOR2_X1 U526 ( .A(n521), .B(n414), .ZN(n376) );
  XNOR2_X1 U527 ( .A(n377), .B(n359), .ZN(G75) );
  NAND2_X1 U528 ( .A1(n644), .A2(n719), .ZN(n377) );
  NAND2_X1 U529 ( .A1(n730), .A2(n661), .ZN(n510) );
  XNOR2_X2 U530 ( .A(n504), .B(KEYINPUT32), .ZN(n730) );
  NOR2_X1 U531 ( .A1(n732), .A2(n731), .ZN(n566) );
  XNOR2_X1 U532 ( .A(n543), .B(n542), .ZN(n637) );
  NOR2_X1 U533 ( .A1(n556), .A2(n385), .ZN(n384) );
  INV_X1 U534 ( .A(n567), .ZN(n385) );
  XNOR2_X2 U535 ( .A(n538), .B(n537), .ZN(n709) );
  NAND2_X1 U536 ( .A1(n467), .A2(n468), .ZN(n469) );
  NAND2_X1 U537 ( .A1(n397), .A2(n396), .ZN(n395) );
  XNOR2_X1 U538 ( .A(n586), .B(KEYINPUT68), .ZN(n396) );
  XNOR2_X1 U539 ( .A(n566), .B(KEYINPUT46), .ZN(n397) );
  NAND2_X1 U540 ( .A1(n592), .A2(n667), .ZN(n565) );
  NAND2_X1 U541 ( .A1(n406), .A2(n544), .ZN(n405) );
  NOR2_X1 U542 ( .A1(n405), .A2(n570), .ZN(n560) );
  XNOR2_X2 U543 ( .A(n410), .B(n409), .ZN(n570) );
  NOR2_X2 U544 ( .A1(n575), .A2(n441), .ZN(n442) );
  NAND2_X1 U545 ( .A1(n600), .A2(n650), .ZN(n653) );
  INV_X1 U546 ( .A(n619), .ZN(n588) );
  NAND2_X1 U547 ( .A1(n619), .A2(n620), .ZN(n521) );
  XNOR2_X2 U548 ( .A(n544), .B(KEYINPUT1), .ZN(n619) );
  XNOR2_X1 U549 ( .A(n467), .B(n417), .ZN(n416) );
  XNOR2_X1 U550 ( .A(n427), .B(n419), .ZN(n418) );
  NOR2_X2 U551 ( .A1(n717), .A2(KEYINPUT2), .ZN(n596) );
  XNOR2_X1 U552 ( .A(n449), .B(n431), .ZN(n432) );
  XOR2_X2 U553 ( .A(G122), .B(G104), .Z(n450) );
  XNOR2_X2 U554 ( .A(n495), .B(n494), .ZN(n544) );
  INV_X1 U555 ( .A(n729), .ZN(n517) );
  AND2_X1 U556 ( .A1(n436), .A2(G210), .ZN(n422) );
  INV_X1 U557 ( .A(n678), .ZN(n593) );
  INV_X1 U558 ( .A(KEYINPUT77), .ZN(n595) );
  AND2_X1 U559 ( .A1(n728), .A2(n593), .ZN(n594) );
  INV_X1 U560 ( .A(n647), .ZN(n648) );
  XNOR2_X1 U561 ( .A(n477), .B(n476), .ZN(n478) );
  NAND2_X1 U562 ( .A1(n603), .A2(n602), .ZN(n607) );
  XNOR2_X1 U563 ( .A(n484), .B(n478), .ZN(n479) );
  INV_X1 U564 ( .A(KEYINPUT40), .ZN(n564) );
  NAND2_X1 U565 ( .A1(G234), .A2(n647), .ZN(n423) );
  XNOR2_X1 U566 ( .A(KEYINPUT20), .B(n423), .ZN(n501) );
  NAND2_X1 U567 ( .A1(n501), .A2(G221), .ZN(n426) );
  XNOR2_X1 U568 ( .A(KEYINPUT87), .B(KEYINPUT21), .ZN(n424) );
  XNOR2_X1 U569 ( .A(n424), .B(KEYINPUT86), .ZN(n425) );
  XOR2_X1 U570 ( .A(n426), .B(n425), .Z(n615) );
  XNOR2_X1 U571 ( .A(n488), .B(n450), .ZN(n427) );
  XNOR2_X1 U572 ( .A(KEYINPUT82), .B(G101), .ZN(n428) );
  XNOR2_X1 U573 ( .A(n353), .B(n428), .ZN(n430) );
  XNOR2_X2 U574 ( .A(G143), .B(G128), .ZN(n457) );
  XOR2_X1 U575 ( .A(KEYINPUT83), .B(KEYINPUT17), .Z(n431) );
  NAND2_X1 U576 ( .A1(G224), .A2(n719), .ZN(n433) );
  XOR2_X1 U577 ( .A(KEYINPUT72), .B(n434), .Z(n436) );
  XNOR2_X2 U578 ( .A(n435), .B(n422), .ZN(n540) );
  NAND2_X1 U579 ( .A1(G214), .A2(n436), .ZN(n602) );
  XNOR2_X1 U580 ( .A(n437), .B(KEYINPUT14), .ZN(n439) );
  NAND2_X1 U581 ( .A1(n439), .A2(G952), .ZN(n635) );
  NOR2_X1 U582 ( .A1(n635), .A2(G953), .ZN(n438) );
  XNOR2_X1 U583 ( .A(n438), .B(KEYINPUT84), .ZN(n549) );
  XNOR2_X1 U584 ( .A(G898), .B(KEYINPUT85), .ZN(n708) );
  NAND2_X1 U585 ( .A1(G953), .A2(n708), .ZN(n704) );
  NAND2_X1 U586 ( .A1(G902), .A2(n439), .ZN(n545) );
  NOR2_X1 U587 ( .A1(n704), .A2(n545), .ZN(n440) );
  NOR2_X1 U588 ( .A1(n549), .A2(n440), .ZN(n441) );
  XNOR2_X1 U589 ( .A(KEYINPUT13), .B(KEYINPUT96), .ZN(n455) );
  NAND2_X1 U590 ( .A1(n471), .A2(G214), .ZN(n443) );
  XNOR2_X1 U591 ( .A(n444), .B(n443), .ZN(n448) );
  XNOR2_X1 U592 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U593 ( .A(n448), .B(n447), .Z(n453) );
  XNOR2_X1 U594 ( .A(G143), .B(n450), .ZN(n451) );
  XNOR2_X1 U595 ( .A(n451), .B(G113), .ZN(n452) );
  NOR2_X1 U596 ( .A1(G902), .A2(n689), .ZN(n454) );
  XNOR2_X1 U597 ( .A(n456), .B(KEYINPUT99), .ZN(n465) );
  XNOR2_X1 U598 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U599 ( .A(n461), .B(n460), .Z(n464) );
  NAND2_X1 U600 ( .A1(G217), .A2(n499), .ZN(n463) );
  NOR2_X1 U601 ( .A1(n695), .A2(G902), .ZN(n466) );
  XOR2_X1 U602 ( .A(n466), .B(G478), .Z(n526) );
  NAND2_X1 U603 ( .A1(G210), .A2(n471), .ZN(n472) );
  XNOR2_X1 U604 ( .A(n473), .B(n472), .ZN(n477) );
  XNOR2_X1 U605 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U606 ( .A(n479), .B(n480), .ZN(n645) );
  NOR2_X1 U607 ( .A1(G902), .A2(n645), .ZN(n482) );
  XNOR2_X1 U608 ( .A(KEYINPUT70), .B(G472), .ZN(n481) );
  XNOR2_X1 U609 ( .A(n482), .B(n481), .ZN(n505) );
  NOR2_X2 U610 ( .A1(n507), .A2(n511), .ZN(n530) );
  INV_X1 U611 ( .A(n498), .ZN(n483) );
  NAND2_X1 U612 ( .A1(n484), .A2(n483), .ZN(n487) );
  INV_X1 U613 ( .A(n484), .ZN(n485) );
  NAND2_X1 U614 ( .A1(n485), .A2(n498), .ZN(n486) );
  NAND2_X1 U615 ( .A1(G227), .A2(n719), .ZN(n491) );
  INV_X1 U616 ( .A(G469), .ZN(n494) );
  XNOR2_X1 U617 ( .A(n497), .B(n496), .ZN(n500) );
  NAND2_X1 U618 ( .A1(n501), .A2(G217), .ZN(n502) );
  XNOR2_X1 U619 ( .A(KEYINPUT100), .B(n570), .ZN(n614) );
  AND2_X1 U620 ( .A1(n619), .A2(n614), .ZN(n503) );
  NAND2_X1 U621 ( .A1(n588), .A2(n556), .ZN(n506) );
  NOR2_X1 U622 ( .A1(n507), .A2(n506), .ZN(n508) );
  NAND2_X1 U623 ( .A1(n509), .A2(n570), .ZN(n661) );
  XNOR2_X1 U624 ( .A(n510), .B(KEYINPUT81), .ZN(n518) );
  INV_X1 U625 ( .A(n511), .ZN(n572) );
  XNOR2_X1 U626 ( .A(KEYINPUT33), .B(KEYINPUT69), .ZN(n512) );
  XNOR2_X1 U627 ( .A(n513), .B(n512), .ZN(n638) );
  NAND2_X1 U628 ( .A1(KEYINPUT34), .A2(n514), .ZN(n515) );
  AND2_X1 U629 ( .A1(n527), .A2(n526), .ZN(n581) );
  XNOR2_X1 U630 ( .A(n516), .B(KEYINPUT35), .ZN(n729) );
  NAND2_X1 U631 ( .A1(n519), .A2(n618), .ZN(n520) );
  NOR2_X1 U632 ( .A1(n618), .A2(n521), .ZN(n626) );
  NAND2_X1 U633 ( .A1(n522), .A2(n626), .ZN(n523) );
  XNOR2_X1 U634 ( .A(n523), .B(KEYINPUT91), .ZN(n524) );
  XNOR2_X1 U635 ( .A(KEYINPUT31), .B(n524), .ZN(n673) );
  NAND2_X1 U636 ( .A1(n657), .A2(n673), .ZN(n525) );
  XNOR2_X1 U637 ( .A(n525), .B(KEYINPUT92), .ZN(n529) );
  INV_X1 U638 ( .A(n526), .ZN(n528) );
  NOR2_X1 U639 ( .A1(n528), .A2(n527), .ZN(n662) );
  INV_X1 U640 ( .A(n662), .ZN(n674) );
  NAND2_X1 U641 ( .A1(n670), .A2(n674), .ZN(n606) );
  NAND2_X1 U642 ( .A1(n529), .A2(n606), .ZN(n533) );
  XOR2_X1 U643 ( .A(n530), .B(KEYINPUT80), .Z(n531) );
  NOR2_X1 U644 ( .A1(n614), .A2(n531), .ZN(n532) );
  NAND2_X1 U645 ( .A1(n588), .A2(n532), .ZN(n655) );
  NAND2_X1 U646 ( .A1(n533), .A2(n655), .ZN(n534) );
  XNOR2_X1 U647 ( .A(KEYINPUT101), .B(n534), .ZN(n535) );
  NAND2_X1 U648 ( .A1(n536), .A2(n535), .ZN(n538) );
  INV_X1 U649 ( .A(KEYINPUT45), .ZN(n537) );
  INV_X1 U650 ( .A(n539), .ZN(n605) );
  INV_X1 U651 ( .A(n544), .ZN(n554) );
  OR2_X1 U652 ( .A1(n719), .A2(n545), .ZN(n546) );
  XNOR2_X1 U653 ( .A(KEYINPUT104), .B(n546), .ZN(n547) );
  NOR2_X1 U654 ( .A1(G900), .A2(n547), .ZN(n548) );
  NOR2_X1 U655 ( .A1(n549), .A2(n548), .ZN(n559) );
  NOR2_X1 U656 ( .A1(n559), .A2(n615), .ZN(n567) );
  INV_X1 U657 ( .A(n570), .ZN(n550) );
  XOR2_X1 U658 ( .A(KEYINPUT28), .B(KEYINPUT108), .Z(n551) );
  NAND2_X1 U659 ( .A1(n637), .A2(n574), .ZN(n555) );
  XOR2_X1 U660 ( .A(KEYINPUT106), .B(KEYINPUT30), .Z(n558) );
  XNOR2_X1 U661 ( .A(n558), .B(n557), .ZN(n562) );
  XOR2_X1 U662 ( .A(KEYINPUT75), .B(n560), .Z(n561) );
  INV_X1 U663 ( .A(n603), .ZN(n563) );
  INV_X1 U664 ( .A(n670), .ZN(n667) );
  NAND2_X1 U665 ( .A1(n567), .A2(n602), .ZN(n568) );
  NAND2_X1 U666 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U667 ( .A(n576), .B(KEYINPUT71), .ZN(n584) );
  NAND2_X1 U668 ( .A1(n577), .A2(KEYINPUT47), .ZN(n582) );
  INV_X1 U669 ( .A(n363), .ZN(n579) );
  NOR2_X1 U670 ( .A1(n579), .A2(n578), .ZN(n580) );
  NAND2_X1 U671 ( .A1(n581), .A2(n580), .ZN(n666) );
  AND2_X1 U672 ( .A1(n582), .A2(n666), .ZN(n583) );
  NAND2_X1 U673 ( .A1(n584), .A2(n583), .ZN(n585) );
  AND2_X1 U674 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U675 ( .A(n589), .B(KEYINPUT43), .ZN(n590) );
  NOR2_X1 U676 ( .A1(n363), .A2(n590), .ZN(n591) );
  XNOR2_X1 U677 ( .A(KEYINPUT105), .B(n591), .ZN(n728) );
  AND2_X1 U678 ( .A1(n662), .A2(n592), .ZN(n678) );
  NAND2_X1 U679 ( .A1(n717), .A2(KEYINPUT2), .ZN(n599) );
  XNOR2_X1 U680 ( .A(KEYINPUT79), .B(n599), .ZN(n600) );
  NAND2_X1 U681 ( .A1(n601), .A2(n653), .ZN(n642) );
  NOR2_X1 U682 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U683 ( .A1(n605), .A2(n604), .ZN(n611) );
  INV_X1 U684 ( .A(n606), .ZN(n608) );
  NOR2_X1 U685 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U686 ( .A(n609), .B(KEYINPUT116), .ZN(n610) );
  NOR2_X1 U687 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U688 ( .A(n612), .B(KEYINPUT117), .ZN(n613) );
  NAND2_X1 U689 ( .A1(n613), .A2(n638), .ZN(n632) );
  XNOR2_X1 U690 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n629) );
  AND2_X1 U691 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U692 ( .A(n616), .B(KEYINPUT49), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n618), .A2(n617), .ZN(n623) );
  NOR2_X1 U694 ( .A1(n620), .A2(n619), .ZN(n621) );
  XNOR2_X1 U695 ( .A(n621), .B(KEYINPUT50), .ZN(n622) );
  NOR2_X1 U696 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U697 ( .A(KEYINPUT113), .B(n624), .Z(n625) );
  NOR2_X1 U698 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U699 ( .A(KEYINPUT51), .B(n627), .Z(n628) );
  XNOR2_X1 U700 ( .A(n629), .B(n628), .ZN(n630) );
  NAND2_X1 U701 ( .A1(n630), .A2(n637), .ZN(n631) );
  NAND2_X1 U702 ( .A1(n632), .A2(n631), .ZN(n633) );
  XOR2_X1 U703 ( .A(KEYINPUT52), .B(n633), .Z(n634) );
  NOR2_X1 U704 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U705 ( .A(n636), .B(KEYINPUT118), .ZN(n640) );
  AND2_X1 U706 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U707 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U708 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U709 ( .A(n643), .B(KEYINPUT119), .ZN(n644) );
  XOR2_X1 U710 ( .A(n647), .B(KEYINPUT78), .Z(n646) );
  NAND2_X1 U711 ( .A1(n646), .A2(KEYINPUT2), .ZN(n652) );
  NAND2_X1 U712 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U713 ( .A1(G472), .A2(n698), .ZN(n654) );
  XNOR2_X1 U714 ( .A(G101), .B(n655), .ZN(G3) );
  NOR2_X1 U715 ( .A1(n657), .A2(n670), .ZN(n656) );
  XOR2_X1 U716 ( .A(G104), .B(n656), .Z(G6) );
  NOR2_X1 U717 ( .A1(n657), .A2(n674), .ZN(n659) );
  XNOR2_X1 U718 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n658) );
  XNOR2_X1 U719 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U720 ( .A(G107), .B(n660), .ZN(G9) );
  XNOR2_X1 U721 ( .A(G110), .B(n661), .ZN(G12) );
  XOR2_X1 U722 ( .A(KEYINPUT111), .B(KEYINPUT29), .Z(n664) );
  NAND2_X1 U723 ( .A1(n668), .A2(n662), .ZN(n663) );
  XNOR2_X1 U724 ( .A(n664), .B(n663), .ZN(n665) );
  XOR2_X1 U725 ( .A(G128), .B(n665), .Z(G30) );
  XNOR2_X1 U726 ( .A(G143), .B(n666), .ZN(G45) );
  NAND2_X1 U727 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U728 ( .A(n669), .B(G146), .ZN(G48) );
  NOR2_X1 U729 ( .A1(n670), .A2(n673), .ZN(n671) );
  XOR2_X1 U730 ( .A(KEYINPUT112), .B(n671), .Z(n672) );
  XNOR2_X1 U731 ( .A(G113), .B(n672), .ZN(G15) );
  NOR2_X1 U732 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U733 ( .A(G116), .B(n675), .Z(G18) );
  XNOR2_X1 U734 ( .A(G125), .B(n676), .ZN(n677) );
  XNOR2_X1 U735 ( .A(n677), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U736 ( .A(G134), .B(n678), .Z(G36) );
  XOR2_X1 U737 ( .A(KEYINPUT121), .B(KEYINPUT54), .Z(n681) );
  XNOR2_X1 U738 ( .A(n679), .B(KEYINPUT55), .ZN(n680) );
  XNOR2_X1 U739 ( .A(KEYINPUT56), .B(n682), .ZN(G51) );
  XOR2_X1 U740 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n684) );
  NAND2_X1 U741 ( .A1(n698), .A2(G469), .ZN(n683) );
  XNOR2_X1 U742 ( .A(n684), .B(n683), .ZN(n686) );
  XNOR2_X1 U743 ( .A(n686), .B(n685), .ZN(n687) );
  NOR2_X1 U744 ( .A1(n702), .A2(n687), .ZN(G54) );
  NAND2_X1 U745 ( .A1(n698), .A2(G475), .ZN(n690) );
  XOR2_X1 U746 ( .A(KEYINPUT59), .B(KEYINPUT65), .Z(n688) );
  NOR2_X2 U747 ( .A1(n702), .A2(n691), .ZN(n693) );
  XNOR2_X1 U748 ( .A(KEYINPUT66), .B(KEYINPUT60), .ZN(n692) );
  XNOR2_X1 U749 ( .A(n693), .B(n692), .ZN(G60) );
  NAND2_X1 U750 ( .A1(G478), .A2(n698), .ZN(n694) );
  XNOR2_X1 U751 ( .A(n695), .B(n694), .ZN(n696) );
  XNOR2_X1 U752 ( .A(n697), .B(KEYINPUT122), .ZN(G63) );
  NAND2_X1 U753 ( .A1(G217), .A2(n698), .ZN(n699) );
  XNOR2_X1 U754 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U755 ( .A1(n702), .A2(n701), .ZN(G66) );
  NAND2_X1 U756 ( .A1(n704), .A2(n703), .ZN(n713) );
  NAND2_X1 U757 ( .A1(G224), .A2(G953), .ZN(n705) );
  XNOR2_X1 U758 ( .A(n705), .B(KEYINPUT123), .ZN(n706) );
  XNOR2_X1 U759 ( .A(n706), .B(KEYINPUT61), .ZN(n707) );
  NOR2_X1 U760 ( .A1(n708), .A2(n707), .ZN(n711) );
  NOR2_X1 U761 ( .A1(G953), .A2(n709), .ZN(n710) );
  NOR2_X1 U762 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U763 ( .A(n713), .B(n712), .ZN(n714) );
  XNOR2_X1 U764 ( .A(KEYINPUT124), .B(n714), .ZN(G69) );
  XNOR2_X1 U765 ( .A(n716), .B(n715), .ZN(n722) );
  XNOR2_X1 U766 ( .A(n722), .B(n717), .ZN(n718) );
  XNOR2_X1 U767 ( .A(n718), .B(KEYINPUT125), .ZN(n720) );
  NAND2_X1 U768 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U769 ( .A(n721), .B(KEYINPUT126), .ZN(n726) );
  XNOR2_X1 U770 ( .A(G227), .B(n722), .ZN(n723) );
  NAND2_X1 U771 ( .A1(n723), .A2(G900), .ZN(n724) );
  NAND2_X1 U772 ( .A1(n724), .A2(G953), .ZN(n725) );
  NAND2_X1 U773 ( .A1(n726), .A2(n725), .ZN(n727) );
  XOR2_X1 U774 ( .A(KEYINPUT127), .B(n727), .Z(G72) );
  XNOR2_X1 U775 ( .A(G140), .B(n728), .ZN(G42) );
  XOR2_X1 U776 ( .A(n729), .B(G122), .Z(G24) );
  XNOR2_X1 U777 ( .A(n730), .B(G119), .ZN(G21) );
  XOR2_X1 U778 ( .A(n731), .B(G131), .Z(G33) );
  XOR2_X1 U779 ( .A(n732), .B(G137), .Z(G39) );
endmodule

