

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(G164), .A2(G1384), .ZN(n710) );
  NOR2_X2 U550 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X2 U551 ( .A1(G2105), .A2(n521), .ZN(n584) );
  NOR2_X4 U552 ( .A1(G2105), .A2(G2104), .ZN(n517) );
  AND2_X2 U553 ( .A1(G2104), .A2(G2105), .ZN(n515) );
  NOR2_X2 U554 ( .A1(n614), .A2(n934), .ZN(n626) );
  AND2_X1 U555 ( .A1(n626), .A2(n927), .ZN(n625) );
  INV_X1 U556 ( .A(KEYINPUT17), .ZN(n516) );
  INV_X1 U557 ( .A(KEYINPUT99), .ZN(n634) );
  INV_X1 U558 ( .A(G2104), .ZN(n521) );
  NOR2_X1 U559 ( .A1(G651), .A2(G543), .ZN(n802) );
  XOR2_X1 U560 ( .A(KEYINPUT1), .B(n527), .Z(n808) );
  NOR2_X1 U561 ( .A1(G651), .A2(n561), .ZN(n806) );
  NAND2_X1 U562 ( .A1(n717), .A2(G137), .ZN(n595) );
  NOR2_X1 U563 ( .A1(n525), .A2(n524), .ZN(G164) );
  XNOR2_X2 U564 ( .A(n517), .B(n516), .ZN(n717) );
  NAND2_X1 U565 ( .A1(n717), .A2(G138), .ZN(n520) );
  NAND2_X1 U566 ( .A1(G114), .A2(n515), .ZN(n518) );
  XOR2_X1 U567 ( .A(KEYINPUT87), .B(n518), .Z(n519) );
  NAND2_X1 U568 ( .A1(n520), .A2(n519), .ZN(n525) );
  BUF_X1 U569 ( .A(n584), .Z(n895) );
  NAND2_X1 U570 ( .A1(G102), .A2(n895), .ZN(n523) );
  AND2_X2 U571 ( .A1(n521), .A2(G2105), .ZN(n898) );
  NAND2_X1 U572 ( .A1(G126), .A2(n898), .ZN(n522) );
  NAND2_X1 U573 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U574 ( .A(KEYINPUT0), .B(G543), .Z(n561) );
  INV_X1 U575 ( .A(G651), .ZN(n526) );
  NOR2_X1 U576 ( .A1(n561), .A2(n526), .ZN(n803) );
  NAND2_X1 U577 ( .A1(G78), .A2(n803), .ZN(n529) );
  NOR2_X1 U578 ( .A1(G543), .A2(n526), .ZN(n527) );
  NAND2_X1 U579 ( .A1(G65), .A2(n808), .ZN(n528) );
  NAND2_X1 U580 ( .A1(n529), .A2(n528), .ZN(n532) );
  NAND2_X1 U581 ( .A1(n802), .A2(G91), .ZN(n530) );
  XOR2_X1 U582 ( .A(KEYINPUT68), .B(n530), .Z(n531) );
  NOR2_X1 U583 ( .A1(n532), .A2(n531), .ZN(n534) );
  NAND2_X1 U584 ( .A1(n806), .A2(G53), .ZN(n533) );
  NAND2_X1 U585 ( .A1(n534), .A2(n533), .ZN(G299) );
  NAND2_X1 U586 ( .A1(G90), .A2(n802), .ZN(n536) );
  NAND2_X1 U587 ( .A1(G77), .A2(n803), .ZN(n535) );
  NAND2_X1 U588 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U589 ( .A(KEYINPUT9), .B(n537), .ZN(n541) );
  NAND2_X1 U590 ( .A1(G64), .A2(n808), .ZN(n539) );
  NAND2_X1 U591 ( .A1(G52), .A2(n806), .ZN(n538) );
  AND2_X1 U592 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U593 ( .A1(n541), .A2(n540), .ZN(G301) );
  INV_X1 U594 ( .A(G301), .ZN(G171) );
  NAND2_X1 U595 ( .A1(G63), .A2(n808), .ZN(n543) );
  NAND2_X1 U596 ( .A1(G51), .A2(n806), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n543), .A2(n542), .ZN(n545) );
  XOR2_X1 U598 ( .A(KEYINPUT73), .B(KEYINPUT6), .Z(n544) );
  XNOR2_X1 U599 ( .A(n545), .B(n544), .ZN(n553) );
  XNOR2_X1 U600 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n551) );
  NAND2_X1 U601 ( .A1(n802), .A2(G89), .ZN(n546) );
  XNOR2_X1 U602 ( .A(n546), .B(KEYINPUT4), .ZN(n548) );
  NAND2_X1 U603 ( .A1(G76), .A2(n803), .ZN(n547) );
  NAND2_X1 U604 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U605 ( .A(n549), .B(KEYINPUT5), .ZN(n550) );
  XNOR2_X1 U606 ( .A(n551), .B(n550), .ZN(n552) );
  NOR2_X1 U607 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U608 ( .A(KEYINPUT7), .B(n554), .Z(G168) );
  XOR2_X1 U609 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U610 ( .A1(G88), .A2(n802), .ZN(n556) );
  NAND2_X1 U611 ( .A1(G75), .A2(n803), .ZN(n555) );
  NAND2_X1 U612 ( .A1(n556), .A2(n555), .ZN(n560) );
  NAND2_X1 U613 ( .A1(G62), .A2(n808), .ZN(n558) );
  NAND2_X1 U614 ( .A1(G50), .A2(n806), .ZN(n557) );
  NAND2_X1 U615 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U616 ( .A1(n560), .A2(n559), .ZN(G166) );
  INV_X1 U617 ( .A(G166), .ZN(G303) );
  NAND2_X1 U618 ( .A1(G49), .A2(n806), .ZN(n563) );
  NAND2_X1 U619 ( .A1(G87), .A2(n561), .ZN(n562) );
  NAND2_X1 U620 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U621 ( .A1(n808), .A2(n564), .ZN(n567) );
  NAND2_X1 U622 ( .A1(G74), .A2(G651), .ZN(n565) );
  XOR2_X1 U623 ( .A(KEYINPUT77), .B(n565), .Z(n566) );
  NAND2_X1 U624 ( .A1(n567), .A2(n566), .ZN(G288) );
  XOR2_X1 U625 ( .A(KEYINPUT78), .B(KEYINPUT2), .Z(n569) );
  NAND2_X1 U626 ( .A1(G73), .A2(n803), .ZN(n568) );
  XNOR2_X1 U627 ( .A(n569), .B(n568), .ZN(n573) );
  NAND2_X1 U628 ( .A1(G86), .A2(n802), .ZN(n571) );
  NAND2_X1 U629 ( .A1(G61), .A2(n808), .ZN(n570) );
  NAND2_X1 U630 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U631 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U632 ( .A(KEYINPUT79), .B(n574), .Z(n576) );
  NAND2_X1 U633 ( .A1(n806), .A2(G48), .ZN(n575) );
  NAND2_X1 U634 ( .A1(n576), .A2(n575), .ZN(G305) );
  NAND2_X1 U635 ( .A1(G85), .A2(n802), .ZN(n578) );
  NAND2_X1 U636 ( .A1(G72), .A2(n803), .ZN(n577) );
  NAND2_X1 U637 ( .A1(n578), .A2(n577), .ZN(n581) );
  NAND2_X1 U638 ( .A1(G47), .A2(n806), .ZN(n579) );
  XOR2_X1 U639 ( .A(KEYINPUT66), .B(n579), .Z(n580) );
  NOR2_X1 U640 ( .A1(n581), .A2(n580), .ZN(n583) );
  NAND2_X1 U641 ( .A1(n808), .A2(G60), .ZN(n582) );
  NAND2_X1 U642 ( .A1(n583), .A2(n582), .ZN(G290) );
  INV_X1 U643 ( .A(KEYINPUT23), .ZN(n586) );
  NAND2_X1 U644 ( .A1(n584), .A2(G101), .ZN(n585) );
  XNOR2_X1 U645 ( .A(n586), .B(n585), .ZN(n588) );
  NAND2_X1 U646 ( .A1(n898), .A2(G125), .ZN(n587) );
  NAND2_X1 U647 ( .A1(n588), .A2(n587), .ZN(n591) );
  INV_X1 U648 ( .A(n591), .ZN(n590) );
  INV_X1 U649 ( .A(KEYINPUT65), .ZN(n589) );
  NAND2_X1 U650 ( .A1(n590), .A2(n589), .ZN(n593) );
  NAND2_X1 U651 ( .A1(KEYINPUT65), .A2(n591), .ZN(n592) );
  NAND2_X1 U652 ( .A1(n593), .A2(n592), .ZN(n765) );
  NAND2_X1 U653 ( .A1(n515), .A2(G113), .ZN(n594) );
  AND2_X1 U654 ( .A1(n595), .A2(n594), .ZN(n766) );
  AND2_X1 U655 ( .A1(G40), .A2(n766), .ZN(n596) );
  NAND2_X1 U656 ( .A1(n765), .A2(n596), .ZN(n597) );
  XNOR2_X1 U657 ( .A(n597), .B(KEYINPUT88), .ZN(n711) );
  INV_X1 U658 ( .A(n710), .ZN(n598) );
  NOR2_X2 U659 ( .A1(n711), .A2(n598), .ZN(n599) );
  XNOR2_X2 U660 ( .A(n599), .B(KEYINPUT64), .ZN(n601) );
  NAND2_X1 U661 ( .A1(n601), .A2(G1996), .ZN(n600) );
  XNOR2_X1 U662 ( .A(n600), .B(KEYINPUT26), .ZN(n603) );
  INV_X2 U663 ( .A(n601), .ZN(n659) );
  NAND2_X1 U664 ( .A1(G1341), .A2(n659), .ZN(n602) );
  NAND2_X1 U665 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U666 ( .A(n604), .B(KEYINPUT98), .ZN(n614) );
  NAND2_X1 U667 ( .A1(G56), .A2(n808), .ZN(n605) );
  XOR2_X1 U668 ( .A(KEYINPUT14), .B(n605), .Z(n611) );
  NAND2_X1 U669 ( .A1(n802), .A2(G81), .ZN(n606) );
  XNOR2_X1 U670 ( .A(n606), .B(KEYINPUT12), .ZN(n608) );
  NAND2_X1 U671 ( .A1(G68), .A2(n803), .ZN(n607) );
  NAND2_X1 U672 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U673 ( .A(KEYINPUT13), .B(n609), .Z(n610) );
  NOR2_X1 U674 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U675 ( .A1(n806), .A2(G43), .ZN(n612) );
  NAND2_X1 U676 ( .A1(n613), .A2(n612), .ZN(n934) );
  NAND2_X1 U677 ( .A1(G92), .A2(n802), .ZN(n616) );
  NAND2_X1 U678 ( .A1(G66), .A2(n808), .ZN(n615) );
  NAND2_X1 U679 ( .A1(n616), .A2(n615), .ZN(n620) );
  NAND2_X1 U680 ( .A1(G79), .A2(n803), .ZN(n618) );
  NAND2_X1 U681 ( .A1(G54), .A2(n806), .ZN(n617) );
  NAND2_X1 U682 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U683 ( .A1(n620), .A2(n619), .ZN(n621) );
  XOR2_X1 U684 ( .A(KEYINPUT15), .B(n621), .Z(n927) );
  OR2_X1 U685 ( .A1(n659), .A2(G2067), .ZN(n623) );
  INV_X1 U686 ( .A(n659), .ZN(n642) );
  OR2_X1 U687 ( .A1(G1348), .A2(n642), .ZN(n622) );
  NAND2_X1 U688 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U689 ( .A1(n625), .A2(n624), .ZN(n628) );
  NOR2_X1 U690 ( .A1(n927), .A2(n626), .ZN(n627) );
  NOR2_X1 U691 ( .A1(n628), .A2(n627), .ZN(n633) );
  NAND2_X1 U692 ( .A1(G2072), .A2(n642), .ZN(n629) );
  XOR2_X1 U693 ( .A(KEYINPUT27), .B(n629), .Z(n631) );
  NAND2_X1 U694 ( .A1(n659), .A2(G1956), .ZN(n630) );
  NAND2_X1 U695 ( .A1(n631), .A2(n630), .ZN(n636) );
  NOR2_X1 U696 ( .A1(n636), .A2(G299), .ZN(n632) );
  NOR2_X1 U697 ( .A1(n633), .A2(n632), .ZN(n635) );
  XNOR2_X1 U698 ( .A(n635), .B(n634), .ZN(n640) );
  XOR2_X1 U699 ( .A(KEYINPUT97), .B(KEYINPUT28), .Z(n638) );
  NAND2_X1 U700 ( .A1(G299), .A2(n636), .ZN(n637) );
  XOR2_X1 U701 ( .A(n638), .B(n637), .Z(n639) );
  XNOR2_X1 U702 ( .A(n641), .B(KEYINPUT29), .ZN(n647) );
  NAND2_X1 U703 ( .A1(n659), .A2(G1961), .ZN(n644) );
  XOR2_X1 U704 ( .A(G2078), .B(KEYINPUT25), .Z(n977) );
  NAND2_X1 U705 ( .A1(n977), .A2(n642), .ZN(n643) );
  NAND2_X1 U706 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U707 ( .A(KEYINPUT96), .B(n645), .Z(n653) );
  NAND2_X1 U708 ( .A1(G171), .A2(n653), .ZN(n646) );
  NAND2_X1 U709 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U710 ( .A(n648), .B(KEYINPUT100), .ZN(n658) );
  NAND2_X1 U711 ( .A1(n659), .A2(G8), .ZN(n705) );
  NOR2_X1 U712 ( .A1(G1966), .A2(n705), .ZN(n672) );
  NOR2_X1 U713 ( .A1(n659), .A2(G2084), .ZN(n674) );
  NOR2_X1 U714 ( .A1(n672), .A2(n674), .ZN(n649) );
  NAND2_X1 U715 ( .A1(G8), .A2(n649), .ZN(n650) );
  XNOR2_X1 U716 ( .A(KEYINPUT30), .B(n650), .ZN(n651) );
  XOR2_X1 U717 ( .A(KEYINPUT101), .B(n651), .Z(n652) );
  NOR2_X1 U718 ( .A1(G168), .A2(n652), .ZN(n655) );
  NOR2_X1 U719 ( .A1(G171), .A2(n653), .ZN(n654) );
  NOR2_X1 U720 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U721 ( .A(KEYINPUT31), .B(n656), .Z(n657) );
  NAND2_X1 U722 ( .A1(n658), .A2(n657), .ZN(n671) );
  NAND2_X1 U723 ( .A1(n671), .A2(G286), .ZN(n667) );
  INV_X1 U724 ( .A(G8), .ZN(n665) );
  NOR2_X1 U725 ( .A1(n659), .A2(G2090), .ZN(n661) );
  NOR2_X1 U726 ( .A1(G1971), .A2(n705), .ZN(n660) );
  NOR2_X1 U727 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U728 ( .A(n662), .B(KEYINPUT102), .ZN(n663) );
  NAND2_X1 U729 ( .A1(n663), .A2(G303), .ZN(n664) );
  OR2_X1 U730 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U731 ( .A1(n667), .A2(n666), .ZN(n669) );
  INV_X1 U732 ( .A(KEYINPUT32), .ZN(n668) );
  XNOR2_X1 U733 ( .A(n669), .B(n668), .ZN(n695) );
  INV_X1 U734 ( .A(n705), .ZN(n670) );
  NAND2_X1 U735 ( .A1(n695), .A2(n670), .ZN(n678) );
  INV_X1 U736 ( .A(n671), .ZN(n673) );
  NOR2_X1 U737 ( .A1(n673), .A2(n672), .ZN(n676) );
  NAND2_X1 U738 ( .A1(G8), .A2(n674), .ZN(n675) );
  NAND2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n697) );
  NAND2_X1 U740 ( .A1(G1976), .A2(G288), .ZN(n932) );
  NAND2_X1 U741 ( .A1(n697), .A2(n932), .ZN(n677) );
  NOR2_X1 U742 ( .A1(n678), .A2(n677), .ZN(n687) );
  INV_X1 U743 ( .A(n932), .ZN(n682) );
  NOR2_X1 U744 ( .A1(G288), .A2(G1976), .ZN(n679) );
  XNOR2_X1 U745 ( .A(n679), .B(KEYINPUT103), .ZN(n689) );
  INV_X1 U746 ( .A(n689), .ZN(n681) );
  NOR2_X1 U747 ( .A1(G1971), .A2(G303), .ZN(n680) );
  NOR2_X1 U748 ( .A1(n681), .A2(n680), .ZN(n926) );
  OR2_X1 U749 ( .A1(n682), .A2(n926), .ZN(n683) );
  OR2_X1 U750 ( .A1(n705), .A2(n683), .ZN(n685) );
  INV_X1 U751 ( .A(KEYINPUT33), .ZN(n684) );
  NAND2_X1 U752 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U753 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U754 ( .A(n688), .B(KEYINPUT104), .ZN(n693) );
  XOR2_X1 U755 ( .A(G1981), .B(G305), .Z(n922) );
  NOR2_X1 U756 ( .A1(n705), .A2(n689), .ZN(n690) );
  NAND2_X1 U757 ( .A1(KEYINPUT33), .A2(n690), .ZN(n691) );
  NAND2_X1 U758 ( .A1(n922), .A2(n691), .ZN(n692) );
  NOR2_X2 U759 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U760 ( .A(n694), .B(KEYINPUT105), .ZN(n709) );
  BUF_X1 U761 ( .A(n695), .Z(n696) );
  NAND2_X1 U762 ( .A1(n697), .A2(n696), .ZN(n700) );
  NOR2_X1 U763 ( .A1(G2090), .A2(G303), .ZN(n698) );
  NAND2_X1 U764 ( .A1(G8), .A2(n698), .ZN(n699) );
  NAND2_X1 U765 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U766 ( .A1(n705), .A2(n701), .ZN(n702) );
  XNOR2_X1 U767 ( .A(KEYINPUT106), .B(n702), .ZN(n707) );
  NOR2_X1 U768 ( .A1(G1981), .A2(G305), .ZN(n703) );
  XOR2_X1 U769 ( .A(n703), .B(KEYINPUT24), .Z(n704) );
  OR2_X1 U770 ( .A1(n705), .A2(n704), .ZN(n706) );
  AND2_X1 U771 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U772 ( .A1(n709), .A2(n708), .ZN(n748) );
  NOR2_X1 U773 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U774 ( .A(KEYINPUT89), .B(n712), .Z(n759) );
  XOR2_X1 U775 ( .A(G2067), .B(KEYINPUT37), .Z(n713) );
  XOR2_X1 U776 ( .A(KEYINPUT90), .B(n713), .Z(n757) );
  NAND2_X1 U777 ( .A1(G128), .A2(n898), .ZN(n715) );
  NAND2_X1 U778 ( .A1(G116), .A2(n515), .ZN(n714) );
  NAND2_X1 U779 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U780 ( .A(n716), .B(KEYINPUT35), .ZN(n722) );
  NAND2_X1 U781 ( .A1(G104), .A2(n895), .ZN(n719) );
  NAND2_X1 U782 ( .A1(G140), .A2(n717), .ZN(n718) );
  NAND2_X1 U783 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U784 ( .A(KEYINPUT34), .B(n720), .Z(n721) );
  NAND2_X1 U785 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U786 ( .A(n723), .B(KEYINPUT36), .Z(n908) );
  OR2_X1 U787 ( .A1(n757), .A2(n908), .ZN(n724) );
  XNOR2_X1 U788 ( .A(n724), .B(KEYINPUT91), .ZN(n1009) );
  NAND2_X1 U789 ( .A1(n759), .A2(n1009), .ZN(n755) );
  INV_X1 U790 ( .A(n755), .ZN(n743) );
  XOR2_X1 U791 ( .A(KEYINPUT93), .B(n759), .Z(n741) );
  NAND2_X1 U792 ( .A1(G119), .A2(n898), .ZN(n726) );
  NAND2_X1 U793 ( .A1(G107), .A2(n515), .ZN(n725) );
  NAND2_X1 U794 ( .A1(n726), .A2(n725), .ZN(n730) );
  NAND2_X1 U795 ( .A1(G95), .A2(n895), .ZN(n728) );
  NAND2_X1 U796 ( .A1(G131), .A2(n717), .ZN(n727) );
  NAND2_X1 U797 ( .A1(n728), .A2(n727), .ZN(n729) );
  OR2_X1 U798 ( .A1(n730), .A2(n729), .ZN(n890) );
  NAND2_X1 U799 ( .A1(G1991), .A2(n890), .ZN(n740) );
  XOR2_X1 U800 ( .A(KEYINPUT38), .B(KEYINPUT92), .Z(n732) );
  NAND2_X1 U801 ( .A1(G105), .A2(n895), .ZN(n731) );
  XNOR2_X1 U802 ( .A(n732), .B(n731), .ZN(n736) );
  NAND2_X1 U803 ( .A1(G129), .A2(n898), .ZN(n734) );
  NAND2_X1 U804 ( .A1(G117), .A2(n515), .ZN(n733) );
  NAND2_X1 U805 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U806 ( .A1(n736), .A2(n735), .ZN(n738) );
  NAND2_X1 U807 ( .A1(n717), .A2(G141), .ZN(n737) );
  NAND2_X1 U808 ( .A1(n738), .A2(n737), .ZN(n888) );
  NAND2_X1 U809 ( .A1(G1996), .A2(n888), .ZN(n739) );
  NAND2_X1 U810 ( .A1(n740), .A2(n739), .ZN(n996) );
  NAND2_X1 U811 ( .A1(n741), .A2(n996), .ZN(n742) );
  XOR2_X1 U812 ( .A(KEYINPUT94), .B(n742), .Z(n752) );
  NOR2_X1 U813 ( .A1(n743), .A2(n752), .ZN(n744) );
  XOR2_X1 U814 ( .A(n744), .B(KEYINPUT95), .Z(n746) );
  XNOR2_X1 U815 ( .A(G1986), .B(G290), .ZN(n931) );
  NAND2_X1 U816 ( .A1(n931), .A2(n759), .ZN(n745) );
  AND2_X1 U817 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U818 ( .A1(n748), .A2(n747), .ZN(n762) );
  NOR2_X1 U819 ( .A1(G1996), .A2(n888), .ZN(n1001) );
  NOR2_X1 U820 ( .A1(G1991), .A2(n890), .ZN(n749) );
  XOR2_X1 U821 ( .A(KEYINPUT107), .B(n749), .Z(n997) );
  NOR2_X1 U822 ( .A1(G1986), .A2(G290), .ZN(n750) );
  NOR2_X1 U823 ( .A1(n997), .A2(n750), .ZN(n751) );
  NOR2_X1 U824 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U825 ( .A1(n1001), .A2(n753), .ZN(n754) );
  XNOR2_X1 U826 ( .A(n754), .B(KEYINPUT39), .ZN(n756) );
  NAND2_X1 U827 ( .A1(n756), .A2(n755), .ZN(n758) );
  NAND2_X1 U828 ( .A1(n757), .A2(n908), .ZN(n1017) );
  NAND2_X1 U829 ( .A1(n758), .A2(n1017), .ZN(n760) );
  NAND2_X1 U830 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U831 ( .A1(n762), .A2(n761), .ZN(n764) );
  XNOR2_X1 U832 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n763) );
  XNOR2_X1 U833 ( .A(n764), .B(n763), .ZN(G329) );
  AND2_X1 U834 ( .A1(n766), .A2(n765), .ZN(G160) );
  XNOR2_X1 U835 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U836 ( .A(G2443), .B(G2446), .Z(n768) );
  XNOR2_X1 U837 ( .A(G2427), .B(G2451), .ZN(n767) );
  XNOR2_X1 U838 ( .A(n768), .B(n767), .ZN(n774) );
  XOR2_X1 U839 ( .A(G2430), .B(G2454), .Z(n770) );
  XNOR2_X1 U840 ( .A(G1348), .B(G1341), .ZN(n769) );
  XNOR2_X1 U841 ( .A(n770), .B(n769), .ZN(n772) );
  XOR2_X1 U842 ( .A(G2435), .B(G2438), .Z(n771) );
  XNOR2_X1 U843 ( .A(n772), .B(n771), .ZN(n773) );
  XOR2_X1 U844 ( .A(n774), .B(n773), .Z(n775) );
  AND2_X1 U845 ( .A1(G14), .A2(n775), .ZN(G401) );
  NAND2_X1 U846 ( .A1(G123), .A2(n898), .ZN(n776) );
  XNOR2_X1 U847 ( .A(n776), .B(KEYINPUT18), .ZN(n783) );
  NAND2_X1 U848 ( .A1(G111), .A2(n515), .ZN(n778) );
  NAND2_X1 U849 ( .A1(G135), .A2(n717), .ZN(n777) );
  NAND2_X1 U850 ( .A1(n778), .A2(n777), .ZN(n781) );
  NAND2_X1 U851 ( .A1(G99), .A2(n895), .ZN(n779) );
  XNOR2_X1 U852 ( .A(KEYINPUT75), .B(n779), .ZN(n780) );
  NOR2_X1 U853 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U854 ( .A1(n783), .A2(n782), .ZN(n998) );
  XNOR2_X1 U855 ( .A(G2096), .B(n998), .ZN(n784) );
  OR2_X1 U856 ( .A1(G2100), .A2(n784), .ZN(G156) );
  INV_X1 U857 ( .A(G132), .ZN(G219) );
  INV_X1 U858 ( .A(G82), .ZN(G220) );
  INV_X1 U859 ( .A(G57), .ZN(G237) );
  INV_X1 U860 ( .A(G120), .ZN(G236) );
  NAND2_X1 U861 ( .A1(G94), .A2(G452), .ZN(n785) );
  XNOR2_X1 U862 ( .A(n785), .B(KEYINPUT67), .ZN(G173) );
  XOR2_X1 U863 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n787) );
  NAND2_X1 U864 ( .A1(G7), .A2(G661), .ZN(n786) );
  XNOR2_X1 U865 ( .A(n787), .B(n786), .ZN(G223) );
  INV_X1 U866 ( .A(G223), .ZN(n846) );
  NAND2_X1 U867 ( .A1(n846), .A2(G567), .ZN(n788) );
  XOR2_X1 U868 ( .A(KEYINPUT11), .B(n788), .Z(G234) );
  INV_X1 U869 ( .A(G860), .ZN(n794) );
  OR2_X1 U870 ( .A1(n934), .A2(n794), .ZN(G153) );
  NOR2_X1 U871 ( .A1(n927), .A2(G868), .ZN(n789) );
  XOR2_X1 U872 ( .A(KEYINPUT70), .B(n789), .Z(n791) );
  NAND2_X1 U873 ( .A1(G868), .A2(G301), .ZN(n790) );
  NAND2_X1 U874 ( .A1(n791), .A2(n790), .ZN(G284) );
  INV_X1 U875 ( .A(G868), .ZN(n824) );
  NOR2_X1 U876 ( .A1(G286), .A2(n824), .ZN(n793) );
  NOR2_X1 U877 ( .A1(G868), .A2(G299), .ZN(n792) );
  NOR2_X1 U878 ( .A1(n793), .A2(n792), .ZN(G297) );
  NAND2_X1 U879 ( .A1(n794), .A2(G559), .ZN(n795) );
  NAND2_X1 U880 ( .A1(n795), .A2(n927), .ZN(n796) );
  XNOR2_X1 U881 ( .A(n796), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U882 ( .A1(G868), .A2(n934), .ZN(n797) );
  XNOR2_X1 U883 ( .A(KEYINPUT74), .B(n797), .ZN(n800) );
  NAND2_X1 U884 ( .A1(G868), .A2(n927), .ZN(n798) );
  NOR2_X1 U885 ( .A1(G559), .A2(n798), .ZN(n799) );
  NOR2_X1 U886 ( .A1(n800), .A2(n799), .ZN(G282) );
  NAND2_X1 U887 ( .A1(n927), .A2(G559), .ZN(n822) );
  XNOR2_X1 U888 ( .A(n934), .B(n822), .ZN(n801) );
  NOR2_X1 U889 ( .A1(n801), .A2(G860), .ZN(n813) );
  NAND2_X1 U890 ( .A1(G93), .A2(n802), .ZN(n805) );
  NAND2_X1 U891 ( .A1(G80), .A2(n803), .ZN(n804) );
  NAND2_X1 U892 ( .A1(n805), .A2(n804), .ZN(n812) );
  NAND2_X1 U893 ( .A1(G55), .A2(n806), .ZN(n807) );
  XNOR2_X1 U894 ( .A(n807), .B(KEYINPUT76), .ZN(n810) );
  NAND2_X1 U895 ( .A1(n808), .A2(G67), .ZN(n809) );
  NAND2_X1 U896 ( .A1(n810), .A2(n809), .ZN(n811) );
  OR2_X1 U897 ( .A1(n812), .A2(n811), .ZN(n825) );
  XOR2_X1 U898 ( .A(n813), .B(n825), .Z(G145) );
  XNOR2_X1 U899 ( .A(KEYINPUT19), .B(KEYINPUT81), .ZN(n815) );
  XNOR2_X1 U900 ( .A(G288), .B(KEYINPUT80), .ZN(n814) );
  XNOR2_X1 U901 ( .A(n815), .B(n814), .ZN(n818) );
  XOR2_X1 U902 ( .A(n825), .B(G290), .Z(n816) );
  XNOR2_X1 U903 ( .A(n816), .B(n934), .ZN(n817) );
  XNOR2_X1 U904 ( .A(n818), .B(n817), .ZN(n820) );
  XNOR2_X1 U905 ( .A(G299), .B(G166), .ZN(n819) );
  XNOR2_X1 U906 ( .A(n820), .B(n819), .ZN(n821) );
  XNOR2_X1 U907 ( .A(n821), .B(G305), .ZN(n911) );
  XNOR2_X1 U908 ( .A(n911), .B(n822), .ZN(n823) );
  NOR2_X1 U909 ( .A1(n824), .A2(n823), .ZN(n827) );
  NOR2_X1 U910 ( .A1(G868), .A2(n825), .ZN(n826) );
  NOR2_X1 U911 ( .A1(n827), .A2(n826), .ZN(G295) );
  NAND2_X1 U912 ( .A1(G2084), .A2(G2078), .ZN(n828) );
  XOR2_X1 U913 ( .A(KEYINPUT20), .B(n828), .Z(n829) );
  NAND2_X1 U914 ( .A1(n829), .A2(G2090), .ZN(n830) );
  XNOR2_X1 U915 ( .A(n830), .B(KEYINPUT21), .ZN(n831) );
  XNOR2_X1 U916 ( .A(KEYINPUT82), .B(n831), .ZN(n832) );
  NAND2_X1 U917 ( .A1(G2072), .A2(n832), .ZN(G158) );
  NOR2_X1 U918 ( .A1(G236), .A2(G237), .ZN(n833) );
  NAND2_X1 U919 ( .A1(G69), .A2(n833), .ZN(n834) );
  XNOR2_X1 U920 ( .A(KEYINPUT83), .B(n834), .ZN(n835) );
  NAND2_X1 U921 ( .A1(n835), .A2(G108), .ZN(n836) );
  XNOR2_X1 U922 ( .A(KEYINPUT84), .B(n836), .ZN(n850) );
  NAND2_X1 U923 ( .A1(n850), .A2(G567), .ZN(n837) );
  XNOR2_X1 U924 ( .A(n837), .B(KEYINPUT85), .ZN(n842) );
  NOR2_X1 U925 ( .A1(G220), .A2(G219), .ZN(n838) );
  XNOR2_X1 U926 ( .A(KEYINPUT22), .B(n838), .ZN(n839) );
  NAND2_X1 U927 ( .A1(n839), .A2(G96), .ZN(n840) );
  OR2_X1 U928 ( .A1(G218), .A2(n840), .ZN(n851) );
  AND2_X1 U929 ( .A1(G2106), .A2(n851), .ZN(n841) );
  NOR2_X1 U930 ( .A1(n842), .A2(n841), .ZN(G319) );
  INV_X1 U931 ( .A(G319), .ZN(n844) );
  NAND2_X1 U932 ( .A1(G483), .A2(G661), .ZN(n843) );
  NOR2_X1 U933 ( .A1(n844), .A2(n843), .ZN(n849) );
  NAND2_X1 U934 ( .A1(n849), .A2(G36), .ZN(n845) );
  XNOR2_X1 U935 ( .A(KEYINPUT86), .B(n845), .ZN(G176) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n846), .ZN(G217) );
  AND2_X1 U937 ( .A1(G15), .A2(G2), .ZN(n847) );
  NAND2_X1 U938 ( .A1(G661), .A2(n847), .ZN(G259) );
  NAND2_X1 U939 ( .A1(G3), .A2(G1), .ZN(n848) );
  NAND2_X1 U940 ( .A1(n849), .A2(n848), .ZN(G188) );
  INV_X1 U942 ( .A(G108), .ZN(G238) );
  INV_X1 U943 ( .A(G96), .ZN(G221) );
  NOR2_X1 U944 ( .A1(n851), .A2(n850), .ZN(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  XOR2_X1 U946 ( .A(KEYINPUT42), .B(G2072), .Z(n853) );
  XNOR2_X1 U947 ( .A(G2084), .B(G2078), .ZN(n852) );
  XNOR2_X1 U948 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U949 ( .A(n854), .B(G2100), .Z(n856) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2090), .ZN(n855) );
  XNOR2_X1 U951 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U952 ( .A(G2096), .B(KEYINPUT43), .Z(n858) );
  XNOR2_X1 U953 ( .A(KEYINPUT109), .B(G2678), .ZN(n857) );
  XNOR2_X1 U954 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U955 ( .A(n860), .B(n859), .Z(G227) );
  XNOR2_X1 U956 ( .A(G1956), .B(KEYINPUT41), .ZN(n870) );
  XOR2_X1 U957 ( .A(G1976), .B(G1971), .Z(n862) );
  XNOR2_X1 U958 ( .A(G1981), .B(G1961), .ZN(n861) );
  XNOR2_X1 U959 ( .A(n862), .B(n861), .ZN(n866) );
  XOR2_X1 U960 ( .A(G1966), .B(G1986), .Z(n864) );
  XNOR2_X1 U961 ( .A(G1996), .B(G1991), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U963 ( .A(n866), .B(n865), .Z(n868) );
  XNOR2_X1 U964 ( .A(KEYINPUT110), .B(G2474), .ZN(n867) );
  XNOR2_X1 U965 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U966 ( .A(n870), .B(n869), .ZN(G229) );
  NAND2_X1 U967 ( .A1(G124), .A2(n898), .ZN(n871) );
  XNOR2_X1 U968 ( .A(n871), .B(KEYINPUT44), .ZN(n874) );
  NAND2_X1 U969 ( .A1(G112), .A2(n515), .ZN(n872) );
  XOR2_X1 U970 ( .A(KEYINPUT111), .B(n872), .Z(n873) );
  NAND2_X1 U971 ( .A1(n874), .A2(n873), .ZN(n878) );
  NAND2_X1 U972 ( .A1(G100), .A2(n895), .ZN(n876) );
  NAND2_X1 U973 ( .A1(G136), .A2(n717), .ZN(n875) );
  NAND2_X1 U974 ( .A1(n876), .A2(n875), .ZN(n877) );
  NOR2_X1 U975 ( .A1(n878), .A2(n877), .ZN(G162) );
  NAND2_X1 U976 ( .A1(G106), .A2(n895), .ZN(n880) );
  NAND2_X1 U977 ( .A1(G142), .A2(n717), .ZN(n879) );
  NAND2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U979 ( .A(n881), .B(KEYINPUT45), .ZN(n883) );
  NAND2_X1 U980 ( .A1(G130), .A2(n898), .ZN(n882) );
  NAND2_X1 U981 ( .A1(n883), .A2(n882), .ZN(n886) );
  NAND2_X1 U982 ( .A1(n515), .A2(G118), .ZN(n884) );
  XOR2_X1 U983 ( .A(KEYINPUT112), .B(n884), .Z(n885) );
  NOR2_X1 U984 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U985 ( .A(G160), .B(n887), .ZN(n907) );
  XNOR2_X1 U986 ( .A(G162), .B(n888), .ZN(n889) );
  XNOR2_X1 U987 ( .A(n889), .B(n998), .ZN(n894) );
  XNOR2_X1 U988 ( .A(KEYINPUT48), .B(KEYINPUT113), .ZN(n892) );
  XNOR2_X1 U989 ( .A(n890), .B(KEYINPUT46), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U991 ( .A(n894), .B(n893), .Z(n905) );
  NAND2_X1 U992 ( .A1(G103), .A2(n895), .ZN(n897) );
  NAND2_X1 U993 ( .A1(G139), .A2(n717), .ZN(n896) );
  NAND2_X1 U994 ( .A1(n897), .A2(n896), .ZN(n903) );
  NAND2_X1 U995 ( .A1(G127), .A2(n898), .ZN(n900) );
  NAND2_X1 U996 ( .A1(G115), .A2(n515), .ZN(n899) );
  NAND2_X1 U997 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U998 ( .A(KEYINPUT47), .B(n901), .Z(n902) );
  NOR2_X1 U999 ( .A1(n903), .A2(n902), .ZN(n1011) );
  XNOR2_X1 U1000 ( .A(G164), .B(n1011), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n909) );
  XOR2_X1 U1003 ( .A(n909), .B(n908), .Z(n910) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n910), .ZN(G395) );
  XOR2_X1 U1005 ( .A(KEYINPUT114), .B(n911), .Z(n913) );
  XNOR2_X1 U1006 ( .A(n927), .B(G286), .ZN(n912) );
  XNOR2_X1 U1007 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1008 ( .A(n914), .B(G171), .ZN(n915) );
  NOR2_X1 U1009 ( .A1(G37), .A2(n915), .ZN(G397) );
  NOR2_X1 U1010 ( .A1(G227), .A2(G229), .ZN(n916) );
  XOR2_X1 U1011 ( .A(KEYINPUT49), .B(n916), .Z(n917) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n917), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(G401), .A2(n918), .ZN(n921) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n919) );
  XOR2_X1 U1015 ( .A(KEYINPUT115), .B(n919), .Z(n920) );
  NAND2_X1 U1016 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1019 ( .A(G1966), .B(G168), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1021 ( .A(KEYINPUT57), .B(n924), .Z(n943) );
  NAND2_X1 U1022 ( .A1(G1971), .A2(G303), .ZN(n925) );
  NAND2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n940) );
  XOR2_X1 U1024 ( .A(G1348), .B(n927), .Z(n929) );
  XOR2_X1 U1025 ( .A(G171), .B(G1961), .Z(n928) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n938) );
  XNOR2_X1 U1027 ( .A(G1956), .B(G299), .ZN(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n933) );
  NAND2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n936) );
  XNOR2_X1 U1030 ( .A(G1341), .B(n934), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(n941), .B(KEYINPUT123), .ZN(n942) );
  NOR2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1036 ( .A(KEYINPUT124), .B(n944), .Z(n946) );
  XNOR2_X1 U1037 ( .A(G16), .B(KEYINPUT56), .ZN(n945) );
  NAND2_X1 U1038 ( .A1(n946), .A2(n945), .ZN(n1026) );
  XNOR2_X1 U1039 ( .A(G5), .B(G1961), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(n947), .B(KEYINPUT125), .ZN(n966) );
  XNOR2_X1 U1041 ( .A(G1986), .B(G24), .ZN(n952) );
  XNOR2_X1 U1042 ( .A(G1971), .B(G22), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(G1976), .B(G23), .ZN(n948) );
  NOR2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(KEYINPUT127), .B(n950), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1047 ( .A(KEYINPUT58), .B(n953), .Z(n964) );
  XOR2_X1 U1048 ( .A(G1348), .B(KEYINPUT59), .Z(n954) );
  XNOR2_X1 U1049 ( .A(G4), .B(n954), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(G6), .B(G1981), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n960) );
  XNOR2_X1 U1052 ( .A(G1956), .B(G20), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(G1341), .B(G19), .ZN(n957) );
  NOR2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(n961), .B(KEYINPUT126), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(KEYINPUT60), .B(n962), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(G21), .B(G1966), .ZN(n967) );
  NOR2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(KEYINPUT61), .B(n969), .ZN(n971) );
  INV_X1 U1063 ( .A(G16), .ZN(n970) );
  NAND2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(n972), .A2(G11), .ZN(n1024) );
  XNOR2_X1 U1066 ( .A(G35), .B(G2090), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(n973), .B(KEYINPUT119), .ZN(n988) );
  XNOR2_X1 U1068 ( .A(KEYINPUT53), .B(KEYINPUT121), .ZN(n986) );
  XNOR2_X1 U1069 ( .A(G2067), .B(G26), .ZN(n975) );
  XNOR2_X1 U1070 ( .A(G2072), .B(G33), .ZN(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1072 ( .A(KEYINPUT120), .B(n976), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(G1996), .B(G32), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(n977), .B(G27), .ZN(n978) );
  NOR2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n984) );
  XOR2_X1 U1077 ( .A(G1991), .B(G25), .Z(n982) );
  NAND2_X1 U1078 ( .A1(G28), .A2(n982), .ZN(n983) );
  NOR2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(n986), .B(n985), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(KEYINPUT122), .B(n989), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(G34), .B(G2084), .ZN(n990) );
  XNOR2_X1 U1084 ( .A(KEYINPUT54), .B(n990), .ZN(n991) );
  NOR2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1086 ( .A1(G29), .A2(n993), .ZN(n994) );
  XNOR2_X1 U1087 ( .A(n994), .B(KEYINPUT55), .ZN(n1022) );
  XNOR2_X1 U1088 ( .A(G2084), .B(G160), .ZN(n995) );
  XNOR2_X1 U1089 ( .A(n995), .B(KEYINPUT116), .ZN(n1007) );
  NOR2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1005) );
  XOR2_X1 U1092 ( .A(G2090), .B(G162), .Z(n1000) );
  NOR2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1094 ( .A(KEYINPUT117), .B(n1002), .Z(n1003) );
  XNOR2_X1 U1095 ( .A(n1003), .B(KEYINPUT51), .ZN(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1099 ( .A(KEYINPUT118), .B(n1010), .Z(n1016) );
  XOR2_X1 U1100 ( .A(G2072), .B(n1011), .Z(n1013) );
  XOR2_X1 U1101 ( .A(G164), .B(G2078), .Z(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1103 ( .A(KEYINPUT50), .B(n1014), .Z(n1015) );
  NOR2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1018) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(KEYINPUT52), .B(n1019), .ZN(n1020) );
  NAND2_X1 U1107 ( .A1(G29), .A2(n1020), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1027), .Z(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

