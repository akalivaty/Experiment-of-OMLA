

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783;

  AND2_X1 U384 ( .A1(n364), .A2(n622), .ZN(n633) );
  XNOR2_X1 U385 ( .A(n519), .B(n462), .ZN(n461) );
  INV_X1 U386 ( .A(G953), .ZN(n709) );
  OR2_X2 U387 ( .A1(n644), .A2(n707), .ZN(n638) );
  XNOR2_X2 U388 ( .A(n686), .B(KEYINPUT109), .ZN(n622) );
  XNOR2_X2 U389 ( .A(n552), .B(n551), .ZN(n653) );
  XNOR2_X2 U390 ( .A(n456), .B(n763), .ZN(n740) );
  NOR2_X1 U391 ( .A1(n606), .A2(n605), .ZN(n730) );
  NOR2_X1 U392 ( .A1(n780), .A2(n779), .ZN(n431) );
  OR2_X1 U393 ( .A1(n600), .A2(n486), .ZN(n485) );
  XNOR2_X1 U394 ( .A(n457), .B(KEYINPUT22), .ZN(n600) );
  XNOR2_X1 U395 ( .A(n634), .B(n443), .ZN(n683) );
  XNOR2_X1 U396 ( .A(G104), .B(G110), .ZN(n438) );
  NAND2_X1 U397 ( .A1(n401), .A2(n400), .ZN(n433) );
  AND2_X1 U398 ( .A1(n403), .A2(n402), .ZN(n401) );
  AND2_X1 U399 ( .A1(G475), .A2(n746), .ZN(n747) );
  NOR2_X1 U400 ( .A1(n389), .A2(n385), .ZN(n711) );
  NAND2_X1 U401 ( .A1(n361), .A2(n369), .ZN(n407) );
  NAND2_X1 U402 ( .A1(n431), .A2(n781), .ZN(n453) );
  XNOR2_X1 U403 ( .A(n599), .B(KEYINPUT111), .ZN(n780) );
  XNOR2_X1 U404 ( .A(n594), .B(n593), .ZN(n779) );
  XNOR2_X1 U405 ( .A(n485), .B(KEYINPUT83), .ZN(n602) );
  NOR2_X1 U406 ( .A1(n610), .A2(n696), .ZN(n613) );
  NOR2_X1 U407 ( .A1(n678), .A2(n677), .ZN(n637) );
  NOR2_X1 U408 ( .A1(n461), .A2(n524), .ZN(n526) );
  XNOR2_X1 U409 ( .A(n596), .B(n445), .ZN(n677) );
  INV_X1 U410 ( .A(n653), .ZN(n688) );
  XNOR2_X1 U411 ( .A(n664), .B(KEYINPUT38), .ZN(n675) );
  XNOR2_X1 U412 ( .A(n536), .B(KEYINPUT10), .ZN(n770) );
  INV_X1 U413 ( .A(n438), .ZN(n514) );
  XNOR2_X1 U414 ( .A(KEYINPUT91), .B(KEYINPUT77), .ZN(n513) );
  NOR2_X2 U415 ( .A1(n753), .A2(n372), .ZN(n426) );
  NOR2_X2 U416 ( .A1(G902), .A2(n742), .ZN(n535) );
  OR2_X1 U417 ( .A1(n740), .A2(n384), .ZN(n383) );
  INV_X1 U418 ( .A(KEYINPUT78), .ZN(n390) );
  XNOR2_X1 U419 ( .A(n584), .B(n482), .ZN(n533) );
  XNOR2_X1 U420 ( .A(KEYINPUT4), .B(KEYINPUT68), .ZN(n482) );
  XNOR2_X1 U421 ( .A(G146), .B(n769), .ZN(n560) );
  INV_X1 U422 ( .A(KEYINPUT1), .ZN(n443) );
  NOR2_X1 U423 ( .A1(n382), .A2(n381), .ZN(n380) );
  INV_X1 U424 ( .A(n674), .ZN(n381) );
  XNOR2_X1 U425 ( .A(n770), .B(n568), .ZN(n575) );
  XNOR2_X1 U426 ( .A(G113), .B(G131), .ZN(n572) );
  XNOR2_X1 U427 ( .A(n591), .B(n590), .ZN(n606) );
  INV_X1 U428 ( .A(KEYINPUT47), .ZN(n450) );
  NOR2_X1 U429 ( .A1(n645), .A2(n614), .ZN(n615) );
  NOR2_X1 U430 ( .A1(n738), .A2(n390), .ZN(n387) );
  NAND2_X1 U431 ( .A1(n670), .A2(n366), .ZN(n388) );
  XNOR2_X1 U432 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n478) );
  NOR2_X1 U433 ( .A1(n496), .A2(n488), .ZN(n487) );
  INV_X1 U434 ( .A(KEYINPUT44), .ZN(n488) );
  NOR2_X1 U435 ( .A1(G953), .A2(G237), .ZN(n569) );
  XOR2_X1 U436 ( .A(KEYINPUT76), .B(KEYINPUT5), .Z(n557) );
  XNOR2_X1 U437 ( .A(n533), .B(n479), .ZN(n769) );
  XNOR2_X1 U438 ( .A(n481), .B(n480), .ZN(n479) );
  XNOR2_X1 U439 ( .A(KEYINPUT70), .B(G131), .ZN(n481) );
  XNOR2_X1 U440 ( .A(G137), .B(G134), .ZN(n480) );
  XNOR2_X1 U441 ( .A(G146), .B(G125), .ZN(n467) );
  XNOR2_X1 U442 ( .A(KEYINPUT69), .B(KEYINPUT87), .ZN(n538) );
  INV_X1 U443 ( .A(n708), .ZN(n501) );
  INV_X1 U444 ( .A(KEYINPUT93), .ZN(n515) );
  INV_X1 U445 ( .A(n631), .ZN(n477) );
  NAND2_X1 U446 ( .A1(n437), .A2(n714), .ZN(n398) );
  XNOR2_X1 U447 ( .A(n713), .B(KEYINPUT66), .ZN(n714) );
  NAND2_X1 U448 ( .A1(n757), .A2(n711), .ZN(n437) );
  XNOR2_X1 U449 ( .A(n512), .B(n395), .ZN(n394) );
  OR2_X2 U450 ( .A1(n710), .A2(n669), .ZN(n746) );
  XNOR2_X1 U451 ( .A(n439), .B(KEYINPUT88), .ZN(n672) );
  NOR2_X1 U452 ( .A1(n653), .A2(n652), .ZN(n661) );
  NAND2_X1 U453 ( .A1(n460), .A2(n458), .ZN(n457) );
  NOR2_X1 U454 ( .A1(n677), .A2(n459), .ZN(n458) );
  INV_X1 U455 ( .A(n664), .ZN(n391) );
  XOR2_X1 U456 ( .A(n579), .B(n578), .Z(n605) );
  NOR2_X1 U457 ( .A1(n748), .A2(G902), .ZN(n579) );
  NAND2_X2 U458 ( .A1(n471), .A2(n468), .ZN(n686) );
  AND2_X1 U459 ( .A1(n473), .A2(n472), .ZN(n471) );
  NAND2_X1 U460 ( .A1(G472), .A2(n470), .ZN(n469) );
  BUF_X1 U461 ( .A(n597), .Z(n610) );
  NOR2_X1 U462 ( .A1(n372), .A2(G472), .ZN(n464) );
  XNOR2_X1 U463 ( .A(n441), .B(n587), .ZN(n751) );
  XNOR2_X1 U464 ( .A(n589), .B(n588), .ZN(n441) );
  AND2_X2 U465 ( .A1(n398), .A2(n746), .ZN(n753) );
  NAND2_X1 U466 ( .A1(n727), .A2(n643), .ZN(n440) );
  XNOR2_X1 U467 ( .A(G113), .B(G101), .ZN(n508) );
  NAND2_X1 U468 ( .A1(n495), .A2(KEYINPUT90), .ZN(n494) );
  INV_X1 U469 ( .A(KEYINPUT75), .ZN(n452) );
  OR2_X1 U470 ( .A1(G237), .A2(G902), .ZN(n518) );
  NAND2_X1 U471 ( .A1(n454), .A2(n547), .ZN(n384) );
  NOR2_X1 U472 ( .A1(n454), .A2(n547), .ZN(n382) );
  XNOR2_X1 U473 ( .A(G143), .B(G122), .ZN(n566) );
  XOR2_X1 U474 ( .A(KEYINPUT99), .B(G104), .Z(n567) );
  XNOR2_X1 U475 ( .A(n446), .B(n571), .ZN(n573) );
  XNOR2_X1 U476 ( .A(n570), .B(n447), .ZN(n446) );
  INV_X1 U477 ( .A(KEYINPUT11), .ZN(n447) );
  XOR2_X1 U478 ( .A(G101), .B(G107), .Z(n528) );
  NAND2_X1 U479 ( .A1(n388), .A2(n386), .ZN(n385) );
  NOR2_X1 U480 ( .A1(n387), .A2(n547), .ZN(n386) );
  INV_X1 U481 ( .A(KEYINPUT72), .ZN(n499) );
  XNOR2_X1 U482 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n395) );
  XNOR2_X1 U483 ( .A(n467), .B(KEYINPUT80), .ZN(n397) );
  NAND2_X1 U484 ( .A1(n675), .A2(n674), .ZN(n678) );
  INV_X1 U485 ( .A(n598), .ZN(n459) );
  INV_X1 U486 ( .A(KEYINPUT108), .ZN(n445) );
  NAND2_X1 U487 ( .A1(n430), .A2(n429), .ZN(n696) );
  INV_X1 U488 ( .A(n609), .ZN(n430) );
  INV_X1 U489 ( .A(G902), .ZN(n470) );
  NAND2_X1 U490 ( .A1(n474), .A2(G902), .ZN(n472) );
  XNOR2_X1 U491 ( .A(n560), .B(n561), .ZN(n715) );
  XNOR2_X1 U492 ( .A(n558), .B(n559), .ZN(n451) );
  BUF_X1 U493 ( .A(n683), .Z(n448) );
  XNOR2_X1 U494 ( .A(n467), .B(n466), .ZN(n536) );
  INV_X1 U495 ( .A(G140), .ZN(n466) );
  XNOR2_X1 U496 ( .A(n538), .B(n537), .ZN(n539) );
  INV_X1 U497 ( .A(KEYINPUT8), .ZN(n537) );
  XNOR2_X1 U498 ( .A(G134), .B(KEYINPUT104), .ZN(n580) );
  XOR2_X1 U499 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n581) );
  OR2_X1 U500 ( .A1(n500), .A2(KEYINPUT121), .ZN(n410) );
  INV_X1 U501 ( .A(KEYINPUT19), .ZN(n462) );
  NAND2_X1 U502 ( .A1(n368), .A2(n379), .ZN(n519) );
  AND2_X1 U503 ( .A1(n626), .A2(n476), .ZN(n641) );
  NOR2_X1 U504 ( .A1(n634), .A2(n607), .ZN(n625) );
  NOR2_X1 U505 ( .A1(n425), .A2(KEYINPUT63), .ZN(n422) );
  XNOR2_X1 U506 ( .A(n418), .B(n374), .ZN(n417) );
  NAND2_X1 U507 ( .A1(n747), .A2(n398), .ZN(n418) );
  INV_X1 U508 ( .A(KEYINPUT121), .ZN(n409) );
  INV_X1 U509 ( .A(KEYINPUT40), .ZN(n629) );
  NOR2_X1 U510 ( .A1(n662), .A2(n656), .ZN(n735) );
  XOR2_X1 U511 ( .A(KEYINPUT32), .B(n602), .Z(n781) );
  NAND2_X1 U512 ( .A1(n601), .A2(n363), .ZN(n486) );
  NAND2_X1 U513 ( .A1(n642), .A2(n391), .ZN(n727) );
  AND2_X1 U514 ( .A1(n641), .A2(n640), .ZN(n642) );
  AND2_X1 U515 ( .A1(n606), .A2(n605), .ZN(n732) );
  XNOR2_X1 U516 ( .A(n484), .B(n483), .ZN(n752) );
  XNOR2_X1 U517 ( .A(n751), .B(n750), .ZN(n483) );
  XNOR2_X1 U518 ( .A(n434), .B(n373), .ZN(n745) );
  INV_X1 U519 ( .A(KEYINPUT56), .ZN(n419) );
  AND2_X1 U520 ( .A1(n410), .A2(n709), .ZN(n361) );
  INV_X1 U521 ( .A(G472), .ZN(n474) );
  AND2_X1 U522 ( .A1(n670), .A2(n738), .ZN(n362) );
  XNOR2_X1 U523 ( .A(n562), .B(n686), .ZN(n363) );
  AND2_X1 U524 ( .A1(n688), .A2(n649), .ZN(n364) );
  AND2_X1 U525 ( .A1(n672), .A2(n409), .ZN(n365) );
  AND2_X1 U526 ( .A1(n738), .A2(n390), .ZN(n366) );
  AND2_X1 U527 ( .A1(n746), .A2(G210), .ZN(n367) );
  INV_X1 U528 ( .A(n686), .ZN(n429) );
  AND2_X1 U529 ( .A1(n383), .A2(n380), .ZN(n368) );
  NAND2_X1 U530 ( .A1(n500), .A2(KEYINPUT121), .ZN(n369) );
  XOR2_X1 U531 ( .A(n435), .B(KEYINPUT74), .Z(n370) );
  OR2_X1 U532 ( .A1(KEYINPUT2), .A2(n362), .ZN(n371) );
  XOR2_X1 U533 ( .A(n715), .B(KEYINPUT62), .Z(n372) );
  INV_X1 U534 ( .A(n756), .ZN(n465) );
  XOR2_X1 U535 ( .A(n744), .B(n743), .Z(n373) );
  XNOR2_X1 U536 ( .A(KEYINPUT15), .B(G902), .ZN(n547) );
  XOR2_X1 U537 ( .A(n748), .B(n504), .Z(n374) );
  XOR2_X1 U538 ( .A(n740), .B(n741), .Z(n375) );
  XOR2_X1 U539 ( .A(n660), .B(KEYINPUT48), .Z(n376) );
  AND2_X1 U540 ( .A1(n372), .A2(G472), .ZN(n377) );
  INV_X1 U541 ( .A(n463), .ZN(n425) );
  NOR2_X1 U542 ( .A1(n464), .A2(n756), .ZN(n463) );
  XOR2_X1 U543 ( .A(n749), .B(KEYINPUT60), .Z(n378) );
  OR2_X1 U544 ( .A1(n740), .A2(n712), .ZN(n455) );
  NAND2_X1 U545 ( .A1(n740), .A2(n517), .ZN(n379) );
  NOR2_X1 U546 ( .A1(n670), .A2(n390), .ZN(n389) );
  XNOR2_X2 U547 ( .A(n667), .B(KEYINPUT89), .ZN(n670) );
  NAND2_X1 U548 ( .A1(n661), .A2(n391), .ZN(n654) );
  XNOR2_X2 U549 ( .A(n455), .B(n517), .ZN(n664) );
  NAND2_X1 U550 ( .A1(n653), .A2(n598), .ZN(n607) );
  XNOR2_X1 U551 ( .A(n754), .B(n755), .ZN(n404) );
  AND2_X1 U552 ( .A1(n746), .A2(n371), .ZN(n673) );
  XNOR2_X1 U553 ( .A(G119), .B(G128), .ZN(n541) );
  XNOR2_X1 U554 ( .A(n533), .B(n397), .ZN(n396) );
  XNOR2_X1 U555 ( .A(n527), .B(n393), .ZN(n456) );
  XNOR2_X1 U556 ( .A(n396), .B(n394), .ZN(n393) );
  XNOR2_X1 U557 ( .A(n421), .B(n375), .ZN(n420) );
  XNOR2_X1 U558 ( .A(n451), .B(n392), .ZN(n561) );
  XNOR2_X2 U559 ( .A(n392), .B(KEYINPUT73), .ZN(n498) );
  XNOR2_X2 U560 ( .A(n510), .B(n509), .ZN(n392) );
  XNOR2_X2 U561 ( .A(n762), .B(n499), .ZN(n527) );
  XNOR2_X2 U562 ( .A(n514), .B(n513), .ZN(n762) );
  NAND2_X1 U563 ( .A1(n367), .A2(n398), .ZN(n421) );
  INV_X1 U564 ( .A(n673), .ZN(n399) );
  NAND2_X1 U565 ( .A1(n408), .A2(n407), .ZN(n403) );
  NAND2_X1 U566 ( .A1(n399), .A2(n407), .ZN(n402) );
  NAND2_X1 U567 ( .A1(n365), .A2(n673), .ZN(n400) );
  NOR2_X1 U568 ( .A1(n404), .A2(n756), .ZN(G66) );
  XNOR2_X1 U569 ( .A(n405), .B(n419), .ZN(G51) );
  NAND2_X1 U570 ( .A1(n420), .A2(n465), .ZN(n405) );
  NAND2_X1 U571 ( .A1(n492), .A2(n491), .ZN(n490) );
  XNOR2_X1 U572 ( .A(n406), .B(n378), .ZN(G60) );
  NAND2_X1 U573 ( .A1(n417), .A2(n465), .ZN(n406) );
  NAND2_X1 U574 ( .A1(n672), .A2(n361), .ZN(n408) );
  NAND2_X1 U575 ( .A1(n411), .A2(n416), .ZN(n415) );
  NAND2_X1 U576 ( .A1(n413), .A2(n412), .ZN(n411) );
  NAND2_X1 U577 ( .A1(n424), .A2(n422), .ZN(n412) );
  INV_X1 U578 ( .A(n426), .ZN(n413) );
  NAND2_X1 U579 ( .A1(n426), .A2(n716), .ZN(n416) );
  NAND2_X1 U580 ( .A1(n415), .A2(n414), .ZN(G57) );
  NAND2_X1 U581 ( .A1(n423), .A2(KEYINPUT63), .ZN(n414) );
  NAND2_X1 U582 ( .A1(n424), .A2(n463), .ZN(n423) );
  NAND2_X1 U583 ( .A1(n753), .A2(n377), .ZN(n424) );
  NAND2_X1 U584 ( .A1(n427), .A2(n494), .ZN(n493) );
  NAND2_X1 U585 ( .A1(n497), .A2(n489), .ZN(n427) );
  BUF_X1 U586 ( .A(n742), .Z(n428) );
  XNOR2_X2 U587 ( .A(n556), .B(n452), .ZN(n609) );
  XNOR2_X1 U588 ( .A(n433), .B(n432), .ZN(G75) );
  INV_X1 U589 ( .A(KEYINPUT53), .ZN(n432) );
  NAND2_X1 U590 ( .A1(n753), .A2(G469), .ZN(n434) );
  NAND2_X1 U591 ( .A1(n648), .A2(n647), .ZN(n435) );
  XNOR2_X1 U592 ( .A(n436), .B(n376), .ZN(n666) );
  NAND2_X1 U593 ( .A1(n658), .A2(n659), .ZN(n436) );
  XNOR2_X1 U594 ( .A(n444), .B(n478), .ZN(n659) );
  NAND2_X1 U595 ( .A1(n622), .A2(n674), .ZN(n624) );
  NAND2_X1 U596 ( .A1(n715), .A2(n474), .ZN(n473) );
  NAND2_X1 U597 ( .A1(n710), .A2(n671), .ZN(n439) );
  XNOR2_X1 U598 ( .A(n440), .B(KEYINPUT85), .ZN(n648) );
  AND2_X1 U599 ( .A1(n625), .A2(n477), .ZN(n476) );
  XNOR2_X1 U600 ( .A(n563), .B(KEYINPUT33), .ZN(n706) );
  NOR2_X1 U601 ( .A1(n706), .A2(n610), .ZN(n565) );
  XNOR2_X2 U602 ( .A(n639), .B(n638), .ZN(n778) );
  NAND2_X1 U603 ( .A1(n683), .A2(n684), .ZN(n556) );
  NAND2_X1 U604 ( .A1(n442), .A2(n502), .ZN(n599) );
  XNOR2_X1 U605 ( .A(n603), .B(KEYINPUT110), .ZN(n442) );
  INV_X1 U606 ( .A(n683), .ZN(n662) );
  XNOR2_X1 U607 ( .A(n574), .B(n575), .ZN(n748) );
  NOR2_X2 U608 ( .A1(n778), .A2(n782), .ZN(n444) );
  NAND2_X1 U609 ( .A1(n646), .A2(n449), .ZN(n647) );
  XNOR2_X1 U610 ( .A(n728), .B(n450), .ZN(n449) );
  INV_X1 U611 ( .A(n622), .ZN(n632) );
  XNOR2_X2 U612 ( .A(n535), .B(G469), .ZN(n634) );
  XNOR2_X1 U613 ( .A(n613), .B(n612), .ZN(n733) );
  NAND2_X1 U614 ( .A1(n453), .A2(KEYINPUT44), .ZN(n497) );
  NOR2_X1 U615 ( .A1(n453), .A2(KEYINPUT44), .ZN(n618) );
  NAND2_X1 U616 ( .A1(n453), .A2(n487), .ZN(n491) );
  INV_X1 U617 ( .A(n517), .ZN(n454) );
  NOR2_X2 U618 ( .A1(n600), .A2(n448), .ZN(n603) );
  INV_X1 U619 ( .A(n597), .ZN(n460) );
  NOR2_X2 U620 ( .A1(n644), .A2(n461), .ZN(n728) );
  OR2_X1 U621 ( .A1(n715), .A2(n469), .ZN(n468) );
  XNOR2_X1 U622 ( .A(n475), .B(KEYINPUT39), .ZN(n628) );
  NAND2_X1 U623 ( .A1(n641), .A2(n675), .ZN(n475) );
  XNOR2_X2 U624 ( .A(G143), .B(G128), .ZN(n584) );
  NAND2_X1 U625 ( .A1(n753), .A2(G478), .ZN(n484) );
  INV_X1 U626 ( .A(n618), .ZN(n492) );
  AND2_X1 U627 ( .A1(n617), .A2(n496), .ZN(n489) );
  NOR2_X2 U628 ( .A1(n493), .A2(n490), .ZN(n619) );
  INV_X1 U629 ( .A(n617), .ZN(n495) );
  INV_X1 U630 ( .A(KEYINPUT90), .ZN(n496) );
  XNOR2_X2 U631 ( .A(n511), .B(n498), .ZN(n763) );
  NOR2_X1 U632 ( .A1(n705), .A2(n501), .ZN(n500) );
  AND2_X1 U633 ( .A1(n632), .A2(n688), .ZN(n502) );
  AND2_X1 U634 ( .A1(n586), .A2(G221), .ZN(n503) );
  XNOR2_X1 U635 ( .A(KEYINPUT59), .B(KEYINPUT65), .ZN(n504) );
  NAND2_X1 U636 ( .A1(n764), .A2(G953), .ZN(n505) );
  XNOR2_X1 U637 ( .A(n557), .B(G116), .ZN(n558) );
  NAND2_X1 U638 ( .A1(n621), .A2(n505), .ZN(n524) );
  INV_X1 U639 ( .A(n584), .ZN(n585) );
  INV_X1 U640 ( .A(KEYINPUT31), .ZN(n611) );
  XNOR2_X1 U641 ( .A(n503), .B(n544), .ZN(n545) );
  XNOR2_X1 U642 ( .A(n611), .B(KEYINPUT98), .ZN(n612) );
  XNOR2_X1 U643 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U644 ( .A(n546), .B(n545), .ZN(n755) );
  NOR2_X1 U645 ( .A1(G952), .A2(n709), .ZN(n756) );
  XNOR2_X1 U646 ( .A(n630), .B(n629), .ZN(n782) );
  INV_X1 U647 ( .A(n547), .ZN(n712) );
  XNOR2_X1 U648 ( .A(G116), .B(G107), .ZN(n506) );
  XNOR2_X1 U649 ( .A(n506), .B(G122), .ZN(n583) );
  XOR2_X1 U650 ( .A(n583), .B(KEYINPUT16), .Z(n511) );
  INV_X1 U651 ( .A(KEYINPUT3), .ZN(n507) );
  XNOR2_X1 U652 ( .A(n508), .B(n507), .ZN(n510) );
  XOR2_X1 U653 ( .A(KEYINPUT92), .B(G119), .Z(n509) );
  NAND2_X1 U654 ( .A1(n709), .A2(G224), .ZN(n512) );
  NAND2_X1 U655 ( .A1(n518), .A2(G210), .ZN(n516) );
  NAND2_X1 U656 ( .A1(G214), .A2(n518), .ZN(n674) );
  NAND2_X1 U657 ( .A1(G234), .A2(G237), .ZN(n520) );
  XNOR2_X1 U658 ( .A(n520), .B(KEYINPUT14), .ZN(n702) );
  NOR2_X1 U659 ( .A1(G902), .A2(n709), .ZN(n522) );
  NOR2_X1 U660 ( .A1(G953), .A2(G952), .ZN(n521) );
  NOR2_X1 U661 ( .A1(n522), .A2(n521), .ZN(n523) );
  AND2_X1 U662 ( .A1(n702), .A2(n523), .ZN(n621) );
  XNOR2_X1 U663 ( .A(G898), .B(KEYINPUT94), .ZN(n764) );
  INV_X1 U664 ( .A(KEYINPUT0), .ZN(n525) );
  XNOR2_X1 U665 ( .A(n526), .B(n525), .ZN(n597) );
  XNOR2_X1 U666 ( .A(n527), .B(KEYINPUT79), .ZN(n532) );
  NAND2_X1 U667 ( .A1(G227), .A2(n709), .ZN(n529) );
  XNOR2_X1 U668 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U669 ( .A(n530), .B(G140), .Z(n531) );
  XNOR2_X1 U670 ( .A(n532), .B(n531), .ZN(n534) );
  XNOR2_X1 U671 ( .A(n534), .B(n560), .ZN(n742) );
  XNOR2_X1 U672 ( .A(n770), .B(KEYINPUT24), .ZN(n546) );
  NAND2_X1 U673 ( .A1(n709), .A2(G234), .ZN(n540) );
  XNOR2_X1 U674 ( .A(n540), .B(n539), .ZN(n586) );
  XOR2_X1 U675 ( .A(G110), .B(G137), .Z(n542) );
  XNOR2_X1 U676 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U677 ( .A(n543), .B(KEYINPUT23), .Z(n544) );
  NOR2_X1 U678 ( .A1(G902), .A2(n755), .ZN(n552) );
  XOR2_X1 U679 ( .A(KEYINPUT95), .B(KEYINPUT25), .Z(n550) );
  NAND2_X1 U680 ( .A1(n547), .A2(G234), .ZN(n548) );
  XNOR2_X1 U681 ( .A(n548), .B(KEYINPUT20), .ZN(n553) );
  NAND2_X1 U682 ( .A1(G217), .A2(n553), .ZN(n549) );
  XNOR2_X1 U683 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U684 ( .A(KEYINPUT96), .B(KEYINPUT21), .Z(n555) );
  NAND2_X1 U685 ( .A1(G221), .A2(n553), .ZN(n554) );
  XOR2_X1 U686 ( .A(n555), .B(n554), .Z(n687) );
  XNOR2_X1 U687 ( .A(KEYINPUT97), .B(n687), .ZN(n598) );
  INV_X1 U688 ( .A(n607), .ZN(n684) );
  XNOR2_X1 U689 ( .A(KEYINPUT6), .B(KEYINPUT107), .ZN(n562) );
  AND2_X1 U690 ( .A1(n569), .A2(G210), .ZN(n559) );
  NOR2_X1 U691 ( .A1(n609), .A2(n363), .ZN(n563) );
  XNOR2_X1 U692 ( .A(KEYINPUT34), .B(KEYINPUT82), .ZN(n564) );
  XNOR2_X1 U693 ( .A(n565), .B(n564), .ZN(n592) );
  XNOR2_X1 U694 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U695 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n571) );
  NAND2_X1 U696 ( .A1(G214), .A2(n569), .ZN(n570) );
  XNOR2_X1 U697 ( .A(n573), .B(n572), .ZN(n574) );
  XOR2_X1 U698 ( .A(KEYINPUT13), .B(KEYINPUT102), .Z(n577) );
  XNOR2_X1 U699 ( .A(KEYINPUT101), .B(G475), .ZN(n576) );
  XNOR2_X1 U700 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U701 ( .A(KEYINPUT105), .B(G478), .ZN(n591) );
  XNOR2_X1 U702 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U703 ( .A(n583), .B(n582), .ZN(n589) );
  XOR2_X1 U704 ( .A(n585), .B(KEYINPUT103), .Z(n588) );
  NAND2_X1 U705 ( .A1(G217), .A2(n586), .ZN(n587) );
  NOR2_X1 U706 ( .A1(G902), .A2(n751), .ZN(n590) );
  INV_X1 U707 ( .A(n606), .ZN(n595) );
  NOR2_X1 U708 ( .A1(n605), .A2(n595), .ZN(n640) );
  NAND2_X1 U709 ( .A1(n592), .A2(n640), .ZN(n594) );
  XOR2_X1 U710 ( .A(KEYINPUT35), .B(KEYINPUT81), .Z(n593) );
  AND2_X1 U711 ( .A1(n595), .A2(n605), .ZN(n596) );
  NOR2_X1 U712 ( .A1(n653), .A2(n662), .ZN(n601) );
  NAND2_X1 U713 ( .A1(n603), .A2(n363), .ZN(n604) );
  NOR2_X1 U714 ( .A1(n688), .A2(n604), .ZN(n717) );
  NOR2_X1 U715 ( .A1(n730), .A2(n732), .ZN(n679) );
  XNOR2_X1 U716 ( .A(KEYINPUT86), .B(n679), .ZN(n645) );
  NAND2_X1 U717 ( .A1(n625), .A2(n686), .ZN(n608) );
  NOR2_X1 U718 ( .A1(n610), .A2(n608), .ZN(n719) );
  NOR2_X1 U719 ( .A1(n719), .A2(n733), .ZN(n614) );
  XNOR2_X1 U720 ( .A(n615), .B(KEYINPUT106), .ZN(n616) );
  NOR2_X1 U721 ( .A1(n717), .A2(n616), .ZN(n617) );
  XNOR2_X2 U722 ( .A(n619), .B(KEYINPUT45), .ZN(n710) );
  NAND2_X1 U723 ( .A1(G953), .A2(G900), .ZN(n620) );
  NAND2_X1 U724 ( .A1(n621), .A2(n620), .ZN(n631) );
  XOR2_X1 U725 ( .A(KEYINPUT30), .B(KEYINPUT112), .Z(n623) );
  XNOR2_X1 U726 ( .A(n624), .B(n623), .ZN(n626) );
  NAND2_X1 U727 ( .A1(n628), .A2(n732), .ZN(n738) );
  NAND2_X1 U728 ( .A1(KEYINPUT2), .A2(n738), .ZN(n627) );
  XOR2_X1 U729 ( .A(KEYINPUT84), .B(n627), .Z(n668) );
  NAND2_X1 U730 ( .A1(n628), .A2(n730), .ZN(n630) );
  XOR2_X1 U731 ( .A(KEYINPUT114), .B(KEYINPUT42), .Z(n639) );
  NOR2_X1 U732 ( .A1(n687), .A2(n631), .ZN(n649) );
  XNOR2_X1 U733 ( .A(n633), .B(KEYINPUT28), .ZN(n636) );
  XNOR2_X1 U734 ( .A(n634), .B(KEYINPUT113), .ZN(n635) );
  NAND2_X1 U735 ( .A1(n636), .A2(n635), .ZN(n644) );
  XNOR2_X1 U736 ( .A(n637), .B(KEYINPUT41), .ZN(n707) );
  NAND2_X1 U737 ( .A1(KEYINPUT47), .A2(n679), .ZN(n643) );
  NAND2_X1 U738 ( .A1(n728), .A2(n645), .ZN(n646) );
  XOR2_X1 U739 ( .A(KEYINPUT36), .B(KEYINPUT115), .Z(n655) );
  NAND2_X1 U740 ( .A1(n649), .A2(n674), .ZN(n650) );
  NOR2_X1 U741 ( .A1(n363), .A2(n650), .ZN(n651) );
  NAND2_X1 U742 ( .A1(n730), .A2(n651), .ZN(n652) );
  XNOR2_X1 U743 ( .A(n655), .B(n654), .ZN(n656) );
  INV_X1 U744 ( .A(n735), .ZN(n657) );
  AND2_X1 U745 ( .A1(n370), .A2(n657), .ZN(n658) );
  INV_X1 U746 ( .A(KEYINPUT71), .ZN(n660) );
  NAND2_X1 U747 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U748 ( .A(n663), .B(KEYINPUT43), .ZN(n665) );
  NAND2_X1 U749 ( .A1(n665), .A2(n664), .ZN(n739) );
  NAND2_X1 U750 ( .A1(n666), .A2(n739), .ZN(n667) );
  NAND2_X1 U751 ( .A1(n668), .A2(n670), .ZN(n669) );
  INV_X1 U752 ( .A(KEYINPUT2), .ZN(n671) );
  NOR2_X1 U753 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U754 ( .A1(n677), .A2(n676), .ZN(n681) );
  NOR2_X1 U755 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U756 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U757 ( .A1(n682), .A2(n706), .ZN(n700) );
  NOR2_X1 U758 ( .A1(n684), .A2(n448), .ZN(n685) );
  XOR2_X1 U759 ( .A(KEYINPUT50), .B(n685), .Z(n694) );
  XOR2_X1 U760 ( .A(KEYINPUT49), .B(KEYINPUT119), .Z(n690) );
  NAND2_X1 U761 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U762 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X1 U763 ( .A1(n429), .A2(n691), .ZN(n692) );
  XNOR2_X1 U764 ( .A(KEYINPUT120), .B(n692), .ZN(n693) );
  NAND2_X1 U765 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U766 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U767 ( .A(KEYINPUT51), .B(n697), .ZN(n698) );
  NOR2_X1 U768 ( .A1(n698), .A2(n707), .ZN(n699) );
  NOR2_X1 U769 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U770 ( .A(KEYINPUT52), .B(n701), .ZN(n704) );
  NAND2_X1 U771 ( .A1(n702), .A2(G952), .ZN(n703) );
  NOR2_X1 U772 ( .A1(n704), .A2(n703), .ZN(n705) );
  OR2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n708) );
  INV_X1 U774 ( .A(KEYINPUT63), .ZN(n716) );
  INV_X1 U775 ( .A(n710), .ZN(n757) );
  NAND2_X1 U776 ( .A1(KEYINPUT2), .A2(n712), .ZN(n713) );
  XOR2_X1 U777 ( .A(G101), .B(n717), .Z(G3) );
  NAND2_X1 U778 ( .A1(n719), .A2(n730), .ZN(n718) );
  XNOR2_X1 U779 ( .A(n718), .B(G104), .ZN(G6) );
  XOR2_X1 U780 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n721) );
  NAND2_X1 U781 ( .A1(n719), .A2(n732), .ZN(n720) );
  XNOR2_X1 U782 ( .A(n721), .B(n720), .ZN(n722) );
  XNOR2_X1 U783 ( .A(G107), .B(n722), .ZN(G9) );
  XOR2_X1 U784 ( .A(KEYINPUT29), .B(KEYINPUT117), .Z(n724) );
  NAND2_X1 U785 ( .A1(n732), .A2(n728), .ZN(n723) );
  XNOR2_X1 U786 ( .A(n724), .B(n723), .ZN(n726) );
  XOR2_X1 U787 ( .A(G128), .B(KEYINPUT116), .Z(n725) );
  XNOR2_X1 U788 ( .A(n726), .B(n725), .ZN(G30) );
  XNOR2_X1 U789 ( .A(n727), .B(G143), .ZN(G45) );
  NAND2_X1 U790 ( .A1(n728), .A2(n730), .ZN(n729) );
  XNOR2_X1 U791 ( .A(n729), .B(G146), .ZN(G48) );
  NAND2_X1 U792 ( .A1(n733), .A2(n730), .ZN(n731) );
  XNOR2_X1 U793 ( .A(n731), .B(G113), .ZN(G15) );
  NAND2_X1 U794 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U795 ( .A(n734), .B(G116), .ZN(G18) );
  XNOR2_X1 U796 ( .A(n735), .B(KEYINPUT118), .ZN(n736) );
  XNOR2_X1 U797 ( .A(n736), .B(KEYINPUT37), .ZN(n737) );
  XNOR2_X1 U798 ( .A(G125), .B(n737), .ZN(G27) );
  XNOR2_X1 U799 ( .A(G134), .B(n738), .ZN(G36) );
  XNOR2_X1 U800 ( .A(G140), .B(n739), .ZN(G42) );
  XOR2_X1 U801 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n741) );
  XNOR2_X1 U802 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n744) );
  XNOR2_X1 U803 ( .A(n428), .B(KEYINPUT57), .ZN(n743) );
  NOR2_X1 U804 ( .A1(n756), .A2(n745), .ZN(G54) );
  XNOR2_X1 U805 ( .A(KEYINPUT67), .B(KEYINPUT123), .ZN(n749) );
  XOR2_X1 U806 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n750) );
  NOR2_X1 U807 ( .A1(n756), .A2(n752), .ZN(G63) );
  NAND2_X1 U808 ( .A1(G217), .A2(n753), .ZN(n754) );
  NAND2_X1 U809 ( .A1(n709), .A2(n757), .ZN(n761) );
  NAND2_X1 U810 ( .A1(G953), .A2(G224), .ZN(n758) );
  XNOR2_X1 U811 ( .A(n758), .B(KEYINPUT61), .ZN(n759) );
  NAND2_X1 U812 ( .A1(n759), .A2(n764), .ZN(n760) );
  NAND2_X1 U813 ( .A1(n761), .A2(n760), .ZN(n768) );
  XOR2_X1 U814 ( .A(n762), .B(n763), .Z(n766) );
  NOR2_X1 U815 ( .A1(n709), .A2(n764), .ZN(n765) );
  NOR2_X1 U816 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U817 ( .A(n768), .B(n767), .ZN(G69) );
  XOR2_X1 U818 ( .A(n770), .B(n769), .Z(n774) );
  XOR2_X1 U819 ( .A(G227), .B(n774), .Z(n771) );
  NAND2_X1 U820 ( .A1(n771), .A2(G900), .ZN(n772) );
  NAND2_X1 U821 ( .A1(n772), .A2(G953), .ZN(n773) );
  XNOR2_X1 U822 ( .A(n773), .B(KEYINPUT126), .ZN(n777) );
  XNOR2_X1 U823 ( .A(n774), .B(n362), .ZN(n775) );
  NAND2_X1 U824 ( .A1(n775), .A2(n709), .ZN(n776) );
  NAND2_X1 U825 ( .A1(n777), .A2(n776), .ZN(G72) );
  XOR2_X1 U826 ( .A(G137), .B(n778), .Z(G39) );
  XOR2_X1 U827 ( .A(n779), .B(G122), .Z(G24) );
  XOR2_X1 U828 ( .A(n780), .B(G110), .Z(G12) );
  XNOR2_X1 U829 ( .A(G119), .B(n781), .ZN(G21) );
  XNOR2_X1 U830 ( .A(G131), .B(KEYINPUT127), .ZN(n783) );
  XNOR2_X1 U831 ( .A(n783), .B(n782), .ZN(G33) );
endmodule

