//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n780, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1021, new_n1022;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  INV_X1    g003(.A(G176gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT26), .ZN(new_n207));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n208), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT26), .ZN(new_n211));
  AOI22_X1  g010(.A1(new_n209), .A2(new_n211), .B1(G183gat), .B2(G190gat), .ZN(new_n212));
  INV_X1    g011(.A(G190gat), .ZN(new_n213));
  INV_X1    g012(.A(G183gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(new_n214), .B2(KEYINPUT27), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT65), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G183gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n216), .A2(new_n218), .A3(KEYINPUT27), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n215), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n216), .A2(new_n218), .A3(KEYINPUT66), .A4(KEYINPUT27), .ZN(new_n222));
  AOI21_X1  g021(.A(KEYINPUT28), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n214), .A2(KEYINPUT27), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT28), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n225), .A2(new_n215), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n212), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT1), .ZN(new_n228));
  INV_X1    g027(.A(G120gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G113gat), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n229), .A2(G113gat), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n228), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G134gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G127gat), .ZN(new_n235));
  INV_X1    g034(.A(G127gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G134gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n238), .B1(new_n235), .B2(new_n237), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n233), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT68), .B(G113gat), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n230), .B1(new_n243), .B2(new_n229), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n235), .A2(new_n237), .A3(new_n228), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  AND3_X1   g046(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n216), .A2(new_n218), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n250), .B1(new_n251), .B2(G190gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n208), .A2(KEYINPUT23), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT23), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n210), .B1(new_n206), .B2(new_n254), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n252), .A2(KEYINPUT25), .A3(new_n253), .A4(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n254), .B1(G169gat), .B2(G176gat), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n253), .B1(new_n257), .B2(new_n208), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT64), .ZN(new_n259));
  NAND2_X1  g058(.A1(G183gat), .A2(G190gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT24), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(G183gat), .A2(G190gat), .ZN(new_n263));
  NOR3_X1   g062(.A1(new_n262), .A2(new_n263), .A3(new_n248), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n249), .A2(new_n259), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n258), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n256), .B1(new_n266), .B2(KEYINPUT25), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n227), .A2(new_n247), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n247), .B1(new_n227), .B2(new_n267), .ZN(new_n269));
  INV_X1    g068(.A(G227gat), .ZN(new_n270));
  INV_X1    g069(.A(G233gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NOR3_X1   g072(.A1(new_n268), .A2(new_n269), .A3(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n203), .B1(new_n274), .B2(KEYINPUT33), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n227), .A2(new_n267), .ZN(new_n276));
  INV_X1    g075(.A(new_n241), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(new_n239), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n278), .A2(new_n233), .B1(new_n244), .B2(new_n245), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n227), .A2(new_n247), .A3(new_n267), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(new_n272), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT33), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(KEYINPUT69), .A3(new_n283), .ZN(new_n284));
  XOR2_X1   g083(.A(G15gat), .B(G43gat), .Z(new_n285));
  XNOR2_X1  g084(.A(new_n285), .B(KEYINPUT70), .ZN(new_n286));
  XNOR2_X1  g085(.A(G71gat), .B(G99gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n286), .B(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n288), .B1(new_n282), .B2(KEYINPUT32), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n275), .A2(new_n284), .A3(new_n289), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n282), .B(KEYINPUT32), .C1(new_n283), .C2(new_n288), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n272), .B1(new_n280), .B2(new_n281), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT34), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(KEYINPUT71), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n297));
  OAI21_X1  g096(.A(KEYINPUT34), .B1(new_n293), .B2(new_n297), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT73), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n292), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n296), .A2(new_n298), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n302), .A2(new_n291), .A3(new_n290), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n300), .B1(new_n292), .B2(new_n299), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n202), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n291), .ZN(new_n307));
  INV_X1    g106(.A(new_n288), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT32), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n308), .B1(new_n274), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT69), .B1(new_n282), .B2(new_n283), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n307), .B1(new_n312), .B2(new_n284), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n302), .B1(new_n313), .B2(KEYINPUT72), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n292), .A2(new_n299), .A3(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(KEYINPUT36), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n306), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT40), .ZN(new_n319));
  XNOR2_X1  g118(.A(G1gat), .B(G29gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n320), .B(KEYINPUT0), .ZN(new_n321));
  XNOR2_X1  g120(.A(G57gat), .B(G85gat), .ZN(new_n322));
  XOR2_X1   g121(.A(new_n321), .B(new_n322), .Z(new_n323));
  NAND2_X1  g122(.A1(G225gat), .A2(G233gat), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT78), .ZN(new_n325));
  INV_X1    g124(.A(G148gat), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n325), .B1(new_n326), .B2(G141gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(G141gat), .ZN(new_n328));
  INV_X1    g127(.A(G141gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n329), .A2(KEYINPUT78), .A3(G148gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n327), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(G155gat), .ZN(new_n336));
  OR2_X1    g135(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n337));
  NAND2_X1  g136(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT2), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n331), .B(new_n335), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n334), .B1(new_n332), .B2(new_n342), .ZN(new_n343));
  NOR3_X1   g142(.A1(KEYINPUT77), .A2(G155gat), .A3(G162gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n326), .A2(G141gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n329), .A2(G148gat), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n340), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n341), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT80), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n341), .A2(new_n349), .A3(KEYINPUT80), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n352), .A2(KEYINPUT3), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT81), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n352), .A2(KEYINPUT81), .A3(KEYINPUT3), .A4(new_n353), .ZN(new_n357));
  XOR2_X1   g156(.A(KEYINPUT82), .B(KEYINPUT3), .Z(new_n358));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n349), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n247), .ZN(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n356), .A2(new_n357), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n338), .ZN(new_n363));
  NOR2_X1   g162(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n364));
  OAI21_X1  g163(.A(G155gat), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n365), .A2(KEYINPUT2), .B1(new_n334), .B2(new_n333), .ZN(new_n366));
  AOI22_X1  g165(.A1(new_n366), .A2(new_n331), .B1(new_n348), .B2(new_n345), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n279), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT4), .B1(new_n247), .B2(new_n350), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n324), .B1(new_n362), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n352), .A2(new_n247), .A3(new_n353), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n279), .A2(new_n367), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n324), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT39), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n323), .B1(new_n372), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n360), .B1(new_n354), .B2(new_n355), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n379), .A2(new_n357), .B1(new_n369), .B2(new_n370), .ZN(new_n380));
  NOR3_X1   g179(.A1(new_n380), .A2(KEYINPUT39), .A3(new_n324), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n319), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT88), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g183(.A(KEYINPUT88), .B(new_n319), .C1(new_n378), .C2(new_n381), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT5), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n362), .A2(new_n387), .A3(new_n324), .A4(new_n371), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n369), .A2(new_n370), .A3(KEYINPUT83), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT83), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n279), .A2(new_n367), .A3(new_n390), .A4(new_n368), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n392), .A2(new_n362), .A3(new_n324), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT84), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n394), .B1(new_n375), .B2(new_n376), .ZN(new_n395));
  AOI211_X1 g194(.A(KEYINPUT84), .B(new_n324), .C1(new_n373), .C2(new_n374), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT5), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n388), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n323), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(G226gat), .A2(G233gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n401), .B(KEYINPUT75), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n276), .A2(new_n402), .ZN(new_n403));
  XOR2_X1   g202(.A(G211gat), .B(G218gat), .Z(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(G197gat), .A2(G204gat), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(G197gat), .A2(G204gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT74), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n411));
  NOR3_X1   g210(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  OR2_X1    g211(.A1(G197gat), .A2(G204gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n406), .ZN(new_n414));
  INV_X1    g213(.A(new_n411), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT74), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n405), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n411), .B1(new_n413), .B2(new_n406), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT74), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n404), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n401), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT29), .B1(new_n227), .B2(new_n267), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n403), .B(new_n421), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  XOR2_X1   g223(.A(G8gat), .B(G36gat), .Z(new_n425));
  XOR2_X1   g224(.A(G64gat), .B(G92gat), .Z(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  AOI21_X1  g226(.A(new_n401), .B1(new_n227), .B2(new_n267), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT29), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n276), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n402), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n424), .B(new_n427), .C1(new_n432), .C2(new_n421), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT30), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n410), .B1(new_n409), .B2(new_n411), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n404), .B1(new_n436), .B2(new_n419), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n412), .A2(new_n405), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n423), .A2(new_n402), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n439), .B1(new_n440), .B2(new_n428), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n441), .A2(KEYINPUT30), .A3(new_n424), .A4(new_n427), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n424), .B1(new_n432), .B2(new_n421), .ZN(new_n443));
  XOR2_X1   g242(.A(new_n427), .B(KEYINPUT76), .Z(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n435), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT39), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n372), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n377), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n449), .B1(new_n380), .B2(new_n324), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n448), .A2(new_n450), .A3(KEYINPUT40), .A4(new_n323), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n400), .A2(new_n446), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n386), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT38), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n427), .B1(new_n443), .B2(KEYINPUT37), .ZN(new_n455));
  XNOR2_X1  g254(.A(KEYINPUT89), .B(KEYINPUT37), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n424), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n454), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n403), .B(new_n439), .C1(new_n422), .C2(new_n423), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n459), .B(KEYINPUT37), .C1(new_n432), .C2(new_n439), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n444), .A2(new_n454), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n457), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n433), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n323), .B(new_n388), .C1(new_n393), .C2(new_n397), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT6), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n392), .A2(new_n362), .A3(new_n324), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n468), .B(KEYINPUT5), .C1(new_n395), .C2(new_n396), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n323), .B1(new_n469), .B2(new_n388), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n400), .A2(new_n466), .A3(new_n465), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n464), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(G228gat), .A2(G233gat), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n429), .B1(new_n437), .B2(new_n438), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n367), .B1(new_n475), .B2(new_n358), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n421), .B1(new_n429), .B2(new_n359), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G22gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n359), .A2(new_n429), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(new_n439), .A3(KEYINPUT85), .ZN(new_n481));
  INV_X1    g280(.A(new_n474), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT3), .B1(new_n421), .B2(new_n429), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n352), .A2(new_n353), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n481), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n477), .A2(KEYINPUT85), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n478), .B(new_n479), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT86), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G78gat), .B(G106gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(KEYINPUT31), .B(G50gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n478), .B1(new_n485), .B2(new_n486), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(G22gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n487), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n495), .A2(KEYINPUT86), .A3(new_n487), .A4(new_n492), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n453), .A2(new_n473), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT87), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n497), .A2(KEYINPUT87), .A3(new_n498), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n446), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n467), .A2(new_n470), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n398), .A2(KEYINPUT6), .A3(new_n399), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n318), .A2(new_n500), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n314), .A2(new_n316), .A3(new_n499), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT35), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n304), .A2(new_n305), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n446), .B1(new_n471), .B2(new_n472), .ZN(new_n514));
  AND2_X1   g313(.A1(new_n497), .A2(new_n498), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n515), .A2(KEYINPUT35), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n513), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT96), .ZN(new_n520));
  INV_X1    g319(.A(G50gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G43gat), .ZN(new_n522));
  INV_X1    g321(.A(G43gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G50gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(new_n524), .A3(KEYINPUT15), .ZN(new_n525));
  NOR3_X1   g324(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n526));
  OR2_X1    g325(.A1(new_n526), .A2(KEYINPUT90), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(KEYINPUT90), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n527), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT91), .B(G29gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(G36gat), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n525), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT93), .ZN(new_n534));
  NAND2_X1  g333(.A1(KEYINPUT92), .A2(G43gat), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  NOR2_X1   g335(.A1(KEYINPUT92), .A2(G43gat), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n534), .B(new_n521), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT15), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT92), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n523), .ZN(new_n541));
  AOI21_X1  g340(.A(G50gat), .B1(new_n541), .B2(new_n535), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n524), .A2(KEYINPUT93), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n538), .B(new_n539), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n526), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(new_n529), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n547), .A2(new_n532), .A3(new_n525), .ZN(new_n548));
  OAI21_X1  g347(.A(KEYINPUT94), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n547), .A2(new_n532), .A3(new_n525), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT94), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(new_n544), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n533), .B1(new_n549), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(G1gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT16), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n479), .A2(G15gat), .ZN(new_n556));
  INV_X1    g355(.A(G15gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(G22gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n559), .A2(KEYINPUT95), .ZN(new_n560));
  XNOR2_X1  g359(.A(G15gat), .B(G22gat), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT95), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n555), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n559), .A2(KEYINPUT95), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n561), .A2(new_n562), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(new_n566), .A3(new_n554), .ZN(new_n567));
  INV_X1    g366(.A(G8gat), .ZN(new_n568));
  AND3_X1   g367(.A1(new_n564), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n568), .B1(new_n564), .B2(new_n567), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n520), .B1(new_n553), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n533), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n550), .A2(new_n544), .A3(new_n551), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n551), .B1(new_n550), .B2(new_n544), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n570), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n564), .A2(new_n568), .A3(new_n567), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n576), .A2(new_n579), .A3(KEYINPUT96), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n572), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G229gat), .A2(G233gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT17), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n576), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g383(.A(KEYINPUT17), .B(new_n573), .C1(new_n574), .C2(new_n575), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(new_n571), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n581), .A2(new_n582), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT18), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n581), .A2(new_n586), .A3(KEYINPUT18), .A4(new_n582), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n553), .A2(new_n571), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n581), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n582), .B(KEYINPUT13), .Z(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n589), .A2(new_n590), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G113gat), .B(G141gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(G197gat), .ZN(new_n597));
  XOR2_X1   g396(.A(KEYINPUT11), .B(G169gat), .Z(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(KEYINPUT12), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n595), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT97), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n589), .A2(new_n594), .A3(new_n600), .A4(new_n590), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n595), .A2(KEYINPUT97), .A3(new_n601), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G85gat), .A2(G92gat), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT7), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NOR2_X1   g409(.A1(G85gat), .A2(G92gat), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G99gat), .A2(G106gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT8), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT101), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT101), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n612), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n610), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(G99gat), .B(G106gat), .Z(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(KEYINPUT103), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n610), .ZN(new_n623));
  INV_X1    g422(.A(new_n618), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n617), .B1(new_n612), .B2(new_n614), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT103), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n626), .A2(new_n627), .A3(new_n620), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n623), .B(new_n621), .C1(new_n624), .C2(new_n625), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n629), .A2(KEYINPUT102), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT102), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n631), .B1(new_n619), .B2(new_n621), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n622), .B(new_n628), .C1(new_n630), .C2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n633), .A2(new_n553), .ZN(new_n634));
  AND2_X1   g433(.A1(G232gat), .A2(G233gat), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n634), .B1(KEYINPUT41), .B2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(G190gat), .B(G218gat), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n584), .A2(new_n585), .A3(new_n633), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G134gat), .B(G162gat), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n638), .B1(new_n636), .B2(new_n639), .ZN(new_n645));
  OR3_X1    g444(.A1(new_n640), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n644), .B1(new_n640), .B2(new_n645), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n626), .A2(new_n620), .ZN(new_n650));
  XOR2_X1   g449(.A(G57gat), .B(G64gat), .Z(new_n651));
  INV_X1    g450(.A(KEYINPUT9), .ZN(new_n652));
  INV_X1    g451(.A(G71gat), .ZN(new_n653));
  INV_X1    g452(.A(G78gat), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT98), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g457(.A(G71gat), .B(G78gat), .Z(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n656), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  OAI211_X1 g460(.A(new_n655), .B(new_n651), .C1(new_n659), .C2(new_n657), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n650), .A2(new_n663), .A3(new_n629), .ZN(new_n664));
  INV_X1    g463(.A(new_n663), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n664), .B1(new_n633), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(G230gat), .A2(G233gat), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT104), .ZN(new_n669));
  AOI211_X1 g468(.A(KEYINPUT10), .B(new_n664), .C1(new_n633), .C2(new_n665), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n663), .A2(KEYINPUT10), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n633), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n667), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(G120gat), .B(G148gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(G176gat), .B(G204gat), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n674), .B(new_n675), .Z(new_n676));
  NAND3_X1  g475(.A1(new_n669), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n676), .ZN(new_n678));
  INV_X1    g477(.A(new_n667), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n633), .A2(new_n665), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT10), .ZN(new_n681));
  INV_X1    g480(.A(new_n664), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n633), .A2(new_n671), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n679), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n678), .B1(new_n685), .B2(new_n668), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n677), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n663), .A2(KEYINPUT21), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n688), .B(new_n689), .Z(new_n690));
  AOI21_X1  g489(.A(new_n579), .B1(KEYINPUT21), .B2(new_n663), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(G127gat), .B(G155gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT20), .ZN(new_n694));
  NAND2_X1  g493(.A1(G231gat), .A2(G233gat), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT99), .Z(new_n696));
  XNOR2_X1  g495(.A(new_n694), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(G183gat), .B(G211gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n692), .B(new_n699), .Z(new_n700));
  NOR4_X1   g499(.A1(new_n607), .A2(new_n649), .A3(new_n687), .A4(new_n700), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n519), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT105), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(KEYINPUT105), .B1(new_n471), .B2(new_n472), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g508(.A(KEYINPUT16), .B(G8gat), .Z(new_n710));
  NAND3_X1  g509(.A1(new_n702), .A2(new_n446), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT42), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n702), .ZN(new_n714));
  OAI21_X1  g513(.A(G8gat), .B1(new_n714), .B2(new_n505), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n711), .A2(new_n712), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n713), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1325gat));
  OAI21_X1  g518(.A(G15gat), .B1(new_n714), .B2(new_n318), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n702), .A2(new_n557), .A3(new_n513), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(G1326gat));
  NAND2_X1  g521(.A1(new_n702), .A2(new_n504), .ZN(new_n723));
  XNOR2_X1  g522(.A(KEYINPUT43), .B(G22gat), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n723), .B(new_n724), .ZN(G1327gat));
  NAND2_X1  g524(.A1(new_n519), .A2(new_n649), .ZN(new_n726));
  INV_X1    g525(.A(new_n700), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n607), .A2(new_n687), .A3(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n531), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n730), .A2(new_n731), .A3(new_n707), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT45), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n515), .B1(new_n386), .B2(new_n452), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n734), .A2(new_n473), .B1(new_n504), .B2(new_n508), .ZN(new_n735));
  AOI22_X1  g534(.A1(new_n735), .A2(new_n318), .B1(new_n512), .B2(new_n517), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT44), .B1(new_n736), .B2(new_n648), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n648), .B1(new_n510), .B2(new_n518), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n729), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n531), .B1(new_n742), .B2(new_n706), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n733), .A2(new_n743), .ZN(G1328gat));
  NOR4_X1   g543(.A1(new_n726), .A2(G36gat), .A3(new_n505), .A4(new_n729), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT46), .ZN(new_n746));
  OAI21_X1  g545(.A(G36gat), .B1(new_n742), .B2(new_n505), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(G1329gat));
  NAND2_X1  g547(.A1(new_n541), .A2(new_n535), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n749), .B1(new_n742), .B2(new_n318), .ZN(new_n750));
  NAND2_X1  g549(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n751));
  NOR2_X1   g550(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n304), .A2(new_n305), .A3(new_n749), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n752), .B1(new_n730), .B2(new_n753), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n750), .A2(new_n751), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n751), .B1(new_n750), .B2(new_n754), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(G1330gat));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n504), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(G50gat), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n730), .A2(new_n521), .A3(new_n504), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n521), .B1(new_n741), .B2(new_n515), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(KEYINPUT48), .ZN(new_n763));
  OAI22_X1  g562(.A1(new_n761), .A2(KEYINPUT48), .B1(new_n762), .B2(new_n763), .ZN(G1331gat));
  NOR2_X1   g563(.A1(new_n649), .A2(new_n700), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n765), .A2(new_n607), .A3(new_n687), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n519), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n707), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g569(.A(new_n446), .B(KEYINPUT109), .Z(new_n771));
  NOR2_X1   g570(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n773));
  AND2_X1   g572(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(new_n772), .B2(new_n773), .ZN(G1333gat));
  OAI21_X1  g575(.A(G71gat), .B1(new_n767), .B2(new_n318), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n513), .A2(new_n653), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n767), .B2(new_n778), .ZN(new_n779));
  XOR2_X1   g578(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n780));
  XNOR2_X1  g579(.A(new_n779), .B(new_n780), .ZN(G1334gat));
  NAND2_X1  g580(.A1(new_n768), .A2(new_n504), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(G78gat), .ZN(G1335gat));
  INV_X1    g582(.A(G85gat), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n737), .A2(new_n740), .ZN(new_n785));
  INV_X1    g584(.A(new_n607), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(new_n727), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(new_n687), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n785), .A2(new_n707), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n784), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n792), .B2(new_n791), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT51), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(new_n726), .B2(new_n788), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n738), .A2(KEYINPUT51), .A3(new_n787), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n798), .A2(new_n784), .A3(new_n687), .A4(new_n707), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n794), .A2(new_n799), .ZN(G1336gat));
  INV_X1    g599(.A(G92gat), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n771), .A2(new_n789), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n798), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(KEYINPUT112), .A2(KEYINPUT52), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n785), .A2(new_n790), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(new_n771), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G92gat), .ZN(new_n808));
  OAI211_X1 g607(.A(new_n803), .B(new_n804), .C1(new_n806), .C2(new_n808), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n798), .A2(new_n801), .A3(new_n802), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n785), .A2(new_n446), .A3(new_n790), .ZN(new_n811));
  AOI22_X1  g610(.A1(new_n810), .A2(KEYINPUT112), .B1(G92gat), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n809), .B1(new_n812), .B2(new_n807), .ZN(G1337gat));
  OAI21_X1  g612(.A(G99gat), .B1(new_n805), .B2(new_n318), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n789), .A2(G99gat), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n798), .A2(new_n513), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(G1338gat));
  OAI21_X1  g616(.A(G106gat), .B1(new_n805), .B2(new_n499), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n789), .A2(G106gat), .A3(new_n499), .ZN(new_n820));
  INV_X1    g619(.A(new_n797), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT51), .B1(new_n738), .B2(new_n787), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n818), .A2(new_n819), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT113), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT44), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n826), .B1(new_n519), .B2(new_n649), .ZN(new_n827));
  INV_X1    g626(.A(new_n739), .ZN(new_n828));
  AOI211_X1 g627(.A(new_n648), .B(new_n828), .C1(new_n510), .C2(new_n518), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n504), .B(new_n790), .C1(new_n827), .C2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(G106gat), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n823), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n825), .B1(new_n832), .B2(KEYINPUT53), .ZN(new_n833));
  AOI211_X1 g632(.A(KEYINPUT113), .B(new_n819), .C1(new_n831), .C2(new_n823), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n824), .B1(new_n833), .B2(new_n834), .ZN(G1339gat));
  INV_X1    g634(.A(new_n771), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n765), .A2(new_n607), .A3(new_n789), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n676), .B1(new_n685), .B2(new_n838), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n683), .A2(KEYINPUT114), .A3(new_n679), .A4(new_n684), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n673), .A2(new_n840), .A3(KEYINPUT54), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n672), .B1(new_n666), .B2(new_n681), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT114), .B1(new_n842), .B2(new_n679), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n839), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n839), .B(KEYINPUT55), .C1(new_n841), .C2(new_n843), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n677), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n592), .A2(new_n593), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n582), .B1(new_n581), .B2(new_n586), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n599), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n646), .A2(new_n604), .A3(new_n647), .A4(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n687), .A2(new_n604), .A3(new_n851), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n854), .B1(new_n607), .B2(new_n848), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n853), .B1(new_n855), .B2(new_n648), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n837), .B1(new_n856), .B2(new_n727), .ZN(new_n857));
  INV_X1    g656(.A(new_n511), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n857), .A2(new_n858), .A3(new_n707), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n847), .A2(new_n677), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n862), .A2(new_n605), .A3(new_n606), .A4(new_n846), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n649), .B1(new_n863), .B2(new_n854), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n700), .B1(new_n864), .B2(new_n853), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n706), .B1(new_n865), .B2(new_n837), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(KEYINPUT115), .A3(new_n858), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n836), .B1(new_n861), .B2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n243), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n869), .A3(new_n786), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n504), .B1(new_n865), .B2(new_n837), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n706), .A2(new_n836), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n513), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(G113gat), .B1(new_n875), .B2(new_n607), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n870), .A2(new_n876), .ZN(G1340gat));
  NOR3_X1   g676(.A1(new_n875), .A2(new_n229), .A3(new_n789), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n868), .A2(new_n687), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(new_n229), .ZN(G1341gat));
  NAND3_X1  g679(.A1(new_n868), .A2(new_n236), .A3(new_n727), .ZN(new_n881));
  OAI21_X1  g680(.A(G127gat), .B1(new_n875), .B2(new_n700), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(G1342gat));
  NAND2_X1  g682(.A1(new_n861), .A2(new_n867), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n648), .A2(new_n446), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n886), .A2(G134gat), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n871), .A2(new_n649), .A3(new_n874), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(G134gat), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT117), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n889), .A2(KEYINPUT117), .A3(G134gat), .ZN(new_n893));
  AOI22_X1  g692(.A1(KEYINPUT56), .A2(new_n888), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n888), .A2(KEYINPUT116), .A3(KEYINPUT56), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT116), .ZN(new_n896));
  INV_X1    g695(.A(new_n887), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n897), .B1(new_n861), .B2(new_n867), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT56), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n894), .B1(new_n895), .B2(new_n900), .ZN(G1343gat));
  NAND2_X1  g700(.A1(new_n872), .A2(new_n318), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n857), .A2(new_n515), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT57), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n504), .A2(KEYINPUT57), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n846), .A2(KEYINPUT118), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n844), .A2(new_n909), .A3(new_n845), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n908), .A2(new_n862), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n854), .B1(new_n911), .B2(new_n607), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n648), .ZN(new_n913));
  INV_X1    g712(.A(new_n853), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n727), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(new_n837), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n907), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n902), .B1(new_n905), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n329), .B1(new_n918), .B2(new_n786), .ZN(new_n919));
  INV_X1    g718(.A(new_n318), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n920), .A2(new_n499), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n786), .A2(new_n329), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT120), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n866), .A2(new_n771), .A3(new_n921), .A4(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT58), .ZN(new_n926));
  AOI211_X1 g725(.A(KEYINPUT121), .B(new_n926), .C1(new_n924), .C2(KEYINPUT119), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n857), .A2(new_n707), .A3(new_n771), .A4(new_n921), .ZN(new_n929));
  INV_X1    g728(.A(new_n923), .ZN(new_n930));
  OAI21_X1  g729(.A(KEYINPUT119), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n928), .B1(new_n931), .B2(KEYINPUT58), .ZN(new_n932));
  OAI22_X1  g731(.A1(new_n919), .A2(new_n925), .B1(new_n927), .B2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n902), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n910), .A2(new_n677), .A3(new_n847), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n786), .A2(new_n935), .A3(new_n908), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n649), .B1(new_n936), .B2(new_n854), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n700), .B1(new_n937), .B2(new_n853), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n906), .B1(new_n938), .B2(new_n837), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT57), .B1(new_n857), .B2(new_n515), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n786), .B(new_n934), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n925), .B1(new_n941), .B2(G141gat), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n931), .A2(KEYINPUT58), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT121), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n931), .A2(new_n928), .A3(KEYINPUT58), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n942), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n933), .A2(new_n946), .ZN(G1344gat));
  INV_X1    g746(.A(new_n929), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n948), .A2(new_n326), .A3(new_n687), .ZN(new_n949));
  AOI211_X1 g748(.A(KEYINPUT59), .B(new_n326), .C1(new_n918), .C2(new_n687), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT59), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n837), .B(KEYINPUT122), .ZN(new_n952));
  OAI211_X1 g751(.A(new_n904), .B(new_n504), .C1(new_n952), .C2(new_n915), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n903), .A2(KEYINPUT57), .ZN(new_n954));
  NAND4_X1  g753(.A1(new_n953), .A2(new_n954), .A3(new_n934), .A4(new_n687), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n951), .B1(new_n955), .B2(G148gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n949), .B1(new_n950), .B2(new_n956), .ZN(G1345gat));
  AOI21_X1  g756(.A(G155gat), .B1(new_n948), .B2(new_n727), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n700), .A2(new_n336), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT123), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n958), .B1(new_n918), .B2(new_n960), .ZN(G1346gat));
  NOR2_X1   g760(.A1(new_n363), .A2(new_n364), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n866), .A2(new_n962), .A3(new_n885), .A4(new_n921), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n918), .A2(new_n649), .ZN(new_n964));
  INV_X1    g763(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n963), .B1(new_n965), .B2(new_n962), .ZN(G1347gat));
  AND3_X1   g765(.A1(new_n706), .A2(new_n513), .A3(new_n446), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n871), .A2(new_n967), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n968), .A2(new_n204), .A3(new_n607), .ZN(new_n969));
  AOI21_X1  g768(.A(KEYINPUT124), .B1(new_n857), .B2(new_n706), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n857), .A2(KEYINPUT124), .A3(new_n706), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n511), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n973), .A2(new_n786), .A3(new_n836), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n969), .B1(new_n974), .B2(new_n204), .ZN(G1348gat));
  NAND3_X1  g774(.A1(new_n973), .A2(new_n205), .A3(new_n802), .ZN(new_n976));
  OAI21_X1  g775(.A(G176gat), .B1(new_n968), .B2(new_n789), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(G1349gat));
  OR2_X1    g777(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n971), .A2(new_n972), .ZN(new_n980));
  OR2_X1    g779(.A1(new_n214), .A2(KEYINPUT27), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n727), .A2(new_n981), .A3(new_n224), .ZN(new_n982));
  INV_X1    g781(.A(new_n982), .ZN(new_n983));
  NAND4_X1  g782(.A1(new_n980), .A2(new_n858), .A3(new_n836), .A4(new_n983), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n871), .A2(new_n727), .A3(new_n967), .ZN(new_n985));
  AOI22_X1  g784(.A1(new_n985), .A2(new_n251), .B1(KEYINPUT125), .B2(KEYINPUT60), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n979), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT124), .ZN(new_n988));
  AOI211_X1 g787(.A(new_n988), .B(new_n707), .C1(new_n865), .C2(new_n837), .ZN(new_n989));
  OAI211_X1 g788(.A(new_n858), .B(new_n836), .C1(new_n989), .C2(new_n970), .ZN(new_n990));
  OAI211_X1 g789(.A(new_n986), .B(new_n979), .C1(new_n990), .C2(new_n982), .ZN(new_n991));
  INV_X1    g790(.A(new_n991), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n987), .A2(new_n992), .ZN(G1350gat));
  OAI21_X1  g792(.A(G190gat), .B1(new_n968), .B2(new_n648), .ZN(new_n994));
  NOR2_X1   g793(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n649), .A2(new_n213), .ZN(new_n997));
  XNOR2_X1  g796(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n998));
  OAI221_X1 g797(.A(new_n996), .B1(new_n990), .B2(new_n997), .C1(new_n994), .C2(new_n998), .ZN(G1351gat));
  NOR3_X1   g798(.A1(new_n707), .A2(new_n920), .A3(new_n505), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n953), .A2(new_n954), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g800(.A(G197gat), .B1(new_n1001), .B2(new_n607), .ZN(new_n1002));
  NOR3_X1   g801(.A1(new_n920), .A2(new_n499), .A3(new_n771), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n980), .A2(new_n1003), .ZN(new_n1004));
  OR2_X1    g803(.A1(new_n607), .A2(G197gat), .ZN(new_n1005));
  OAI21_X1  g804(.A(new_n1002), .B1(new_n1004), .B2(new_n1005), .ZN(G1352gat));
  NAND4_X1  g805(.A1(new_n953), .A2(new_n954), .A3(new_n1000), .A4(new_n687), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n789), .A2(G204gat), .ZN(new_n1008));
  OAI211_X1 g807(.A(new_n1003), .B(new_n1008), .C1(new_n989), .C2(new_n970), .ZN(new_n1009));
  AOI22_X1  g808(.A1(new_n1007), .A2(G204gat), .B1(new_n1009), .B2(KEYINPUT62), .ZN(new_n1010));
  NOR2_X1   g809(.A1(new_n1009), .A2(KEYINPUT62), .ZN(new_n1011));
  INV_X1    g810(.A(KEYINPUT127), .ZN(new_n1012));
  NOR2_X1   g811(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NOR3_X1   g812(.A1(new_n1009), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1010), .B1(new_n1013), .B2(new_n1014), .ZN(G1353gat));
  NAND4_X1  g814(.A1(new_n953), .A2(new_n954), .A3(new_n1000), .A4(new_n727), .ZN(new_n1016));
  AND3_X1   g815(.A1(new_n1016), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1017));
  AOI21_X1  g816(.A(KEYINPUT63), .B1(new_n1016), .B2(G211gat), .ZN(new_n1018));
  OR2_X1    g817(.A1(new_n700), .A2(G211gat), .ZN(new_n1019));
  OAI22_X1  g818(.A1(new_n1017), .A2(new_n1018), .B1(new_n1004), .B2(new_n1019), .ZN(G1354gat));
  OAI21_X1  g819(.A(G218gat), .B1(new_n1001), .B2(new_n648), .ZN(new_n1021));
  OR2_X1    g820(.A1(new_n648), .A2(G218gat), .ZN(new_n1022));
  OAI21_X1  g821(.A(new_n1021), .B1(new_n1004), .B2(new_n1022), .ZN(G1355gat));
endmodule


