

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U550 ( .A1(n570), .A2(n569), .ZN(n963) );
  NOR2_X2 U551 ( .A1(G543), .A2(n530), .ZN(n528) );
  NOR2_X1 U552 ( .A1(n567), .A2(n566), .ZN(n568) );
  AND2_X2 U553 ( .A1(n521), .A2(G2104), .ZN(n894) );
  NOR2_X1 U554 ( .A1(G651), .A2(n628), .ZN(n637) );
  NOR2_X1 U555 ( .A1(n773), .A2(n759), .ZN(n514) );
  XNOR2_X1 U556 ( .A(n718), .B(KEYINPUT30), .ZN(n719) );
  XNOR2_X1 U557 ( .A(n720), .B(n719), .ZN(n721) );
  AND2_X1 U558 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U559 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U560 ( .A1(n527), .A2(n526), .ZN(G160) );
  XOR2_X1 U561 ( .A(KEYINPUT68), .B(KEYINPUT23), .Z(n516) );
  INV_X1 U562 ( .A(G2105), .ZN(n521) );
  NAND2_X1 U563 ( .A1(G101), .A2(n894), .ZN(n515) );
  XNOR2_X1 U564 ( .A(n516), .B(n515), .ZN(n520) );
  INV_X1 U565 ( .A(G2105), .ZN(n517) );
  NOR2_X4 U566 ( .A1(G2104), .A2(n517), .ZN(n901) );
  NAND2_X1 U567 ( .A1(G125), .A2(n901), .ZN(n518) );
  XOR2_X1 U568 ( .A(n518), .B(KEYINPUT67), .Z(n519) );
  NAND2_X1 U569 ( .A1(n520), .A2(n519), .ZN(n527) );
  AND2_X1 U570 ( .A1(G2104), .A2(G2105), .ZN(n899) );
  NAND2_X1 U571 ( .A1(n899), .A2(G113), .ZN(n525) );
  XNOR2_X1 U572 ( .A(KEYINPUT69), .B(KEYINPUT17), .ZN(n523) );
  NOR2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n522) );
  XNOR2_X1 U574 ( .A(n523), .B(n522), .ZN(n539) );
  NAND2_X1 U575 ( .A1(n539), .A2(G137), .ZN(n524) );
  NAND2_X1 U576 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U577 ( .A(G651), .B(KEYINPUT70), .Z(n530) );
  XOR2_X2 U578 ( .A(KEYINPUT1), .B(n528), .Z(n639) );
  NAND2_X1 U579 ( .A1(G64), .A2(n639), .ZN(n529) );
  XNOR2_X1 U580 ( .A(n529), .B(KEYINPUT71), .ZN(n538) );
  XOR2_X1 U581 ( .A(G543), .B(KEYINPUT0), .Z(n628) );
  NOR2_X1 U582 ( .A1(n628), .A2(n530), .ZN(n643) );
  NAND2_X1 U583 ( .A1(n643), .A2(G77), .ZN(n533) );
  NOR2_X1 U584 ( .A1(G543), .A2(G651), .ZN(n531) );
  XNOR2_X1 U585 ( .A(n531), .B(KEYINPUT66), .ZN(n640) );
  NAND2_X1 U586 ( .A1(G90), .A2(n640), .ZN(n532) );
  NAND2_X1 U587 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U588 ( .A(n534), .B(KEYINPUT9), .ZN(n536) );
  NAND2_X1 U589 ( .A1(G52), .A2(n637), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U591 ( .A1(n538), .A2(n537), .ZN(G171) );
  AND2_X1 U592 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U593 ( .A(G132), .ZN(G219) );
  INV_X1 U594 ( .A(G82), .ZN(G220) );
  INV_X1 U595 ( .A(G120), .ZN(G236) );
  INV_X1 U596 ( .A(G69), .ZN(G235) );
  INV_X1 U597 ( .A(G108), .ZN(G238) );
  NAND2_X1 U598 ( .A1(G102), .A2(n894), .ZN(n542) );
  INV_X1 U599 ( .A(n539), .ZN(n540) );
  INV_X1 U600 ( .A(n540), .ZN(n895) );
  NAND2_X1 U601 ( .A1(G138), .A2(n895), .ZN(n541) );
  NAND2_X1 U602 ( .A1(n542), .A2(n541), .ZN(n546) );
  NAND2_X1 U603 ( .A1(G126), .A2(n901), .ZN(n544) );
  NAND2_X1 U604 ( .A1(G114), .A2(n899), .ZN(n543) );
  NAND2_X1 U605 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U606 ( .A1(n546), .A2(n545), .ZN(G164) );
  NAND2_X1 U607 ( .A1(G63), .A2(n639), .ZN(n548) );
  NAND2_X1 U608 ( .A1(G51), .A2(n637), .ZN(n547) );
  NAND2_X1 U609 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U610 ( .A(KEYINPUT6), .B(n549), .ZN(n555) );
  NAND2_X1 U611 ( .A1(G89), .A2(n640), .ZN(n550) );
  XNOR2_X1 U612 ( .A(n550), .B(KEYINPUT4), .ZN(n552) );
  NAND2_X1 U613 ( .A1(G76), .A2(n643), .ZN(n551) );
  NAND2_X1 U614 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U615 ( .A(n553), .B(KEYINPUT5), .Z(n554) );
  NOR2_X1 U616 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U617 ( .A(KEYINPUT77), .B(n556), .Z(n557) );
  XOR2_X1 U618 ( .A(KEYINPUT7), .B(n557), .Z(G168) );
  XOR2_X1 U619 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U620 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n559) );
  NAND2_X1 U621 ( .A1(G7), .A2(G661), .ZN(n558) );
  XNOR2_X1 U622 ( .A(n559), .B(n558), .ZN(G223) );
  INV_X1 U623 ( .A(G223), .ZN(n828) );
  NAND2_X1 U624 ( .A1(n828), .A2(G567), .ZN(n560) );
  XOR2_X1 U625 ( .A(KEYINPUT11), .B(n560), .Z(G234) );
  NAND2_X1 U626 ( .A1(n639), .A2(G56), .ZN(n561) );
  XOR2_X1 U627 ( .A(KEYINPUT14), .B(n561), .Z(n567) );
  NAND2_X1 U628 ( .A1(G81), .A2(n640), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(KEYINPUT12), .ZN(n564) );
  NAND2_X1 U630 ( .A1(G68), .A2(n643), .ZN(n563) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U632 ( .A(KEYINPUT13), .B(n565), .Z(n566) );
  XNOR2_X1 U633 ( .A(n568), .B(KEYINPUT74), .ZN(n570) );
  NAND2_X1 U634 ( .A1(G43), .A2(n637), .ZN(n569) );
  INV_X1 U635 ( .A(G860), .ZN(n590) );
  OR2_X1 U636 ( .A1(n963), .A2(n590), .ZN(G153) );
  INV_X1 U637 ( .A(G171), .ZN(G301) );
  NAND2_X1 U638 ( .A1(G868), .A2(G301), .ZN(n581) );
  NAND2_X1 U639 ( .A1(G54), .A2(n637), .ZN(n571) );
  XNOR2_X1 U640 ( .A(n571), .B(KEYINPUT76), .ZN(n578) );
  NAND2_X1 U641 ( .A1(G79), .A2(n643), .ZN(n573) );
  NAND2_X1 U642 ( .A1(G66), .A2(n639), .ZN(n572) );
  NAND2_X1 U643 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U644 ( .A1(G92), .A2(n640), .ZN(n574) );
  XNOR2_X1 U645 ( .A(KEYINPUT75), .B(n574), .ZN(n575) );
  NOR2_X1 U646 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U647 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U648 ( .A(KEYINPUT15), .B(n579), .Z(n954) );
  INV_X1 U649 ( .A(G868), .ZN(n656) );
  NAND2_X1 U650 ( .A1(n954), .A2(n656), .ZN(n580) );
  NAND2_X1 U651 ( .A1(n581), .A2(n580), .ZN(G284) );
  NAND2_X1 U652 ( .A1(G65), .A2(n639), .ZN(n583) );
  NAND2_X1 U653 ( .A1(G53), .A2(n637), .ZN(n582) );
  NAND2_X1 U654 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U655 ( .A1(n643), .A2(G78), .ZN(n585) );
  NAND2_X1 U656 ( .A1(G91), .A2(n640), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U658 ( .A1(n587), .A2(n586), .ZN(n953) );
  XOR2_X1 U659 ( .A(n953), .B(KEYINPUT72), .Z(G299) );
  NOR2_X1 U660 ( .A1(G299), .A2(G868), .ZN(n589) );
  NOR2_X1 U661 ( .A1(G286), .A2(n656), .ZN(n588) );
  NOR2_X1 U662 ( .A1(n589), .A2(n588), .ZN(G297) );
  NAND2_X1 U663 ( .A1(n590), .A2(G559), .ZN(n591) );
  INV_X1 U664 ( .A(n954), .ZN(n607) );
  NAND2_X1 U665 ( .A1(n591), .A2(n607), .ZN(n592) );
  XNOR2_X1 U666 ( .A(n592), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U667 ( .A1(n954), .A2(n656), .ZN(n593) );
  XOR2_X1 U668 ( .A(KEYINPUT78), .B(n593), .Z(n594) );
  NOR2_X1 U669 ( .A1(G559), .A2(n594), .ZN(n596) );
  NOR2_X1 U670 ( .A1(G868), .A2(n963), .ZN(n595) );
  NOR2_X1 U671 ( .A1(n596), .A2(n595), .ZN(G282) );
  NAND2_X1 U672 ( .A1(G123), .A2(n901), .ZN(n597) );
  XOR2_X1 U673 ( .A(KEYINPUT18), .B(n597), .Z(n598) );
  XNOR2_X1 U674 ( .A(n598), .B(KEYINPUT79), .ZN(n600) );
  NAND2_X1 U675 ( .A1(G111), .A2(n899), .ZN(n599) );
  NAND2_X1 U676 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U677 ( .A1(G99), .A2(n894), .ZN(n602) );
  NAND2_X1 U678 ( .A1(G135), .A2(n895), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U680 ( .A1(n604), .A2(n603), .ZN(n1004) );
  XNOR2_X1 U681 ( .A(n1004), .B(G2096), .ZN(n606) );
  INV_X1 U682 ( .A(G2100), .ZN(n605) );
  NAND2_X1 U683 ( .A1(n606), .A2(n605), .ZN(G156) );
  NAND2_X1 U684 ( .A1(G559), .A2(n607), .ZN(n608) );
  XNOR2_X1 U685 ( .A(n963), .B(n608), .ZN(n654) );
  NOR2_X1 U686 ( .A1(n654), .A2(G860), .ZN(n617) );
  NAND2_X1 U687 ( .A1(n643), .A2(G80), .ZN(n610) );
  NAND2_X1 U688 ( .A1(G93), .A2(n640), .ZN(n609) );
  NAND2_X1 U689 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U690 ( .A1(G55), .A2(n637), .ZN(n611) );
  XNOR2_X1 U691 ( .A(KEYINPUT81), .B(n611), .ZN(n612) );
  NOR2_X1 U692 ( .A1(n613), .A2(n612), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n639), .A2(G67), .ZN(n614) );
  NAND2_X1 U694 ( .A1(n615), .A2(n614), .ZN(n657) );
  XOR2_X1 U695 ( .A(n657), .B(KEYINPUT80), .Z(n616) );
  XNOR2_X1 U696 ( .A(n617), .B(n616), .ZN(G145) );
  NAND2_X1 U697 ( .A1(n643), .A2(G75), .ZN(n619) );
  NAND2_X1 U698 ( .A1(G88), .A2(n640), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n619), .A2(n618), .ZN(n624) );
  NAND2_X1 U700 ( .A1(G62), .A2(n639), .ZN(n620) );
  XOR2_X1 U701 ( .A(KEYINPUT83), .B(n620), .Z(n622) );
  NAND2_X1 U702 ( .A1(n637), .A2(G50), .ZN(n621) );
  NAND2_X1 U703 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U704 ( .A1(n624), .A2(n623), .ZN(G166) );
  NAND2_X1 U705 ( .A1(G49), .A2(n637), .ZN(n626) );
  NAND2_X1 U706 ( .A1(G74), .A2(G651), .ZN(n625) );
  NAND2_X1 U707 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U708 ( .A1(n639), .A2(n627), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n628), .A2(G87), .ZN(n629) );
  NAND2_X1 U710 ( .A1(n630), .A2(n629), .ZN(G288) );
  AND2_X1 U711 ( .A1(n643), .A2(G72), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n637), .A2(G47), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G85), .A2(n640), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U715 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n639), .A2(G60), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(G290) );
  NAND2_X1 U718 ( .A1(G48), .A2(n637), .ZN(n638) );
  XNOR2_X1 U719 ( .A(n638), .B(KEYINPUT82), .ZN(n648) );
  NAND2_X1 U720 ( .A1(n639), .A2(G61), .ZN(n642) );
  NAND2_X1 U721 ( .A1(G86), .A2(n640), .ZN(n641) );
  NAND2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U723 ( .A1(n643), .A2(G73), .ZN(n644) );
  XOR2_X1 U724 ( .A(KEYINPUT2), .B(n644), .Z(n645) );
  NOR2_X1 U725 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U726 ( .A1(n648), .A2(n647), .ZN(G305) );
  XNOR2_X1 U727 ( .A(G166), .B(G299), .ZN(n653) );
  XNOR2_X1 U728 ( .A(KEYINPUT19), .B(G288), .ZN(n649) );
  XNOR2_X1 U729 ( .A(n649), .B(n657), .ZN(n650) );
  XNOR2_X1 U730 ( .A(n650), .B(G290), .ZN(n651) );
  XNOR2_X1 U731 ( .A(n651), .B(G305), .ZN(n652) );
  XNOR2_X1 U732 ( .A(n653), .B(n652), .ZN(n911) );
  XNOR2_X1 U733 ( .A(n911), .B(n654), .ZN(n655) );
  NOR2_X1 U734 ( .A1(n656), .A2(n655), .ZN(n659) );
  NOR2_X1 U735 ( .A1(G868), .A2(n657), .ZN(n658) );
  NOR2_X1 U736 ( .A1(n659), .A2(n658), .ZN(G295) );
  NAND2_X1 U737 ( .A1(G2084), .A2(G2078), .ZN(n661) );
  XOR2_X1 U738 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n660) );
  XNOR2_X1 U739 ( .A(n661), .B(n660), .ZN(n662) );
  NAND2_X1 U740 ( .A1(G2090), .A2(n662), .ZN(n663) );
  XNOR2_X1 U741 ( .A(KEYINPUT21), .B(n663), .ZN(n664) );
  NAND2_X1 U742 ( .A1(n664), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U743 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U744 ( .A1(G235), .A2(G236), .ZN(n665) );
  XOR2_X1 U745 ( .A(KEYINPUT86), .B(n665), .Z(n666) );
  NOR2_X1 U746 ( .A1(G238), .A2(n666), .ZN(n667) );
  NAND2_X1 U747 ( .A1(G57), .A2(n667), .ZN(n924) );
  NAND2_X1 U748 ( .A1(G567), .A2(n924), .ZN(n673) );
  NOR2_X1 U749 ( .A1(G220), .A2(G219), .ZN(n668) );
  XNOR2_X1 U750 ( .A(KEYINPUT22), .B(n668), .ZN(n669) );
  NAND2_X1 U751 ( .A1(n669), .A2(G96), .ZN(n670) );
  NOR2_X1 U752 ( .A1(n670), .A2(G218), .ZN(n671) );
  XNOR2_X1 U753 ( .A(n671), .B(KEYINPUT85), .ZN(n925) );
  NAND2_X1 U754 ( .A1(G2106), .A2(n925), .ZN(n672) );
  NAND2_X1 U755 ( .A1(n673), .A2(n672), .ZN(n832) );
  NAND2_X1 U756 ( .A1(G661), .A2(G483), .ZN(n674) );
  NOR2_X1 U757 ( .A1(n832), .A2(n674), .ZN(n675) );
  XOR2_X1 U758 ( .A(KEYINPUT87), .B(n675), .Z(n831) );
  NAND2_X1 U759 ( .A1(n831), .A2(G36), .ZN(G176) );
  INV_X1 U760 ( .A(G166), .ZN(G303) );
  INV_X1 U761 ( .A(KEYINPUT90), .ZN(n677) );
  NAND2_X1 U762 ( .A1(G40), .A2(G160), .ZN(n676) );
  XOR2_X1 U763 ( .A(n676), .B(KEYINPUT88), .Z(n779) );
  NOR2_X1 U764 ( .A1(G164), .A2(G1384), .ZN(n777) );
  NAND2_X2 U765 ( .A1(n779), .A2(n777), .ZN(n690) );
  XNOR2_X2 U766 ( .A(n690), .B(KEYINPUT64), .ZN(n739) );
  NOR2_X1 U767 ( .A1(n739), .A2(G2084), .ZN(n678) );
  NAND2_X1 U768 ( .A1(n677), .A2(n678), .ZN(n714) );
  INV_X1 U769 ( .A(n678), .ZN(n679) );
  NAND2_X1 U770 ( .A1(n679), .A2(KEYINPUT90), .ZN(n715) );
  AND2_X1 U771 ( .A1(n714), .A2(n715), .ZN(n680) );
  NAND2_X1 U772 ( .A1(n680), .A2(G8), .ZN(n732) );
  NAND2_X1 U773 ( .A1(n739), .A2(G8), .ZN(n773) );
  NOR2_X1 U774 ( .A1(G1966), .A2(n773), .ZN(n730) );
  INV_X1 U775 ( .A(n739), .ZN(n698) );
  NOR2_X1 U776 ( .A1(G1961), .A2(n698), .ZN(n682) );
  XOR2_X1 U777 ( .A(KEYINPUT25), .B(G2078), .Z(n932) );
  NOR2_X1 U778 ( .A1(n739), .A2(n932), .ZN(n681) );
  NOR2_X1 U779 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U780 ( .A(KEYINPUT91), .B(n683), .ZN(n722) );
  NAND2_X1 U781 ( .A1(n722), .A2(G171), .ZN(n733) );
  NAND2_X1 U782 ( .A1(G2072), .A2(n698), .ZN(n684) );
  XNOR2_X1 U783 ( .A(n684), .B(KEYINPUT27), .ZN(n686) );
  INV_X1 U784 ( .A(G1956), .ZN(n970) );
  NOR2_X1 U785 ( .A1(n698), .A2(n970), .ZN(n685) );
  NOR2_X1 U786 ( .A1(n686), .A2(n685), .ZN(n701) );
  NOR2_X1 U787 ( .A1(n701), .A2(n953), .ZN(n688) );
  XOR2_X1 U788 ( .A(KEYINPUT92), .B(KEYINPUT28), .Z(n687) );
  XNOR2_X1 U789 ( .A(n688), .B(n687), .ZN(n711) );
  INV_X1 U790 ( .A(KEYINPUT64), .ZN(n689) );
  XNOR2_X1 U791 ( .A(n690), .B(n689), .ZN(n691) );
  NAND2_X1 U792 ( .A1(n691), .A2(G1996), .ZN(n692) );
  XNOR2_X1 U793 ( .A(n692), .B(KEYINPUT26), .ZN(n694) );
  NAND2_X1 U794 ( .A1(n739), .A2(G1341), .ZN(n693) );
  NAND2_X1 U795 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U796 ( .A1(n695), .A2(n963), .ZN(n696) );
  XNOR2_X1 U797 ( .A(n696), .B(KEYINPUT65), .ZN(n706) );
  NOR2_X1 U798 ( .A1(n954), .A2(n706), .ZN(n697) );
  XNOR2_X1 U799 ( .A(n697), .B(KEYINPUT93), .ZN(n704) );
  NOR2_X1 U800 ( .A1(n698), .A2(G1348), .ZN(n700) );
  NOR2_X1 U801 ( .A1(G2067), .A2(n739), .ZN(n699) );
  NOR2_X1 U802 ( .A1(n700), .A2(n699), .ZN(n702) );
  NAND2_X1 U803 ( .A1(n701), .A2(n953), .ZN(n705) );
  AND2_X1 U804 ( .A1(n702), .A2(n705), .ZN(n703) );
  NAND2_X1 U805 ( .A1(n704), .A2(n703), .ZN(n709) );
  AND2_X1 U806 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U807 ( .A1(n954), .A2(n707), .ZN(n708) );
  AND2_X1 U808 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U809 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U810 ( .A(n712), .B(KEYINPUT29), .ZN(n713) );
  INV_X1 U811 ( .A(n713), .ZN(n735) );
  NAND2_X1 U812 ( .A1(n733), .A2(n735), .ZN(n727) );
  INV_X1 U813 ( .A(KEYINPUT31), .ZN(n726) );
  NAND2_X1 U814 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U815 ( .A1(G8), .A2(n716), .ZN(n717) );
  NOR2_X1 U816 ( .A1(n730), .A2(n717), .ZN(n720) );
  INV_X1 U817 ( .A(KEYINPUT94), .ZN(n718) );
  NOR2_X1 U818 ( .A1(n721), .A2(G168), .ZN(n724) );
  NOR2_X1 U819 ( .A1(G171), .A2(n722), .ZN(n723) );
  NOR2_X1 U820 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U821 ( .A(n726), .B(n725), .ZN(n736) );
  NAND2_X1 U822 ( .A1(n727), .A2(n736), .ZN(n728) );
  XNOR2_X1 U823 ( .A(KEYINPUT95), .B(n728), .ZN(n729) );
  NOR2_X1 U824 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U825 ( .A1(n732), .A2(n731), .ZN(n751) );
  AND2_X1 U826 ( .A1(n733), .A2(G286), .ZN(n734) );
  NAND2_X1 U827 ( .A1(n735), .A2(n734), .ZN(n747) );
  INV_X1 U828 ( .A(G286), .ZN(n737) );
  OR2_X1 U829 ( .A1(n737), .A2(n736), .ZN(n745) );
  NOR2_X1 U830 ( .A1(G1971), .A2(n773), .ZN(n738) );
  XNOR2_X1 U831 ( .A(n738), .B(KEYINPUT96), .ZN(n741) );
  NOR2_X1 U832 ( .A1(n739), .A2(G2090), .ZN(n740) );
  NOR2_X1 U833 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U834 ( .A1(n742), .A2(G303), .ZN(n743) );
  XOR2_X1 U835 ( .A(KEYINPUT97), .B(n743), .Z(n744) );
  NAND2_X1 U836 ( .A1(n748), .A2(G8), .ZN(n749) );
  XNOR2_X1 U837 ( .A(n749), .B(KEYINPUT32), .ZN(n750) );
  NAND2_X1 U838 ( .A1(n751), .A2(n750), .ZN(n758) );
  NOR2_X1 U839 ( .A1(G2090), .A2(G303), .ZN(n752) );
  NAND2_X1 U840 ( .A1(G8), .A2(n752), .ZN(n753) );
  NAND2_X1 U841 ( .A1(n758), .A2(n753), .ZN(n754) );
  NAND2_X1 U842 ( .A1(n754), .A2(n773), .ZN(n769) );
  NOR2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n760) );
  NOR2_X1 U844 ( .A1(G1971), .A2(G303), .ZN(n755) );
  NOR2_X1 U845 ( .A1(n760), .A2(n755), .ZN(n958) );
  INV_X1 U846 ( .A(KEYINPUT33), .ZN(n756) );
  AND2_X1 U847 ( .A1(n958), .A2(n756), .ZN(n757) );
  NAND2_X1 U848 ( .A1(n758), .A2(n757), .ZN(n767) );
  NAND2_X1 U849 ( .A1(G1976), .A2(G288), .ZN(n957) );
  INV_X1 U850 ( .A(n957), .ZN(n759) );
  OR2_X1 U851 ( .A1(KEYINPUT33), .A2(n514), .ZN(n763) );
  NAND2_X1 U852 ( .A1(n760), .A2(KEYINPUT33), .ZN(n761) );
  OR2_X1 U853 ( .A1(n773), .A2(n761), .ZN(n762) );
  NAND2_X1 U854 ( .A1(n763), .A2(n762), .ZN(n765) );
  XOR2_X1 U855 ( .A(G1981), .B(G305), .Z(n945) );
  INV_X1 U856 ( .A(n945), .ZN(n764) );
  NOR2_X1 U857 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U858 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U859 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U860 ( .A(n770), .B(KEYINPUT98), .ZN(n775) );
  NOR2_X1 U861 ( .A1(G1981), .A2(G305), .ZN(n771) );
  XOR2_X1 U862 ( .A(n771), .B(KEYINPUT24), .Z(n772) );
  NOR2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X2 U864 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U865 ( .A(n776), .B(KEYINPUT99), .ZN(n810) );
  INV_X1 U866 ( .A(n777), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n805) );
  INV_X1 U868 ( .A(n805), .ZN(n822) );
  XNOR2_X1 U869 ( .A(G2067), .B(KEYINPUT37), .ZN(n820) );
  NAND2_X1 U870 ( .A1(G104), .A2(n894), .ZN(n781) );
  NAND2_X1 U871 ( .A1(G140), .A2(n895), .ZN(n780) );
  NAND2_X1 U872 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U873 ( .A(KEYINPUT34), .B(n782), .ZN(n788) );
  NAND2_X1 U874 ( .A1(G128), .A2(n901), .ZN(n784) );
  NAND2_X1 U875 ( .A1(G116), .A2(n899), .ZN(n783) );
  NAND2_X1 U876 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U877 ( .A(KEYINPUT35), .B(n785), .ZN(n786) );
  XNOR2_X1 U878 ( .A(KEYINPUT89), .B(n786), .ZN(n787) );
  NOR2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U880 ( .A(KEYINPUT36), .B(n789), .ZN(n907) );
  NOR2_X1 U881 ( .A1(n820), .A2(n907), .ZN(n1005) );
  NAND2_X1 U882 ( .A1(n822), .A2(n1005), .ZN(n818) );
  NAND2_X1 U883 ( .A1(G119), .A2(n901), .ZN(n791) );
  NAND2_X1 U884 ( .A1(G131), .A2(n895), .ZN(n790) );
  NAND2_X1 U885 ( .A1(n791), .A2(n790), .ZN(n795) );
  NAND2_X1 U886 ( .A1(G95), .A2(n894), .ZN(n793) );
  NAND2_X1 U887 ( .A1(G107), .A2(n899), .ZN(n792) );
  NAND2_X1 U888 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U889 ( .A1(n795), .A2(n794), .ZN(n889) );
  INV_X1 U890 ( .A(G1991), .ZN(n811) );
  NOR2_X1 U891 ( .A1(n889), .A2(n811), .ZN(n804) );
  NAND2_X1 U892 ( .A1(G129), .A2(n901), .ZN(n797) );
  NAND2_X1 U893 ( .A1(G141), .A2(n895), .ZN(n796) );
  NAND2_X1 U894 ( .A1(n797), .A2(n796), .ZN(n800) );
  NAND2_X1 U895 ( .A1(n894), .A2(G105), .ZN(n798) );
  XOR2_X1 U896 ( .A(KEYINPUT38), .B(n798), .Z(n799) );
  NOR2_X1 U897 ( .A1(n800), .A2(n799), .ZN(n802) );
  NAND2_X1 U898 ( .A1(n899), .A2(G117), .ZN(n801) );
  NAND2_X1 U899 ( .A1(n802), .A2(n801), .ZN(n882) );
  AND2_X1 U900 ( .A1(G1996), .A2(n882), .ZN(n803) );
  NOR2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n1015) );
  NOR2_X1 U902 ( .A1(n1015), .A2(n805), .ZN(n814) );
  INV_X1 U903 ( .A(n814), .ZN(n806) );
  AND2_X1 U904 ( .A1(n818), .A2(n806), .ZN(n808) );
  XNOR2_X1 U905 ( .A(G1986), .B(G290), .ZN(n952) );
  NAND2_X1 U906 ( .A1(n952), .A2(n822), .ZN(n807) );
  AND2_X1 U907 ( .A1(n808), .A2(n807), .ZN(n809) );
  NAND2_X1 U908 ( .A1(n810), .A2(n809), .ZN(n825) );
  NOR2_X1 U909 ( .A1(G1996), .A2(n882), .ZN(n1010) );
  NOR2_X1 U910 ( .A1(G1986), .A2(G290), .ZN(n812) );
  AND2_X1 U911 ( .A1(n811), .A2(n889), .ZN(n1003) );
  NOR2_X1 U912 ( .A1(n812), .A2(n1003), .ZN(n813) );
  NOR2_X1 U913 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U914 ( .A(n815), .B(KEYINPUT100), .ZN(n816) );
  NOR2_X1 U915 ( .A1(n1010), .A2(n816), .ZN(n817) );
  XNOR2_X1 U916 ( .A(n817), .B(KEYINPUT39), .ZN(n819) );
  NAND2_X1 U917 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U918 ( .A1(n820), .A2(n907), .ZN(n1014) );
  NAND2_X1 U919 ( .A1(n821), .A2(n1014), .ZN(n823) );
  NAND2_X1 U920 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U921 ( .A1(n825), .A2(n824), .ZN(n827) );
  XOR2_X1 U922 ( .A(KEYINPUT40), .B(KEYINPUT101), .Z(n826) );
  XNOR2_X1 U923 ( .A(n827), .B(n826), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n828), .ZN(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n829) );
  NAND2_X1 U926 ( .A1(G661), .A2(n829), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n830) );
  NAND2_X1 U928 ( .A1(n831), .A2(n830), .ZN(G188) );
  XNOR2_X1 U929 ( .A(KEYINPUT105), .B(n832), .ZN(G319) );
  XNOR2_X1 U930 ( .A(G2427), .B(G2451), .ZN(n842) );
  XOR2_X1 U931 ( .A(KEYINPUT103), .B(G2443), .Z(n834) );
  XNOR2_X1 U932 ( .A(G2435), .B(G2438), .ZN(n833) );
  XNOR2_X1 U933 ( .A(n834), .B(n833), .ZN(n838) );
  XOR2_X1 U934 ( .A(G2454), .B(G2430), .Z(n836) );
  XNOR2_X1 U935 ( .A(G1348), .B(G1341), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U937 ( .A(n838), .B(n837), .Z(n840) );
  XNOR2_X1 U938 ( .A(KEYINPUT102), .B(G2446), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(n843) );
  NAND2_X1 U941 ( .A1(n843), .A2(G14), .ZN(n844) );
  XOR2_X1 U942 ( .A(KEYINPUT104), .B(n844), .Z(G401) );
  XOR2_X1 U943 ( .A(KEYINPUT109), .B(G1956), .Z(n846) );
  XNOR2_X1 U944 ( .A(G1981), .B(G1966), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U946 ( .A(n847), .B(KEYINPUT41), .Z(n849) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1991), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U949 ( .A(G1976), .B(G1971), .Z(n851) );
  XNOR2_X1 U950 ( .A(G1986), .B(G1961), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U952 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U953 ( .A(KEYINPUT108), .B(G2474), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(G229) );
  XOR2_X1 U955 ( .A(G2100), .B(KEYINPUT107), .Z(n857) );
  XNOR2_X1 U956 ( .A(G2678), .B(KEYINPUT43), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U958 ( .A(KEYINPUT42), .B(G2072), .Z(n859) );
  XNOR2_X1 U959 ( .A(G2067), .B(G2090), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U961 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U962 ( .A(KEYINPUT106), .B(G2096), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(n865) );
  XOR2_X1 U964 ( .A(G2084), .B(G2078), .Z(n864) );
  XNOR2_X1 U965 ( .A(n865), .B(n864), .ZN(G227) );
  NAND2_X1 U966 ( .A1(G124), .A2(n901), .ZN(n866) );
  XNOR2_X1 U967 ( .A(n866), .B(KEYINPUT44), .ZN(n867) );
  XNOR2_X1 U968 ( .A(n867), .B(KEYINPUT110), .ZN(n869) );
  NAND2_X1 U969 ( .A1(G112), .A2(n899), .ZN(n868) );
  NAND2_X1 U970 ( .A1(n869), .A2(n868), .ZN(n873) );
  NAND2_X1 U971 ( .A1(G100), .A2(n894), .ZN(n871) );
  NAND2_X1 U972 ( .A1(G136), .A2(n895), .ZN(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U974 ( .A1(n873), .A2(n872), .ZN(G162) );
  NAND2_X1 U975 ( .A1(G130), .A2(n901), .ZN(n875) );
  NAND2_X1 U976 ( .A1(G118), .A2(n899), .ZN(n874) );
  NAND2_X1 U977 ( .A1(n875), .A2(n874), .ZN(n881) );
  NAND2_X1 U978 ( .A1(n894), .A2(G106), .ZN(n876) );
  XOR2_X1 U979 ( .A(KEYINPUT111), .B(n876), .Z(n878) );
  NAND2_X1 U980 ( .A1(n895), .A2(G142), .ZN(n877) );
  NAND2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U982 ( .A(KEYINPUT45), .B(n879), .Z(n880) );
  NOR2_X1 U983 ( .A1(n881), .A2(n880), .ZN(n893) );
  XOR2_X1 U984 ( .A(G162), .B(n1004), .Z(n884) );
  XOR2_X1 U985 ( .A(G164), .B(n882), .Z(n883) );
  XNOR2_X1 U986 ( .A(n884), .B(n883), .ZN(n888) );
  XOR2_X1 U987 ( .A(KEYINPUT115), .B(KEYINPUT112), .Z(n886) );
  XNOR2_X1 U988 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n885) );
  XNOR2_X1 U989 ( .A(n886), .B(n885), .ZN(n887) );
  XOR2_X1 U990 ( .A(n888), .B(n887), .Z(n891) );
  XNOR2_X1 U991 ( .A(G160), .B(n889), .ZN(n890) );
  XNOR2_X1 U992 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U993 ( .A(n893), .B(n892), .ZN(n909) );
  NAND2_X1 U994 ( .A1(G103), .A2(n894), .ZN(n897) );
  NAND2_X1 U995 ( .A1(G139), .A2(n895), .ZN(n896) );
  NAND2_X1 U996 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U997 ( .A(KEYINPUT113), .B(n898), .Z(n906) );
  NAND2_X1 U998 ( .A1(n899), .A2(G115), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n900), .B(KEYINPUT114), .ZN(n903) );
  NAND2_X1 U1000 ( .A1(G127), .A2(n901), .ZN(n902) );
  NAND2_X1 U1001 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1002 ( .A(KEYINPUT47), .B(n904), .Z(n905) );
  NOR2_X1 U1003 ( .A1(n906), .A2(n905), .ZN(n998) );
  XNOR2_X1 U1004 ( .A(n907), .B(n998), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n910), .ZN(G395) );
  XNOR2_X1 U1007 ( .A(G286), .B(n911), .ZN(n914) );
  XNOR2_X1 U1008 ( .A(KEYINPUT116), .B(G301), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(n912), .B(n954), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n915) );
  XOR2_X1 U1011 ( .A(n915), .B(n963), .Z(n916) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n916), .ZN(G397) );
  INV_X1 U1013 ( .A(G401), .ZN(n917) );
  NAND2_X1 U1014 ( .A1(G319), .A2(n917), .ZN(n921) );
  NOR2_X1 U1015 ( .A1(G229), .A2(G227), .ZN(n918) );
  XOR2_X1 U1016 ( .A(KEYINPUT49), .B(n918), .Z(n919) );
  XNOR2_X1 U1017 ( .A(n919), .B(KEYINPUT117), .ZN(n920) );
  NOR2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(G395), .A2(G397), .ZN(n922) );
  NAND2_X1 U1020 ( .A1(n923), .A2(n922), .ZN(G225) );
  XOR2_X1 U1021 ( .A(KEYINPUT118), .B(G225), .Z(G308) );
  INV_X1 U1023 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(G325) );
  INV_X1 U1025 ( .A(G325), .ZN(G261) );
  INV_X1 U1026 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1027 ( .A(G2072), .B(G33), .Z(n926) );
  NAND2_X1 U1028 ( .A1(n926), .A2(G28), .ZN(n929) );
  XOR2_X1 U1029 ( .A(G25), .B(G1991), .Z(n927) );
  XNOR2_X1 U1030 ( .A(KEYINPUT123), .B(n927), .ZN(n928) );
  NOR2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n936) );
  XOR2_X1 U1032 ( .A(G2067), .B(G26), .Z(n931) );
  XOR2_X1 U1033 ( .A(G1996), .B(G32), .Z(n930) );
  NAND2_X1 U1034 ( .A1(n931), .A2(n930), .ZN(n934) );
  XNOR2_X1 U1035 ( .A(G27), .B(n932), .ZN(n933) );
  NOR2_X1 U1036 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1038 ( .A(KEYINPUT53), .B(n937), .ZN(n941) );
  XOR2_X1 U1039 ( .A(KEYINPUT124), .B(G34), .Z(n939) );
  XNOR2_X1 U1040 ( .A(G2084), .B(KEYINPUT54), .ZN(n938) );
  XNOR2_X1 U1041 ( .A(n939), .B(n938), .ZN(n940) );
  NAND2_X1 U1042 ( .A1(n941), .A2(n940), .ZN(n943) );
  XNOR2_X1 U1043 ( .A(G35), .B(G2090), .ZN(n942) );
  NOR2_X1 U1044 ( .A1(n943), .A2(n942), .ZN(n1030) );
  NAND2_X1 U1045 ( .A1(KEYINPUT55), .A2(n1030), .ZN(n944) );
  NAND2_X1 U1046 ( .A1(G11), .A2(n944), .ZN(n1029) );
  XNOR2_X1 U1047 ( .A(G16), .B(KEYINPUT56), .ZN(n969) );
  XNOR2_X1 U1048 ( .A(G1966), .B(G168), .ZN(n946) );
  NAND2_X1 U1049 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1050 ( .A(n947), .B(KEYINPUT57), .ZN(n948) );
  XOR2_X1 U1051 ( .A(KEYINPUT125), .B(n948), .Z(n967) );
  XNOR2_X1 U1052 ( .A(G1961), .B(G171), .ZN(n950) );
  NAND2_X1 U1053 ( .A1(G1971), .A2(G303), .ZN(n949) );
  NAND2_X1 U1054 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1055 ( .A1(n952), .A2(n951), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(n953), .B(G1956), .ZN(n956) );
  XOR2_X1 U1057 ( .A(G1348), .B(n954), .Z(n955) );
  NAND2_X1 U1058 ( .A1(n956), .A2(n955), .ZN(n960) );
  NAND2_X1 U1059 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1060 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1061 ( .A1(n962), .A2(n961), .ZN(n965) );
  XNOR2_X1 U1062 ( .A(G1341), .B(n963), .ZN(n964) );
  NOR2_X1 U1063 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1065 ( .A1(n969), .A2(n968), .ZN(n995) );
  INV_X1 U1066 ( .A(G16), .ZN(n993) );
  XNOR2_X1 U1067 ( .A(G20), .B(n970), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(G1981), .B(G6), .ZN(n972) );
  XNOR2_X1 U1069 ( .A(G1341), .B(G19), .ZN(n971) );
  NOR2_X1 U1070 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n977) );
  XOR2_X1 U1072 ( .A(KEYINPUT59), .B(G1348), .Z(n975) );
  XNOR2_X1 U1073 ( .A(G4), .B(n975), .ZN(n976) );
  NOR2_X1 U1074 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1075 ( .A(KEYINPUT60), .B(n978), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(G1966), .B(G21), .ZN(n980) );
  XNOR2_X1 U1077 ( .A(G5), .B(G1961), .ZN(n979) );
  NOR2_X1 U1078 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1079 ( .A1(n982), .A2(n981), .ZN(n989) );
  XNOR2_X1 U1080 ( .A(G1971), .B(G22), .ZN(n984) );
  XNOR2_X1 U1081 ( .A(G23), .B(G1976), .ZN(n983) );
  NOR2_X1 U1082 ( .A1(n984), .A2(n983), .ZN(n986) );
  XOR2_X1 U1083 ( .A(G1986), .B(G24), .Z(n985) );
  NAND2_X1 U1084 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1085 ( .A(KEYINPUT58), .B(n987), .ZN(n988) );
  NOR2_X1 U1086 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1087 ( .A(n990), .B(KEYINPUT61), .ZN(n991) );
  XNOR2_X1 U1088 ( .A(n991), .B(KEYINPUT126), .ZN(n992) );
  NAND2_X1 U1089 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1090 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1091 ( .A(KEYINPUT127), .B(n996), .ZN(n1027) );
  XNOR2_X1 U1092 ( .A(G164), .B(G2078), .ZN(n997) );
  XNOR2_X1 U1093 ( .A(n997), .B(KEYINPUT121), .ZN(n1000) );
  XOR2_X1 U1094 ( .A(G2072), .B(n998), .Z(n999) );
  NOR2_X1 U1095 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1096 ( .A(KEYINPUT50), .B(n1001), .Z(n1020) );
  XOR2_X1 U1097 ( .A(G160), .B(G2084), .Z(n1002) );
  NOR2_X1 U1098 ( .A1(n1003), .A2(n1002), .ZN(n1007) );
  NOR2_X1 U1099 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1100 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1101 ( .A(n1008), .B(KEYINPUT119), .ZN(n1013) );
  XOR2_X1 U1102 ( .A(G2090), .B(G162), .Z(n1009) );
  NOR2_X1 U1103 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1104 ( .A(KEYINPUT51), .B(n1011), .Z(n1012) );
  NAND2_X1 U1105 ( .A1(n1013), .A2(n1012), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1108 ( .A(KEYINPUT120), .B(n1018), .Z(n1019) );
  NOR2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1110 ( .A(KEYINPUT122), .B(n1021), .ZN(n1022) );
  XNOR2_X1 U1111 ( .A(n1022), .B(KEYINPUT52), .ZN(n1024) );
  INV_X1 U1112 ( .A(KEYINPUT55), .ZN(n1023) );
  NAND2_X1 U1113 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1114 ( .A1(G29), .A2(n1025), .ZN(n1026) );
  NAND2_X1 U1115 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1116 ( .A1(n1029), .A2(n1028), .ZN(n1034) );
  INV_X1 U1117 ( .A(n1030), .ZN(n1032) );
  NOR2_X1 U1118 ( .A1(G29), .A2(KEYINPUT55), .ZN(n1031) );
  NAND2_X1 U1119 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1120 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XOR2_X1 U1121 ( .A(KEYINPUT62), .B(n1035), .Z(G311) );
  INV_X1 U1122 ( .A(G311), .ZN(G150) );
endmodule

