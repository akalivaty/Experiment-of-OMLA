//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:34 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G50), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  OAI21_X1  g0006(.A(KEYINPUT64), .B1(new_n202), .B2(G50), .ZN(new_n207));
  AND3_X1   g0007(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n217), .A2(G50), .A3(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(new_n211), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(KEYINPUT66), .B(G244), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n224), .A2(new_n206), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G58), .A2(G232), .ZN(new_n229));
  NAND4_X1  g0029(.A1(new_n226), .A2(new_n227), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n213), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n216), .B(new_n223), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G264), .B(G270), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  INV_X1    g0044(.A(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(G68), .ZN(new_n246));
  INV_X1    g0046(.A(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n244), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n221), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT8), .ZN(new_n255));
  INV_X1    g0055(.A(G58), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n255), .B1(new_n256), .B2(KEYINPUT70), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT70), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(KEYINPUT8), .A3(G58), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n211), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT71), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  OR3_X1    g0063(.A1(new_n263), .A2(KEYINPUT71), .A3(G20), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n260), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G150), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n265), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n211), .B1(new_n205), .B2(new_n207), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n254), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n210), .A2(G13), .A3(G20), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(G50), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n254), .B1(new_n210), .B2(G20), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n273), .B1(new_n274), .B2(G50), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT9), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n271), .A2(KEYINPUT9), .A3(new_n275), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT10), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT67), .A2(G41), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT67), .A2(G41), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G274), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(G1), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(G1), .A3(G13), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G41), .ZN(new_n294));
  AOI21_X1  g0094(.A(G1), .B1(new_n294), .B2(new_n286), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n290), .B1(G226), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g0097(.A(KEYINPUT3), .B(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G1698), .ZN(new_n299));
  INV_X1    g0099(.A(G223), .ZN(new_n300));
  OAI22_X1  g0100(.A1(new_n299), .A2(new_n300), .B1(new_n206), .B2(new_n298), .ZN(new_n301));
  OR2_X1    g0101(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT3), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G33), .ZN(new_n305));
  NAND2_X1  g0105(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n306));
  NAND4_X1  g0106(.A1(new_n302), .A2(new_n303), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G222), .ZN(new_n308));
  OR3_X1    g0108(.A1(new_n307), .A2(KEYINPUT69), .A3(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT69), .B1(new_n307), .B2(new_n308), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n301), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n297), .B1(new_n311), .B2(new_n292), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G200), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n297), .B(G190), .C1(new_n311), .C2(new_n292), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n280), .A2(new_n281), .A3(new_n313), .A4(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n278), .A2(new_n314), .A3(new_n279), .ZN(new_n316));
  INV_X1    g0116(.A(new_n313), .ZN(new_n317));
  OAI21_X1  g0117(.A(KEYINPUT10), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n276), .ZN(new_n320));
  INV_X1    g0120(.A(G169), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n320), .B1(new_n321), .B2(new_n312), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(G179), .B2(new_n312), .ZN(new_n323));
  INV_X1    g0123(.A(new_n224), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n290), .B1(new_n324), .B2(new_n296), .ZN(new_n325));
  INV_X1    g0125(.A(G238), .ZN(new_n326));
  INV_X1    g0126(.A(G107), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n299), .A2(new_n326), .B1(new_n327), .B2(new_n298), .ZN(new_n328));
  INV_X1    g0128(.A(new_n306), .ZN(new_n329));
  NOR2_X1   g0129(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n331), .A2(new_n298), .A3(G232), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n293), .B1(new_n328), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n325), .A2(G190), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT72), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n334), .B(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(G20), .A2(G77), .ZN(new_n337));
  XNOR2_X1  g0137(.A(KEYINPUT15), .B(G87), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT8), .B(G58), .ZN(new_n339));
  OAI221_X1 g0139(.A(new_n337), .B1(new_n338), .B2(new_n261), .C1(new_n268), .C2(new_n339), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n340), .A2(new_n254), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n274), .A2(G77), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(G77), .B2(new_n272), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n325), .A2(new_n333), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n345), .B1(G200), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n336), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G179), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n325), .A2(new_n349), .A3(new_n333), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT73), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n350), .B(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n344), .B1(new_n321), .B2(new_n346), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  AND4_X1   g0154(.A1(new_n319), .A2(new_n323), .A3(new_n348), .A4(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n254), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT16), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G58), .A2(G68), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT76), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n202), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(G20), .B1(G159), .B2(new_n267), .ZN(new_n361));
  AOI21_X1  g0161(.A(G20), .B1(new_n303), .B2(new_n305), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT77), .B1(new_n362), .B2(KEYINPUT7), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT77), .ZN(new_n364));
  INV_X1    g0164(.A(KEYINPUT7), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n364), .B(new_n365), .C1(new_n298), .C2(G20), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n305), .A2(KEYINPUT78), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n211), .A2(KEYINPUT7), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n298), .A2(KEYINPUT78), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n363), .A2(new_n366), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n357), .B(new_n361), .C1(new_n371), .C2(new_n247), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n267), .A2(G159), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT76), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n358), .B(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n375), .A2(new_n201), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n373), .B1(new_n376), .B2(new_n211), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n362), .A2(KEYINPUT7), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n365), .B1(new_n298), .B2(G20), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n247), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT16), .B1(new_n377), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n356), .B1(new_n372), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n272), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n210), .A2(G20), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n260), .A2(new_n384), .ZN(new_n385));
  AOI211_X1 g0185(.A(new_n383), .B(new_n254), .C1(new_n385), .C2(KEYINPUT79), .ZN(new_n386));
  OR2_X1    g0186(.A1(new_n385), .A2(KEYINPUT79), .ZN(new_n387));
  INV_X1    g0187(.A(new_n260), .ZN(new_n388));
  AOI22_X1  g0188(.A1(new_n386), .A2(new_n387), .B1(new_n383), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n382), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n303), .A2(new_n305), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n302), .A2(G223), .A3(new_n306), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G226), .A2(G1698), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(G87), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n263), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n293), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n296), .A2(G232), .B1(new_n287), .B2(new_n289), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G190), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n402), .B1(G200), .B2(new_n400), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n391), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT17), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n391), .A2(KEYINPUT17), .A3(new_n403), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n321), .B1(new_n398), .B2(new_n399), .ZN(new_n409));
  INV_X1    g0209(.A(new_n400), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n409), .B1(new_n410), .B2(G179), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n357), .B(new_n373), .C1(new_n376), .C2(new_n211), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n363), .A2(new_n366), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n369), .A2(new_n370), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n412), .B1(new_n415), .B2(G68), .ZN(new_n416));
  INV_X1    g0216(.A(new_n380), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n357), .B1(new_n417), .B2(new_n361), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n254), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n411), .B1(new_n419), .B2(new_n389), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT81), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n420), .A2(new_n421), .A3(KEYINPUT18), .ZN(new_n422));
  INV_X1    g0222(.A(new_n409), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n349), .B2(new_n400), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n424), .B1(new_n382), .B2(new_n390), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT81), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n424), .B(KEYINPUT18), .C1(new_n382), .C2(new_n390), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT80), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n419), .A2(new_n389), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT80), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n431), .A2(new_n432), .A3(KEYINPUT18), .A4(new_n424), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n408), .B1(new_n428), .B2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n303), .A2(new_n305), .A3(G232), .A4(G1698), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G97), .ZN(new_n437));
  INV_X1    g0237(.A(G226), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n436), .B(new_n437), .C1(new_n307), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n293), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n296), .A2(G238), .B1(new_n287), .B2(new_n289), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT13), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n442), .B1(new_n440), .B2(new_n441), .ZN(new_n445));
  OAI21_X1  g0245(.A(G169), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT14), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT14), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n448), .B(G169), .C1(new_n444), .C2(new_n445), .ZN(new_n449));
  INV_X1    g0249(.A(new_n445), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n450), .A2(G179), .A3(new_n443), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n447), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n383), .A2(new_n247), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT12), .ZN(new_n454));
  XNOR2_X1  g0254(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n264), .A2(new_n262), .A3(G77), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n267), .A2(G50), .B1(G20), .B2(new_n247), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n356), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n455), .B1(new_n458), .B2(KEYINPUT11), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n458), .A2(KEYINPUT11), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n274), .A2(KEYINPUT74), .A3(G68), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT74), .B1(new_n274), .B2(G68), .ZN(new_n462));
  OR2_X1    g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n459), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT75), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n459), .A2(KEYINPUT75), .A3(new_n463), .A4(new_n460), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n452), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n466), .A2(new_n467), .ZN(new_n470));
  OAI21_X1  g0270(.A(G200), .B1(new_n444), .B2(new_n445), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n450), .A2(G190), .A3(new_n443), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n355), .A2(new_n435), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n327), .A2(KEYINPUT6), .A3(G97), .ZN(new_n477));
  INV_X1    g0277(.A(G97), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(new_n327), .ZN(new_n479));
  NOR2_X1   g0279(.A1(G97), .A2(G107), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n477), .B1(new_n481), .B2(KEYINPUT6), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n482), .A2(G20), .B1(G77), .B2(new_n267), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n371), .B2(new_n327), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n254), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n383), .A2(new_n478), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n210), .A2(G33), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n356), .A2(new_n272), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n486), .B1(new_n488), .B2(new_n478), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n485), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT4), .ZN(new_n492));
  INV_X1    g0292(.A(G244), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n492), .B1(new_n307), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(G33), .A2(G283), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n331), .A2(new_n298), .A3(KEYINPUT4), .A4(G244), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n298), .A2(G250), .A3(G1698), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n494), .A2(new_n495), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n293), .ZN(new_n499));
  OR2_X1    g0299(.A1(KEYINPUT67), .A2(G41), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT5), .B1(new_n500), .B2(new_n282), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT5), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n210), .B(G45), .C1(new_n502), .C2(G41), .ZN(new_n503));
  OAI211_X1 g0303(.A(G257), .B(new_n292), .C1(new_n501), .C2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n502), .B1(new_n283), .B2(new_n284), .ZN(new_n505));
  INV_X1    g0305(.A(new_n503), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n505), .A2(new_n506), .A3(G274), .A4(new_n292), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(G169), .B1(new_n499), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n508), .B1(new_n498), .B2(new_n293), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n349), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n491), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n489), .B1(new_n484), .B2(new_n254), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n499), .A2(G190), .A3(new_n509), .ZN(new_n516));
  INV_X1    g0316(.A(G200), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n515), .B(new_n516), .C1(new_n517), .C2(new_n512), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n303), .A2(new_n305), .A3(G257), .A4(G1698), .ZN(new_n519));
  NAND2_X1  g0319(.A1(G33), .A2(G294), .ZN(new_n520));
  INV_X1    g0320(.A(G250), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n519), .B(new_n520), .C1(new_n307), .C2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n293), .B1(new_n505), .B2(new_n506), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n522), .A2(new_n293), .B1(new_n523), .B2(G264), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n507), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n321), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n524), .A2(new_n349), .A3(new_n507), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n303), .A2(new_n305), .A3(new_n211), .A4(G87), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT87), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(new_n529), .A3(KEYINPUT22), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n529), .A2(KEYINPUT22), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n298), .A2(new_n211), .A3(G87), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G116), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(G20), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT23), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(new_n211), .B2(G107), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n327), .A2(KEYINPUT23), .A3(G20), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n533), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(KEYINPUT24), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT24), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n533), .A2(new_n542), .A3(new_n539), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n356), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT25), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(new_n272), .B2(G107), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n272), .A2(new_n545), .A3(G107), .ZN(new_n548));
  OAI22_X1  g0348(.A1(new_n488), .A2(new_n327), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n526), .B(new_n527), .C1(new_n544), .C2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n543), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n542), .B1(new_n533), .B2(new_n539), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n254), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n525), .A2(G200), .ZN(new_n554));
  INV_X1    g0354(.A(new_n549), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n524), .A2(G190), .A3(new_n507), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n553), .A2(new_n554), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n514), .A2(new_n518), .A3(new_n550), .A4(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n272), .A2(G116), .ZN(new_n559));
  INV_X1    g0359(.A(new_n488), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n559), .B1(new_n560), .B2(G116), .ZN(new_n561));
  AOI21_X1  g0361(.A(G20), .B1(G33), .B2(G283), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n263), .A2(G97), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT86), .ZN(new_n565));
  XNOR2_X1  g0365(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(G116), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n253), .A2(new_n221), .B1(G20), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT20), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n564), .A2(new_n565), .ZN(new_n570));
  AOI21_X1  g0370(.A(KEYINPUT86), .B1(new_n562), .B2(new_n563), .ZN(new_n571));
  OAI211_X1 g0371(.A(KEYINPUT20), .B(new_n568), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n561), .B1(new_n569), .B2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n331), .A2(new_n298), .A3(G257), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n298), .A2(G264), .A3(G1698), .ZN(new_n577));
  INV_X1    g0377(.A(G303), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n576), .B(new_n577), .C1(new_n578), .C2(new_n298), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n293), .ZN(new_n580));
  OAI211_X1 g0380(.A(G270), .B(new_n292), .C1(new_n501), .C2(new_n503), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n581), .A2(new_n507), .A3(KEYINPUT85), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT85), .B1(new_n581), .B2(new_n507), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n580), .B(G190), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n581), .A2(new_n507), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT85), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n581), .A2(new_n507), .A3(KEYINPUT85), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n587), .A2(new_n588), .B1(new_n293), .B2(new_n579), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n575), .B(new_n584), .C1(new_n589), .C2(new_n517), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n580), .B1(new_n582), .B2(new_n583), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n591), .A2(new_n574), .A3(G169), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT21), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n591), .A2(new_n574), .A3(KEYINPUT21), .A4(G169), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n589), .A2(G179), .A3(new_n574), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n590), .A2(new_n594), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n338), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n598), .A2(new_n272), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n488), .A2(new_n338), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n303), .A2(new_n305), .A3(new_n211), .A4(G68), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT19), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n261), .B2(new_n478), .ZN(new_n603));
  NAND3_X1  g0403(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n211), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n396), .A2(new_n478), .A3(new_n327), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n605), .A2(KEYINPUT83), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(KEYINPUT83), .B1(new_n605), .B2(new_n606), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n601), .B(new_n603), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT84), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n356), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n601), .A2(new_n603), .ZN(new_n612));
  INV_X1    g0412(.A(new_n608), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n605), .A2(KEYINPUT83), .A3(new_n606), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT84), .ZN(new_n616));
  AOI211_X1 g0416(.A(new_n599), .B(new_n600), .C1(new_n611), .C2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n307), .A2(new_n326), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n303), .A2(new_n305), .A3(G244), .A4(G1698), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n534), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n293), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n521), .B1(new_n210), .B2(G45), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n292), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT82), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n622), .A2(new_n292), .A3(KEYINPUT82), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n210), .A2(G45), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n625), .A2(new_n626), .B1(G274), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n621), .A2(new_n629), .A3(new_n349), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(G274), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n622), .A2(new_n292), .A3(KEYINPUT82), .ZN(new_n632));
  AOI21_X1  g0432(.A(KEYINPUT82), .B1(new_n622), .B2(new_n292), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n331), .A2(new_n298), .A3(G238), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n635), .A2(new_n619), .A3(new_n534), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n634), .B1(new_n293), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n630), .B1(new_n637), .B2(G169), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n560), .A2(G87), .ZN(new_n639));
  INV_X1    g0439(.A(new_n599), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n254), .B1(new_n615), .B2(KEYINPUT84), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n609), .A2(new_n610), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n639), .B(new_n640), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n621), .A2(new_n629), .A3(G190), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n644), .B1(new_n637), .B2(new_n517), .ZN(new_n645));
  OAI22_X1  g0445(.A1(new_n617), .A2(new_n638), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n558), .A2(new_n597), .A3(new_n646), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n476), .A2(new_n647), .ZN(G372));
  NAND2_X1  g0448(.A1(new_n425), .A2(new_n426), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n429), .ZN(new_n650));
  INV_X1    g0450(.A(new_n354), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n651), .A2(new_n473), .B1(new_n468), .B2(new_n452), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n650), .B1(new_n652), .B2(new_n408), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n319), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n323), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT88), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n619), .A2(new_n534), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n292), .B1(new_n658), .B2(new_n635), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n657), .B(new_n321), .C1(new_n659), .C2(new_n634), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n630), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n621), .A2(new_n629), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n657), .B1(new_n662), .B2(new_n321), .ZN(new_n663));
  OAI21_X1  g0463(.A(KEYINPUT89), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT88), .B1(new_n637), .B2(G169), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT89), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n665), .A2(new_n666), .A3(new_n630), .A4(new_n660), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n617), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n643), .A2(new_n645), .ZN(new_n669));
  NOR4_X1   g0469(.A1(new_n668), .A2(KEYINPUT26), .A3(new_n514), .A4(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT26), .B1(new_n646), .B2(new_n514), .ZN(new_n671));
  INV_X1    g0471(.A(new_n617), .ZN(new_n672));
  AOI21_X1  g0472(.A(G169), .B1(new_n621), .B2(new_n629), .ZN(new_n673));
  AOI22_X1  g0473(.A1(new_n657), .A2(new_n673), .B1(new_n637), .B2(new_n349), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n666), .B1(new_n674), .B2(new_n665), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n661), .A2(new_n663), .A3(KEYINPUT89), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n672), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n671), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n670), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n664), .A2(new_n667), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n669), .B1(new_n680), .B2(new_n672), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n516), .B1(new_n517), .B2(new_n512), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n491), .ZN(new_n683));
  AOI211_X1 g0483(.A(G179), .B(new_n508), .C1(new_n498), .C2(new_n293), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n515), .A2(new_n684), .A3(new_n510), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n681), .A2(KEYINPUT90), .A3(new_n686), .A4(new_n557), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n550), .A2(new_n594), .A3(new_n595), .A4(new_n596), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n557), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n668), .A2(new_n669), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(KEYINPUT90), .B1(new_n691), .B2(new_n686), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n679), .B1(new_n689), .B2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n656), .B1(new_n694), .B2(new_n475), .ZN(G369));
  NAND3_X1  g0495(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n210), .A2(new_n211), .A3(G13), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n697), .A2(KEYINPUT27), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(KEYINPUT27), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n698), .A2(G213), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(G343), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n575), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n696), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n705), .B1(new_n597), .B2(new_n704), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(G330), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n550), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n702), .B1(new_n544), .B2(new_n549), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n711), .B1(new_n557), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n550), .A2(new_n702), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n710), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n696), .A2(new_n703), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(new_n714), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n717), .A2(new_n720), .ZN(G399));
  INV_X1    g0521(.A(new_n214), .ZN(new_n722));
  INV_X1    g0522(.A(new_n285), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n606), .A2(G116), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(G1), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n219), .B2(new_n725), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT28), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT29), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n693), .A2(new_n730), .A3(new_n703), .ZN(new_n731));
  INV_X1    g0531(.A(new_n669), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n677), .A2(KEYINPUT26), .A3(new_n732), .A4(new_n685), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT26), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(new_n646), .B2(new_n514), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT94), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OAI211_X1 g0537(.A(KEYINPUT94), .B(new_n734), .C1(new_n646), .C2(new_n514), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n733), .A2(new_n737), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT95), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n683), .B2(new_n685), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n514), .A2(new_n518), .A3(KEYINPUT95), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n741), .A2(new_n688), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n677), .A2(new_n732), .A3(new_n557), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n677), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n703), .B1(new_n739), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(KEYINPUT29), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n731), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT31), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT93), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n662), .A2(new_n349), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n750), .B1(new_n589), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n499), .A2(new_n509), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n591), .A2(KEYINPUT93), .A3(new_n349), .A4(new_n662), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n752), .A2(new_n753), .A3(new_n754), .A4(new_n525), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n522), .A2(new_n293), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n523), .A2(G264), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(KEYINPUT91), .B1(new_n758), .B2(new_n662), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT91), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n637), .A2(new_n760), .A3(new_n524), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  OAI211_X1 g0562(.A(new_n580), .B(G179), .C1(new_n582), .C2(new_n583), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n753), .ZN(new_n764));
  AOI21_X1  g0564(.A(KEYINPUT92), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT30), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n755), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI211_X1 g0567(.A(KEYINPUT92), .B(KEYINPUT30), .C1(new_n762), .C2(new_n764), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n702), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n749), .A2(new_n769), .B1(new_n647), .B2(new_n703), .ZN(new_n770));
  OAI211_X1 g0570(.A(KEYINPUT31), .B(new_n702), .C1(new_n767), .C2(new_n768), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n708), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n748), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n729), .B1(new_n773), .B2(G1), .ZN(G364));
  AND2_X1   g0574(.A1(new_n211), .A2(G13), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n210), .B1(new_n775), .B2(G45), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n724), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G13), .A2(G33), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT97), .Z(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n707), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n211), .A2(G190), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n787), .A2(KEYINPUT98), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n517), .A2(G179), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n787), .A2(KEYINPUT98), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G179), .A2(G200), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n788), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G283), .A2(new_n792), .B1(new_n795), .B2(G329), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n349), .A2(new_n517), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n211), .A2(new_n401), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n349), .A2(G200), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G326), .A2(new_n800), .B1(new_n803), .B2(G322), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n798), .A2(new_n789), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n786), .A2(new_n801), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G303), .A2(new_n806), .B1(new_n808), .B2(G311), .ZN(new_n809));
  XOR2_X1   g0609(.A(KEYINPUT33), .B(G317), .Z(new_n810));
  NAND2_X1  g0610(.A1(new_n797), .A2(new_n786), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n392), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n211), .B1(new_n793), .B2(G190), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n812), .B1(G294), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n796), .A2(new_n804), .A3(new_n809), .A4(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT99), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n795), .A2(G159), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT32), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n791), .A2(new_n327), .ZN(new_n820));
  INV_X1    g0620(.A(new_n811), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G68), .A2(new_n821), .B1(new_n808), .B2(G77), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n822), .B1(new_n245), .B2(new_n799), .C1(new_n396), .C2(new_n805), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n298), .B1(new_n813), .B2(new_n478), .C1(new_n256), .C2(new_n802), .ZN(new_n824));
  NOR4_X1   g0624(.A1(new_n819), .A2(new_n820), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n817), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n221), .B1(G20), .B2(new_n321), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n784), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n722), .A2(new_n298), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(G45), .B2(new_n219), .ZN(new_n830));
  OR2_X1    g0630(.A1(new_n830), .A2(KEYINPUT96), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(KEYINPUT96), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n831), .B(new_n832), .C1(new_n286), .C2(new_n251), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n722), .A2(new_n392), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n834), .A2(G355), .B1(new_n567), .B2(new_n722), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n826), .A2(new_n827), .B1(new_n828), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n779), .B1(new_n785), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n706), .B(G330), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n838), .B1(new_n839), .B2(new_n779), .ZN(new_n840));
  XOR2_X1   g0640(.A(KEYINPUT100), .B(KEYINPUT101), .Z(new_n841));
  XNOR2_X1  g0641(.A(new_n840), .B(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G396));
  OAI21_X1  g0643(.A(new_n348), .B1(new_n344), .B2(new_n703), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n354), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n651), .A2(new_n703), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n693), .A2(new_n703), .A3(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n769), .A2(new_n749), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n558), .A2(new_n646), .ZN(new_n853));
  INV_X1    g0653(.A(new_n597), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n853), .A2(new_n854), .A3(new_n703), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n852), .A2(new_n771), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(G330), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n849), .B1(new_n693), .B2(new_n703), .ZN(new_n858));
  OR3_X1    g0658(.A1(new_n851), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n857), .B1(new_n851), .B2(new_n858), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n859), .A2(new_n779), .A3(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(G132), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n298), .B1(new_n794), .B2(new_n862), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT103), .Z(new_n864));
  AOI22_X1  g0664(.A1(G137), .A2(new_n800), .B1(new_n821), .B2(G150), .ZN(new_n865));
  AOI22_X1  g0665(.A1(G143), .A2(new_n803), .B1(new_n808), .B2(G159), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(KEYINPUT34), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n792), .A2(G68), .ZN(new_n869));
  AOI22_X1  g0669(.A1(new_n806), .A2(G50), .B1(new_n814), .B2(G58), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n867), .A2(KEYINPUT34), .ZN(new_n872));
  NOR3_X1   g0672(.A1(new_n864), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(G311), .ZN(new_n874));
  OAI22_X1  g0674(.A1(new_n396), .A2(new_n791), .B1(new_n794), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(G294), .ZN(new_n876));
  XNOR2_X1  g0676(.A(KEYINPUT102), .B(G283), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n876), .A2(new_n802), .B1(new_n811), .B2(new_n877), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n805), .A2(new_n327), .B1(new_n807), .B2(new_n567), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n392), .B1(new_n813), .B2(new_n478), .C1(new_n799), .C2(new_n578), .ZN(new_n880));
  NOR4_X1   g0680(.A1(new_n875), .A2(new_n878), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n827), .B1(new_n873), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n827), .A2(new_n780), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n779), .B1(new_n206), .B2(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n882), .B(new_n884), .C1(new_n849), .C2(new_n781), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n861), .A2(new_n885), .ZN(G384));
  OR2_X1    g0686(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n887), .A2(G116), .A3(new_n222), .A4(new_n888), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n889), .B(KEYINPUT36), .Z(new_n890));
  NAND3_X1  g0690(.A1(new_n220), .A2(G77), .A3(new_n359), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n210), .B(G13), .C1(new_n891), .C2(new_n246), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n655), .B1(new_n748), .B2(new_n476), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT106), .ZN(new_n895));
  INV_X1    g0695(.A(new_n700), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n431), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT37), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n404), .A2(new_n897), .A3(new_n898), .A4(new_n425), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n403), .A2(new_n389), .A3(new_n419), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n417), .B(new_n361), .C1(KEYINPUT105), .C2(KEYINPUT16), .ZN(new_n901));
  NOR2_X1   g0701(.A1(KEYINPUT105), .A2(KEYINPUT16), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n377), .B2(new_n380), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n901), .A2(new_n254), .A3(new_n903), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n904), .A2(new_n389), .B1(new_n411), .B2(new_n700), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT37), .B1(new_n900), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n899), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n904), .A2(new_n389), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n896), .ZN(new_n910));
  OAI211_X1 g0710(.A(new_n908), .B(KEYINPUT38), .C1(new_n435), .C2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT38), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n421), .B1(new_n420), .B2(KEYINPUT18), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n425), .A2(KEYINPUT81), .A3(new_n426), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n913), .A2(new_n914), .A3(new_n430), .A4(new_n433), .ZN(new_n915));
  INV_X1    g0715(.A(new_n407), .ZN(new_n916));
  AOI21_X1  g0716(.A(KEYINPUT17), .B1(new_n391), .B2(new_n403), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n910), .B1(new_n915), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n912), .B1(new_n919), .B2(new_n907), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n911), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n466), .A2(new_n467), .A3(new_n702), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n469), .A2(new_n473), .A3(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT104), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n452), .A2(new_n468), .A3(new_n702), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n925), .B1(new_n924), .B2(new_n926), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n929), .B1(new_n850), .B2(new_n847), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n922), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT39), .ZN(new_n932));
  NOR3_X1   g0732(.A1(new_n919), .A2(new_n912), .A3(new_n907), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n649), .A2(new_n429), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n431), .B(new_n896), .C1(new_n408), .C2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n404), .A2(new_n897), .A3(new_n425), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(KEYINPUT37), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n937), .A2(new_n899), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT38), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n932), .B1(new_n933), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n911), .A2(new_n920), .A3(KEYINPUT39), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n469), .A2(new_n702), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n934), .A2(new_n700), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n931), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n895), .B(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT40), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n927), .A2(new_n928), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(new_n856), .A3(new_n849), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n947), .B1(new_n921), .B2(new_n949), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n948), .A2(new_n849), .ZN(new_n951));
  INV_X1    g0751(.A(new_n938), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n897), .B1(new_n918), .B2(new_n650), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n912), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n911), .A2(new_n954), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n951), .A2(new_n955), .A3(KEYINPUT40), .A4(new_n856), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n950), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n476), .A2(new_n856), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n959), .A2(G330), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n946), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n210), .B2(new_n775), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n946), .A2(new_n961), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n893), .B1(new_n963), .B2(new_n964), .ZN(G367));
  OAI21_X1  g0765(.A(new_n828), .B1(new_n214), .B2(new_n338), .ZN(new_n966));
  INV_X1    g0766(.A(new_n829), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n967), .A2(new_n240), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n778), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  AOI22_X1  g0769(.A1(G77), .A2(new_n792), .B1(new_n795), .B2(G137), .ZN(new_n970));
  AOI22_X1  g0770(.A1(G143), .A2(new_n800), .B1(new_n806), .B2(G58), .ZN(new_n971));
  AOI22_X1  g0771(.A1(G159), .A2(new_n821), .B1(new_n808), .B2(G50), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n813), .A2(new_n247), .ZN(new_n973));
  AOI211_X1 g0773(.A(new_n392), .B(new_n973), .C1(G150), .C2(new_n803), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n970), .A2(new_n971), .A3(new_n972), .A4(new_n974), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT109), .Z(new_n976));
  INV_X1    g0776(.A(new_n877), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n800), .A2(G311), .B1(new_n808), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(KEYINPUT108), .B(G317), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n978), .B1(new_n578), .B2(new_n802), .C1(new_n794), .C2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n805), .A2(new_n567), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n392), .B1(new_n876), .B2(new_n811), .C1(new_n981), .C2(KEYINPUT46), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(KEYINPUT46), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n327), .B2(new_n813), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n791), .A2(new_n478), .ZN(new_n985));
  NOR4_X1   g0785(.A1(new_n980), .A2(new_n982), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n976), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT47), .ZN(new_n988));
  INV_X1    g0788(.A(new_n827), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n643), .A2(new_n702), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n677), .A2(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n681), .B2(new_n991), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n969), .B(new_n990), .C1(new_n784), .C2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n741), .A2(new_n742), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(new_n491), .B2(new_n702), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n514), .A2(new_n703), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n719), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT42), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  AND2_X1   g0801(.A1(new_n996), .A2(new_n711), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n703), .B1(new_n1002), .B2(new_n685), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1004), .A2(KEYINPUT107), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT107), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1001), .A2(new_n1006), .A3(new_n1003), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT43), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n993), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n716), .A2(new_n998), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n993), .B(new_n1009), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1005), .A2(new_n1007), .A3(new_n1013), .ZN(new_n1014));
  AND3_X1   g0814(.A1(new_n1011), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1012), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n773), .ZN(new_n1018));
  OR2_X1    g0818(.A1(new_n720), .A2(new_n998), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT44), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n720), .A2(new_n998), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT45), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n716), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1022), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT44), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1019), .B(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1024), .A2(new_n1026), .A3(new_n717), .ZN(new_n1027));
  AND2_X1   g0827(.A1(new_n1023), .A2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n715), .B(new_n718), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(new_n709), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1018), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n724), .B(KEYINPUT41), .Z(new_n1032));
  OAI21_X1  g0832(.A(new_n776), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n994), .B1(new_n1017), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(G387));
  AOI21_X1  g0835(.A(new_n725), .B1(new_n773), .B2(new_n1030), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n773), .B2(new_n1030), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n805), .A2(new_n206), .B1(new_n807), .B2(new_n247), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1038), .B(new_n985), .C1(G159), .C2(new_n800), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n298), .B1(new_n813), .B2(new_n338), .C1(new_n245), .C2(new_n802), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(new_n260), .B2(new_n821), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1039), .B(new_n1041), .C1(new_n266), .C2(new_n794), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n298), .B1(new_n795), .B2(G326), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G294), .A2(new_n806), .B1(new_n814), .B2(new_n977), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT110), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n811), .A2(new_n874), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n802), .A2(new_n979), .B1(new_n807), .B2(new_n578), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(G322), .C2(new_n800), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1046), .B1(new_n1049), .B2(KEYINPUT48), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(KEYINPUT48), .C2(new_n1049), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT49), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1043), .B1(new_n567), .B2(new_n791), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1042), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n827), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n726), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n834), .A2(new_n1058), .B1(new_n327), .B2(new_n722), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n237), .A2(new_n286), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n339), .A2(G50), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT50), .Z(new_n1062));
  OAI211_X1 g0862(.A(new_n726), .B(new_n286), .C1(new_n247), .C2(new_n206), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n829), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1059), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n779), .B1(new_n1065), .B2(new_n828), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1057), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n715), .B2(new_n784), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n1030), .B2(new_n777), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1037), .A2(new_n1069), .ZN(G393));
  NAND3_X1  g0870(.A1(new_n1023), .A2(new_n1027), .A3(new_n777), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n828), .B1(new_n478), .B2(new_n214), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n967), .A2(new_n244), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n778), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G87), .A2(new_n792), .B1(new_n795), .B2(G143), .ZN(new_n1075));
  INV_X1    g0875(.A(G159), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n799), .A2(new_n266), .B1(new_n802), .B2(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT51), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n813), .A2(new_n206), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n811), .A2(new_n245), .B1(new_n807), .B2(new_n339), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n392), .B(new_n1081), .C1(G68), .C2(new_n806), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1075), .A2(new_n1078), .A3(new_n1080), .A4(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n392), .B1(new_n807), .B2(new_n876), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1084), .B(new_n820), .C1(new_n806), .C2(new_n977), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G317), .A2(new_n800), .B1(new_n803), .B2(G311), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT52), .Z(new_n1087));
  NAND2_X1  g0887(.A1(new_n795), .A2(G322), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n811), .A2(new_n578), .B1(new_n813), .B2(new_n567), .ZN(new_n1090));
  XOR2_X1   g0890(.A(new_n1090), .B(KEYINPUT111), .Z(new_n1091));
  OAI21_X1  g0891(.A(new_n1083), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1074), .B1(new_n1092), .B2(new_n827), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n998), .B2(new_n783), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1071), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT112), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1071), .A2(KEYINPUT112), .A3(new_n1094), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1023), .A2(new_n1027), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n773), .A2(new_n1030), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1102), .A2(new_n724), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1099), .A2(new_n1104), .ZN(G390));
  NAND2_X1  g0905(.A1(new_n748), .A2(new_n476), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n857), .A2(new_n475), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1106), .A2(new_n656), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT114), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n894), .A2(KEYINPUT114), .A3(new_n1108), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT115), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n850), .A2(new_n847), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n948), .B1(new_n772), .B2(new_n849), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n856), .A2(G330), .A3(new_n849), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1117), .A2(new_n929), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1114), .B(new_n1115), .C1(new_n1116), .C2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n847), .B1(new_n746), .B2(new_n846), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n772), .A2(new_n849), .A3(new_n948), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1117), .A2(new_n929), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1119), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1114), .B1(new_n1126), .B2(new_n1115), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1125), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n940), .A2(new_n941), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n930), .B2(new_n942), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1122), .A2(KEYINPUT113), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n942), .B1(new_n911), .B2(new_n954), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n1121), .B2(new_n929), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1130), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1132), .B1(new_n1130), .B2(new_n1134), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1113), .A2(new_n1128), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(KEYINPUT114), .B1(new_n894), .B2(new_n1108), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n475), .B1(new_n731), .B2(new_n747), .ZN(new_n1140));
  NOR4_X1   g0940(.A1(new_n1140), .A2(new_n1110), .A3(new_n655), .A4(new_n1107), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1130), .A2(new_n1134), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n1131), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1115), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(KEYINPUT115), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1146), .A2(new_n1119), .A3(new_n1124), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1142), .A2(new_n1135), .A3(new_n1144), .A4(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1138), .A2(new_n1148), .A3(new_n724), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1144), .A2(new_n777), .A3(new_n1135), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n883), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n778), .B1(new_n260), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n869), .B1(new_n876), .B2(new_n794), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(G107), .A2(new_n821), .B1(new_n803), .B2(G116), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n800), .A2(G283), .B1(new_n808), .B2(G97), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n298), .B1(new_n806), .B2(G87), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1154), .A2(new_n1155), .A3(new_n1080), .A4(new_n1156), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1153), .A2(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(G132), .A2(new_n803), .B1(new_n821), .B2(G137), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT54), .B(G143), .ZN(new_n1160));
  INV_X1    g0960(.A(G125), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1159), .B1(new_n807), .B2(new_n1160), .C1(new_n794), .C2(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n805), .A2(new_n266), .ZN(new_n1163));
  XOR2_X1   g0963(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(G128), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1166), .B(new_n298), .C1(new_n1167), .C2(new_n799), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n1163), .A2(new_n1165), .B1(new_n1076), .B2(new_n813), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n791), .A2(new_n245), .ZN(new_n1170));
  NOR4_X1   g0970(.A1(new_n1162), .A2(new_n1168), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1158), .B1(new_n1172), .B2(KEYINPUT117), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(KEYINPUT117), .B2(new_n1172), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1152), .B1(new_n1174), .B2(new_n827), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1129), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1175), .B1(new_n1176), .B2(new_n781), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(KEYINPUT118), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT118), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1179), .B(new_n1175), .C1(new_n1176), .C2(new_n781), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n1150), .A2(KEYINPUT119), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT119), .B1(new_n1150), .B2(new_n1181), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1149), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT120), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1149), .B(KEYINPUT120), .C1(new_n1182), .C2(new_n1183), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(G378));
  INV_X1    g0988(.A(KEYINPUT57), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT122), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1144), .A2(new_n1135), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1190), .B(new_n1142), .C1(new_n1191), .C2(new_n1128), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n950), .A2(G330), .A3(new_n956), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n319), .A2(new_n323), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n320), .A2(new_n700), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  OR3_X1    g0999(.A1(new_n1196), .A2(new_n1197), .A3(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1199), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1193), .A2(new_n1203), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n950), .A2(new_n956), .A3(G330), .A4(new_n1202), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n945), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n945), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1208), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1192), .A2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1190), .B1(new_n1148), .B2(new_n1142), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1189), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1142), .B1(new_n1191), .B2(new_n1128), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(KEYINPUT122), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1215), .A2(KEYINPUT57), .A3(new_n1192), .A4(new_n1210), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1213), .A2(new_n724), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n776), .B1(new_n1207), .B2(new_n1209), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT121), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n779), .B1(new_n245), .B2(new_n883), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n799), .A2(new_n1161), .B1(new_n811), .B2(new_n862), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n808), .A2(G137), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1222), .B1(new_n1167), .B2(new_n802), .C1(new_n805), .C2(new_n1160), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1221), .B(new_n1223), .C1(G150), .C2(new_n814), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  OR2_X1    g1025(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(KEYINPUT59), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n792), .A2(G159), .ZN(new_n1228));
  AOI211_X1 g1028(.A(G33), .B(G41), .C1(new_n795), .C2(G124), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(G116), .A2(new_n800), .B1(new_n803), .B2(G107), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n791), .A2(new_n256), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G283), .B2(new_n795), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n298), .B(new_n723), .C1(new_n821), .C2(G97), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n807), .A2(new_n338), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n973), .B(new_n1235), .C1(G77), .C2(new_n806), .ZN(new_n1236));
  AND4_X1   g1036(.A1(new_n1231), .A2(new_n1233), .A3(new_n1234), .A4(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT58), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1237), .A2(KEYINPUT58), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n245), .B1(G33), .B2(G41), .C1(new_n723), .C2(new_n298), .ZN(new_n1240));
  AND4_X1   g1040(.A1(new_n1230), .A2(new_n1238), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1220), .B1(new_n989), .B2(new_n1241), .C1(new_n1202), .C2(new_n781), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  OR3_X1    g1043(.A1(new_n1218), .A2(new_n1219), .A3(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1219), .B1(new_n1218), .B2(new_n1243), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1217), .A2(new_n1246), .ZN(G375));
  AOI21_X1  g1047(.A(new_n779), .B1(new_n247), .B2(new_n883), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n799), .A2(new_n862), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT124), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1232), .B(new_n1250), .C1(G128), .C2(new_n795), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n1076), .A2(new_n805), .B1(new_n811), .B2(new_n1160), .ZN(new_n1252));
  OAI221_X1 g1052(.A(new_n298), .B1(new_n813), .B2(new_n245), .C1(new_n266), .C2(new_n807), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1252), .B(new_n1253), .C1(G137), .C2(new_n803), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n392), .B1(new_n813), .B2(new_n338), .C1(new_n567), .C2(new_n811), .ZN(new_n1255));
  INV_X1    g1055(.A(G283), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n802), .A2(new_n1256), .B1(new_n807), .B2(new_n327), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n799), .A2(new_n876), .B1(new_n805), .B2(new_n478), .ZN(new_n1258));
  NOR3_X1   g1058(.A1(new_n1255), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(G77), .A2(new_n792), .B1(new_n795), .B2(G303), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n1251), .A2(new_n1254), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1261));
  OAI221_X1 g1061(.A(new_n1248), .B1(new_n989), .B2(new_n1261), .C1(new_n948), .C2(new_n781), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n776), .B(KEYINPUT123), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1263), .B1(new_n1147), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1032), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(new_n1113), .B2(new_n1128), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1142), .A2(new_n1147), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1266), .B1(new_n1268), .B2(new_n1269), .ZN(G381));
  NAND3_X1  g1070(.A1(new_n1149), .A2(new_n1181), .A3(new_n1150), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(G375), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(G390), .ZN(new_n1274));
  INV_X1    g1074(.A(G384), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(G393), .A2(G396), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1034), .A2(new_n1274), .A3(new_n1275), .A4(new_n1276), .ZN(new_n1277));
  OR3_X1    g1077(.A1(new_n1273), .A2(G381), .A3(new_n1277), .ZN(G407));
  OAI211_X1 g1078(.A(G407), .B(G213), .C1(G343), .C2(new_n1273), .ZN(G409));
  NAND3_X1  g1079(.A1(G378), .A2(new_n1217), .A3(new_n1246), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1215), .A2(new_n1267), .A3(new_n1192), .A4(new_n1210), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1243), .B1(new_n1210), .B2(new_n1265), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1271), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1280), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(G213), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1286), .A2(G343), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT60), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1289), .B1(new_n1142), .B2(new_n1147), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1290), .A2(new_n1269), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1113), .A2(new_n1128), .A3(KEYINPUT60), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1292), .A2(new_n724), .ZN(new_n1293));
  OAI21_X1  g1093(.A(new_n1266), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT125), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1275), .A2(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1294), .A2(new_n1295), .A3(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(KEYINPUT60), .B1(new_n1113), .B2(new_n1128), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1113), .A2(new_n1128), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1301), .A2(new_n724), .A3(new_n1292), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1302), .A2(new_n1296), .A3(new_n1275), .A4(new_n1266), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1298), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1285), .A2(new_n1288), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(KEYINPUT62), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT61), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1287), .A2(G2897), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1304), .A2(new_n1308), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1298), .A2(new_n1303), .A3(G2897), .A4(new_n1287), .ZN(new_n1310));
  AND2_X1   g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1215), .A2(new_n1192), .A3(new_n1210), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n725), .B1(new_n1312), .B2(new_n1189), .ZN(new_n1313));
  AOI22_X1  g1113(.A1(new_n1313), .A2(new_n1216), .B1(new_n1245), .B2(new_n1244), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1283), .B1(new_n1314), .B2(G378), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1311), .B1(new_n1315), .B2(new_n1287), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1287), .B1(new_n1280), .B2(new_n1284), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT62), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1317), .A2(new_n1318), .A3(new_n1304), .ZN(new_n1319));
  NAND4_X1  g1119(.A1(new_n1306), .A2(new_n1307), .A3(new_n1316), .A4(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n842), .B1(new_n1037), .B2(new_n1069), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1276), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(G390), .A2(new_n1322), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n1099), .B(new_n1104), .C1(new_n1276), .C2(new_n1321), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1323), .A2(new_n1034), .A3(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1034), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1320), .A2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1330));
  OAI211_X1 g1130(.A(new_n1327), .B(new_n1307), .C1(new_n1317), .C2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1331), .ZN(new_n1332));
  AND2_X1   g1132(.A1(new_n1298), .A2(new_n1303), .ZN(new_n1333));
  AOI211_X1 g1133(.A(new_n1287), .B(new_n1333), .C1(new_n1280), .C2(new_n1284), .ZN(new_n1334));
  OAI21_X1  g1134(.A(KEYINPUT126), .B1(new_n1334), .B2(KEYINPUT63), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1334), .A2(KEYINPUT63), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT126), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT63), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1305), .A2(new_n1337), .A3(new_n1338), .ZN(new_n1339));
  NAND4_X1  g1139(.A1(new_n1332), .A2(new_n1335), .A3(new_n1336), .A4(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1329), .A2(new_n1340), .ZN(G405));
  INV_X1    g1141(.A(new_n1271), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(G375), .A2(new_n1342), .ZN(new_n1343));
  AND3_X1   g1143(.A1(new_n1343), .A2(new_n1280), .A3(new_n1304), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1304), .B1(new_n1343), .B2(new_n1280), .ZN(new_n1345));
  OR4_X1    g1145(.A1(KEYINPUT127), .A2(new_n1344), .A3(new_n1345), .A4(new_n1327), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT127), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1328), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1327), .A2(KEYINPUT127), .ZN(new_n1349));
  OAI211_X1 g1149(.A(new_n1348), .B(new_n1349), .C1(new_n1344), .C2(new_n1345), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1346), .A2(new_n1350), .ZN(G402));
endmodule


