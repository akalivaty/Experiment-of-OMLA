//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 1 1 0 1 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 0 1 0 1 1 1 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n814, new_n815, new_n816, new_n817, new_n819, new_n820, new_n821,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n948, new_n949, new_n950;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT24), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n203), .A2(G183gat), .A3(G190gat), .ZN(new_n204));
  INV_X1    g003(.A(G183gat), .ZN(new_n205));
  INV_X1    g004(.A(G190gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n204), .B1(new_n207), .B2(new_n203), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n205), .A2(new_n206), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G169gat), .ZN(new_n211));
  INV_X1    g010(.A(G176gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n213), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n214), .A2(KEYINPUT23), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n202), .B1(new_n210), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n214), .B(KEYINPUT65), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT23), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(G190gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(new_n205), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(new_n208), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n222), .A2(new_n225), .A3(KEYINPUT25), .A4(new_n217), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n220), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT27), .B(G183gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT28), .ZN(new_n230));
  XNOR2_X1  g029(.A(new_n229), .B(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT26), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n221), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n213), .B1(KEYINPUT26), .B2(new_n215), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n207), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(new_n235), .A3(KEYINPUT67), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT67), .B1(new_n231), .B2(new_n235), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n227), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(G113gat), .B(G120gat), .Z(new_n240));
  INV_X1    g039(.A(KEYINPUT1), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G127gat), .B(G134gat), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n240), .A2(new_n241), .A3(new_n243), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n239), .A2(new_n247), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n220), .A2(new_n226), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n235), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n249), .B1(new_n252), .B2(new_n236), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n245), .A2(new_n246), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n248), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G227gat), .A2(G233gat), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT32), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT33), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(G15gat), .B(G43gat), .Z(new_n263));
  XNOR2_X1  g062(.A(G71gat), .B(G99gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n260), .A2(new_n262), .A3(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n255), .A3(new_n257), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n267), .A2(KEYINPUT34), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(KEYINPUT34), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n268), .B1(KEYINPUT68), .B2(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n257), .B1(new_n248), .B2(new_n255), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n265), .B1(new_n271), .B2(KEYINPUT33), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT32), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n267), .A2(new_n276), .A3(KEYINPUT34), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n266), .A2(new_n270), .A3(new_n275), .A4(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n269), .A2(KEYINPUT68), .ZN(new_n279));
  OR2_X1    g078(.A1(new_n267), .A2(KEYINPUT34), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n279), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n272), .A2(new_n274), .ZN(new_n282));
  AOI221_X4 g081(.A(new_n273), .B1(KEYINPUT33), .B2(new_n265), .C1(new_n256), .C2(new_n258), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n278), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT69), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT36), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n278), .A2(KEYINPUT69), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT85), .ZN(new_n291));
  XNOR2_X1  g090(.A(G141gat), .B(G148gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT79), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT2), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(new_n293), .B2(new_n292), .ZN(new_n295));
  NAND2_X1  g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT78), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n296), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n299), .B1(new_n298), .B2(new_n297), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n295), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT80), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT81), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT2), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n297), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n302), .A2(new_n292), .B1(new_n305), .B2(new_n296), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n296), .A2(KEYINPUT2), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(new_n303), .ZN(new_n308));
  OAI211_X1 g107(.A(new_n306), .B(new_n308), .C1(new_n302), .C2(new_n292), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n301), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT3), .ZN(new_n311));
  XOR2_X1   g110(.A(KEYINPUT83), .B(KEYINPUT3), .Z(new_n312));
  NAND3_X1  g111(.A1(new_n301), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n254), .A2(KEYINPUT82), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT82), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n247), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g115(.A1(new_n311), .A2(new_n313), .A3(new_n314), .A4(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G225gat), .A2(G233gat), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT5), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n254), .A2(new_n309), .A3(new_n301), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT84), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n254), .A2(new_n301), .A3(KEYINPUT84), .A4(new_n309), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(KEYINPUT4), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT4), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n321), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n319), .A2(new_n320), .A3(new_n326), .A4(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n314), .A2(new_n310), .A3(new_n316), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n323), .A2(new_n330), .A3(new_n324), .ZN(new_n331));
  INV_X1    g130(.A(new_n318), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n320), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n323), .A2(new_n327), .A3(new_n324), .ZN(new_n334));
  INV_X1    g133(.A(new_n310), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(KEYINPUT4), .A3(new_n254), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n334), .A2(new_n317), .A3(new_n318), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n329), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G1gat), .B(G29gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(KEYINPUT0), .ZN(new_n341));
  XNOR2_X1  g140(.A(G57gat), .B(G85gat), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n341), .B(new_n342), .Z(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n291), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n339), .A2(new_n344), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT6), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n329), .A2(new_n338), .A3(KEYINPUT85), .A4(new_n343), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n345), .A2(new_n346), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n339), .A2(KEYINPUT6), .A3(new_n344), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n226), .A2(new_n220), .B1(new_n231), .B2(new_n235), .ZN(new_n352));
  NAND2_X1  g151(.A1(G226gat), .A2(G233gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT72), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n354), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT29), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n355), .B1(new_n253), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G211gat), .B(G218gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT70), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n362));
  INV_X1    g161(.A(G197gat), .ZN(new_n363));
  INV_X1    g162(.A(G204gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G197gat), .A2(G204gat), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n362), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OR2_X1    g166(.A1(new_n367), .A2(KEYINPUT71), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n361), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT70), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n360), .B(new_n370), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n367), .A2(KEYINPUT71), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT73), .B1(new_n359), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n239), .A2(new_n357), .A3(new_n356), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT73), .ZN(new_n377));
  INV_X1    g176(.A(new_n374), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n376), .A2(new_n377), .A3(new_n378), .A4(new_n355), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n356), .B1(new_n352), .B2(KEYINPUT29), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n381), .B(new_n374), .C1(new_n253), .C2(new_n356), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT74), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n239), .A2(new_n354), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n385), .A2(KEYINPUT74), .A3(new_n374), .A4(new_n381), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G8gat), .B(G36gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(G64gat), .B(G92gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n380), .A2(new_n387), .A3(KEYINPUT30), .A4(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT77), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI22_X1  g195(.A1(new_n375), .A2(new_n379), .B1(new_n384), .B2(new_n386), .ZN(new_n397));
  NAND4_X1  g196(.A1(new_n397), .A2(KEYINPUT77), .A3(KEYINPUT30), .A4(new_n393), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n393), .B1(new_n380), .B2(new_n387), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n397), .A2(new_n393), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT30), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n351), .A2(new_n399), .A3(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT31), .B(G50gat), .ZN(new_n405));
  INV_X1    g204(.A(G106gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G228gat), .A2(G233gat), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n369), .A2(new_n373), .A3(new_n357), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n310), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT87), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n409), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n412), .A2(KEYINPUT87), .A3(new_n310), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n374), .B1(new_n357), .B2(new_n313), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n417), .A2(KEYINPUT88), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT88), .ZN(new_n419));
  AOI211_X1 g218(.A(new_n419), .B(new_n374), .C1(new_n357), .C2(new_n313), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n415), .B(new_n416), .C1(new_n418), .C2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G22gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n361), .A2(KEYINPUT86), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT86), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n371), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(new_n425), .A3(new_n367), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n426), .B(new_n357), .C1(new_n367), .C2(new_n425), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n335), .B1(new_n427), .B2(new_n312), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n409), .B1(new_n428), .B2(new_n417), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n421), .A2(new_n422), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n422), .B1(new_n421), .B2(new_n429), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n431), .A2(G78gat), .A3(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(G78gat), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n421), .A2(new_n429), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(G22gat), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n434), .B1(new_n436), .B2(new_n430), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n408), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(G78gat), .B1(new_n431), .B2(new_n432), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n436), .A2(new_n434), .A3(new_n430), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(new_n440), .A3(new_n407), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n404), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n285), .A2(KEYINPUT36), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n290), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n349), .A2(new_n350), .A3(new_n401), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT37), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n380), .A2(new_n387), .A3(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n385), .A2(new_n378), .A3(new_n381), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n449), .B(KEYINPUT37), .C1(new_n378), .C2(new_n359), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n392), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT38), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n380), .A2(new_n387), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT37), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n455), .A2(KEYINPUT38), .A3(new_n392), .A4(new_n448), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n446), .A2(new_n457), .ZN(new_n458));
  AND2_X1   g257(.A1(new_n438), .A2(new_n441), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n399), .A2(new_n403), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n326), .A2(new_n317), .A3(new_n328), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n332), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n331), .A2(new_n332), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT39), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n344), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  XOR2_X1   g265(.A(KEYINPUT89), .B(KEYINPUT39), .Z(new_n467));
  NAND3_X1  g266(.A1(new_n461), .A2(new_n332), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(KEYINPUT40), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n346), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT40), .B1(new_n466), .B2(new_n468), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n460), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n458), .A2(new_n459), .A3(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n438), .A2(new_n278), .A3(new_n284), .A4(new_n441), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT35), .B1(new_n475), .B2(new_n404), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT69), .B1(new_n278), .B2(new_n284), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n278), .A2(KEYINPUT69), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n351), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(new_n460), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT35), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n438), .A2(new_n482), .A3(new_n441), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n445), .A2(new_n474), .B1(new_n476), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(G43gat), .A2(G50gat), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(G43gat), .A2(G50gat), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT15), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OR3_X1    g288(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n488), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT15), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n493), .A2(new_n494), .A3(new_n486), .ZN(new_n495));
  INV_X1    g294(.A(G29gat), .ZN(new_n496));
  INV_X1    g295(.A(G36gat), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  AND4_X1   g298(.A1(new_n489), .A2(new_n492), .A3(new_n495), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n491), .A2(KEYINPUT90), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT90), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n502), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n501), .A2(new_n490), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n489), .B1(new_n504), .B2(new_n499), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT91), .B1(new_n500), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT91), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n492), .A2(new_n495), .A3(new_n489), .A4(new_n499), .ZN(new_n508));
  NOR3_X1   g307(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n509), .B1(KEYINPUT90), .B2(new_n491), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n498), .B1(new_n510), .B2(new_n503), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n507), .B(new_n508), .C1(new_n511), .C2(new_n489), .ZN(new_n512));
  XNOR2_X1  g311(.A(G15gat), .B(G22gat), .ZN(new_n513));
  INV_X1    g312(.A(G1gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT16), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n516), .B1(G1gat), .B2(new_n513), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(G8gat), .ZN(new_n518));
  INV_X1    g317(.A(G8gat), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n516), .B(new_n519), .C1(G1gat), .C2(new_n513), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n506), .A2(new_n512), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT93), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n506), .A2(new_n512), .A3(new_n521), .A4(KEYINPUT93), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n506), .A2(new_n512), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n526), .B1(new_n528), .B2(new_n521), .ZN(new_n529));
  NAND2_X1  g328(.A1(G229gat), .A2(G233gat), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n530), .B(KEYINPUT13), .Z(new_n531));
  NAND2_X1  g330(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT18), .ZN(new_n533));
  XOR2_X1   g332(.A(KEYINPUT92), .B(KEYINPUT17), .Z(new_n534));
  NAND3_X1  g333(.A1(new_n506), .A2(new_n512), .A3(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n500), .A2(new_n505), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n521), .B1(KEYINPUT17), .B2(new_n536), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n524), .A2(new_n525), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  AOI211_X1 g337(.A(KEYINPUT94), .B(new_n533), .C1(new_n538), .C2(new_n530), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n535), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n526), .A2(new_n530), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT94), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT18), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n532), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G113gat), .B(G141gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n545), .B(G197gat), .ZN(new_n546));
  XOR2_X1   g345(.A(KEYINPUT11), .B(G169gat), .Z(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n548), .B(KEYINPUT12), .Z(new_n549));
  NAND2_X1  g348(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n549), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n532), .B(new_n551), .C1(new_n539), .C2(new_n543), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G71gat), .A2(G78gat), .ZN(new_n555));
  INV_X1    g354(.A(G71gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(new_n434), .ZN(new_n557));
  XNOR2_X1  g356(.A(G57gat), .B(G64gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT9), .ZN(new_n559));
  OAI211_X1 g358(.A(new_n555), .B(new_n557), .C1(new_n558), .C2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT95), .ZN(new_n561));
  INV_X1    g360(.A(G57gat), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n561), .B1(new_n562), .B2(G64gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(G64gat), .ZN(new_n564));
  INV_X1    g363(.A(G64gat), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n565), .A2(KEYINPUT95), .A3(G57gat), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n555), .B1(new_n557), .B2(new_n559), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n560), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT21), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT96), .ZN(new_n573));
  XOR2_X1   g372(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(G183gat), .B(G211gat), .Z(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT98), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n575), .B(new_n577), .ZN(new_n578));
  AND2_X1   g377(.A1(new_n560), .A2(new_n569), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n521), .B1(KEYINPUT21), .B2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT97), .ZN(new_n581));
  XNOR2_X1  g380(.A(G127gat), .B(G155gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n581), .B(new_n584), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n578), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n578), .A2(new_n585), .ZN(new_n587));
  AND2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G230gat), .A2(G233gat), .ZN(new_n590));
  XOR2_X1   g389(.A(KEYINPUT103), .B(KEYINPUT10), .Z(new_n591));
  XNOR2_X1  g390(.A(G99gat), .B(G106gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G85gat), .A2(G92gat), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT7), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n594), .B1(new_n595), .B2(KEYINPUT100), .ZN(new_n596));
  NAND2_X1  g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(KEYINPUT8), .ZN(new_n598));
  OR2_X1    g397(.A1(G85gat), .A2(G92gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n595), .A2(KEYINPUT101), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n596), .A2(new_n598), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NOR4_X1   g400(.A1(new_n594), .A2(new_n595), .A3(KEYINPUT100), .A4(KEYINPUT101), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n593), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT8), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n604), .B1(G99gat), .B2(G106gat), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT101), .ZN(new_n606));
  OAI22_X1  g405(.A1(new_n606), .A2(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n595), .A2(KEYINPUT100), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n609), .A2(new_n606), .A3(G85gat), .A4(G92gat), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n608), .A2(new_n592), .A3(new_n610), .A4(new_n596), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n603), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(KEYINPUT102), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(new_n613), .A3(new_n579), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n611), .B(new_n603), .C1(new_n570), .C2(KEYINPUT102), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n591), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT10), .ZN(new_n617));
  NOR3_X1   g416(.A1(new_n612), .A2(new_n617), .A3(new_n570), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n590), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G120gat), .B(G148gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(G176gat), .B(G204gat), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n620), .B(new_n621), .Z(new_n622));
  NAND2_X1  g421(.A1(new_n614), .A2(new_n615), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n619), .B(new_n622), .C1(new_n590), .C2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n590), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n619), .A2(KEYINPUT104), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT104), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n627), .B(new_n590), .C1(new_n616), .C2(new_n618), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n625), .B1(new_n626), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n624), .B1(new_n629), .B2(new_n622), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT105), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT105), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n632), .B(new_n624), .C1(new_n629), .C2(new_n622), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n536), .A2(KEYINPUT17), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n535), .A2(new_n636), .A3(new_n612), .ZN(new_n637));
  AND2_X1   g436(.A1(G232gat), .A2(G233gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT41), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n637), .B(new_n639), .C1(new_n527), .C2(new_n612), .ZN(new_n640));
  XOR2_X1   g439(.A(G190gat), .B(G218gat), .Z(new_n641));
  OR2_X1    g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n638), .A2(KEYINPUT41), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT99), .ZN(new_n644));
  XNOR2_X1  g443(.A(G134gat), .B(G162gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n640), .A2(new_n641), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n642), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n646), .B1(new_n642), .B2(new_n647), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n589), .A2(new_n635), .A3(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n485), .A2(new_n554), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n480), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(G1gat), .ZN(G1324gat));
  INV_X1    g454(.A(KEYINPUT42), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n653), .A2(new_n460), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT106), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT16), .B(G8gat), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n656), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(G8gat), .ZN(new_n661));
  OR3_X1    g460(.A1(new_n657), .A2(new_n656), .A3(new_n659), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(G1325gat));
  INV_X1    g462(.A(G15gat), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n653), .A2(new_n664), .A3(new_n479), .ZN(new_n665));
  AND2_X1   g464(.A1(new_n290), .A2(new_n444), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n653), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n665), .B1(new_n668), .B2(new_n664), .ZN(G1326gat));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n442), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT43), .B(G22gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1327gat));
  NAND4_X1  g471(.A1(new_n474), .A2(new_n444), .A3(new_n290), .A4(new_n443), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n484), .A2(new_n476), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n651), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n589), .A2(new_n554), .A3(new_n634), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n675), .A2(new_n496), .A3(new_n480), .A4(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n677), .B(KEYINPUT107), .Z(new_n678));
  OR2_X1    g477(.A1(new_n678), .A2(KEYINPUT45), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n675), .A2(KEYINPUT108), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n675), .A2(KEYINPUT108), .A3(KEYINPUT44), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n676), .ZN(new_n685));
  OAI21_X1  g484(.A(G29gat), .B1(new_n685), .B2(new_n351), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n678), .A2(KEYINPUT45), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n679), .A2(new_n686), .A3(new_n687), .ZN(G1328gat));
  INV_X1    g487(.A(new_n460), .ZN(new_n689));
  OAI21_X1  g488(.A(G36gat), .B1(new_n685), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n676), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n691), .A2(G36gat), .A3(new_n689), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n690), .A2(new_n694), .ZN(G1329gat));
  INV_X1    g494(.A(new_n479), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n691), .A2(G43gat), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT110), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n682), .A2(new_n667), .A3(new_n683), .A4(new_n676), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(G43gat), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT47), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n698), .A2(KEYINPUT47), .A3(new_n700), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(G1330gat));
  INV_X1    g504(.A(KEYINPUT111), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n691), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n459), .A2(G50gat), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT48), .ZN(new_n709));
  AOI22_X1  g508(.A1(new_n707), .A2(new_n708), .B1(KEYINPUT112), .B2(new_n709), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n709), .A2(KEYINPUT112), .ZN(new_n711));
  NAND4_X1  g510(.A1(new_n682), .A2(new_n442), .A3(new_n683), .A4(new_n676), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(G50gat), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n711), .B1(new_n710), .B2(new_n713), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(G1331gat));
  NAND3_X1  g515(.A1(new_n589), .A2(new_n554), .A3(new_n651), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n485), .A2(new_n635), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n480), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n460), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n721), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT49), .B(G64gat), .Z(new_n723));
  OAI21_X1  g522(.A(new_n722), .B1(new_n721), .B2(new_n723), .ZN(G1333gat));
  AOI21_X1  g523(.A(new_n556), .B1(new_n718), .B2(new_n667), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n696), .A2(G71gat), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(new_n718), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g527(.A1(new_n718), .A2(new_n442), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g529(.A1(new_n589), .A2(new_n635), .A3(new_n553), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n684), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(G85gat), .B1(new_n732), .B2(new_n351), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n589), .A2(new_n553), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT113), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n675), .B2(new_n735), .ZN(new_n736));
  AOI211_X1 g535(.A(KEYINPUT113), .B(new_n651), .C1(new_n673), .C2(new_n674), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT51), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT113), .B1(new_n485), .B2(new_n651), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n675), .A2(new_n735), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT51), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n739), .A2(new_n740), .A3(new_n741), .A4(new_n734), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n351), .A2(new_n635), .A3(G85gat), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n733), .A2(new_n745), .ZN(G1336gat));
  NAND4_X1  g545(.A1(new_n682), .A2(new_n460), .A3(new_n683), .A4(new_n731), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G92gat), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n689), .A2(new_n635), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(G92gat), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n736), .B2(new_n737), .ZN(new_n754));
  INV_X1    g553(.A(new_n753), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n739), .A2(new_n740), .A3(new_n734), .A4(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n752), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT115), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n748), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AOI211_X1 g558(.A(KEYINPUT115), .B(new_n752), .C1(new_n754), .C2(new_n756), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT52), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n743), .A2(new_n751), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n762), .A2(new_n763), .A3(new_n748), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n764), .ZN(G1337gat));
  OAI21_X1  g564(.A(G99gat), .B1(new_n732), .B2(new_n666), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n696), .A2(G99gat), .A3(new_n635), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n743), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n768), .ZN(G1338gat));
  NAND4_X1  g568(.A1(new_n682), .A2(new_n442), .A3(new_n683), .A4(new_n731), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(G106gat), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(KEYINPUT53), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n459), .A2(G106gat), .A3(new_n635), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n738), .A2(new_n742), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT116), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n738), .A2(new_n742), .A3(new_n776), .A4(new_n773), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n772), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n773), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n780), .B1(new_n754), .B2(new_n756), .ZN(new_n781));
  OAI21_X1  g580(.A(KEYINPUT53), .B1(new_n771), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n782), .ZN(G1339gat));
  NOR2_X1   g582(.A1(new_n717), .A2(new_n634), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n529), .A2(new_n531), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n538), .A2(new_n530), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n548), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n552), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n634), .A2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n626), .A2(new_n628), .A3(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n622), .ZN(new_n793));
  OR3_X1    g592(.A1(new_n616), .A2(new_n590), .A3(new_n618), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(KEYINPUT54), .A3(new_n619), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n792), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n792), .A2(new_n795), .A3(KEYINPUT55), .A4(new_n793), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(new_n624), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n553), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n650), .B1(new_n790), .B2(new_n802), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n801), .A2(new_n789), .A3(new_n650), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n588), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n785), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n480), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n807), .A2(new_n460), .A3(new_n475), .ZN(new_n808));
  AOI21_X1  g607(.A(G113gat), .B1(new_n808), .B2(new_n553), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(new_n459), .A3(new_n479), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n810), .A2(new_n351), .A3(new_n460), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n553), .A2(G113gat), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n809), .B1(new_n811), .B2(new_n812), .ZN(G1340gat));
  INV_X1    g612(.A(G120gat), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n814), .B1(new_n811), .B2(new_n634), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT117), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n808), .A2(new_n814), .A3(new_n634), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1341gat));
  NAND2_X1  g617(.A1(new_n811), .A2(new_n589), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n588), .A2(G127gat), .ZN(new_n820));
  AOI22_X1  g619(.A1(new_n819), .A2(G127gat), .B1(new_n808), .B2(new_n820), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n821), .B(KEYINPUT118), .ZN(G1342gat));
  INV_X1    g621(.A(G134gat), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n823), .A3(new_n650), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n824), .A2(KEYINPUT56), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n823), .B1(new_n811), .B2(new_n650), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n827), .B1(KEYINPUT56), .B2(new_n824), .ZN(G1343gat));
  NOR2_X1   g627(.A1(new_n807), .A2(KEYINPUT122), .ZN(new_n829));
  NOR4_X1   g628(.A1(new_n829), .A2(new_n460), .A3(new_n459), .A4(new_n667), .ZN(new_n830));
  INV_X1    g629(.A(G141gat), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n807), .A2(KEYINPUT122), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n830), .A2(new_n831), .A3(new_n553), .A4(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n460), .A2(new_n351), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n666), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n442), .A2(KEYINPUT57), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT119), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n796), .A2(new_n797), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n799), .A2(new_n624), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n798), .A2(KEYINPUT119), .A3(new_n624), .A4(new_n799), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n553), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n790), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(KEYINPUT120), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT120), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n843), .A2(new_n846), .A3(new_n790), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n651), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n804), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n650), .B1(new_n844), .B2(KEYINPUT120), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(KEYINPUT121), .A3(new_n847), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n589), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n837), .B1(new_n853), .B2(new_n784), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n459), .B1(new_n785), .B2(new_n805), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(KEYINPUT57), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  AOI211_X1 g656(.A(new_n554), .B(new_n835), .C1(new_n854), .C2(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n833), .B1(new_n858), .B2(new_n831), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n860), .B1(new_n858), .B2(new_n831), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n859), .A2(new_n861), .A3(KEYINPUT58), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT58), .ZN(new_n863));
  OAI221_X1 g662(.A(new_n833), .B1(new_n860), .B2(new_n863), .C1(new_n858), .C2(new_n831), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(G1344gat));
  AND2_X1   g664(.A1(new_n830), .A2(new_n832), .ZN(new_n866));
  INV_X1    g665(.A(G148gat), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n867), .A3(new_n634), .ZN(new_n868));
  INV_X1    g667(.A(new_n835), .ZN(new_n869));
  AND4_X1   g668(.A1(new_n552), .A2(new_n631), .A3(new_n633), .A4(new_n788), .ZN(new_n870));
  AOI22_X1  g669(.A1(new_n800), .A2(new_n838), .B1(new_n550), .B2(new_n552), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n842), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n651), .B1(new_n872), .B2(new_n846), .ZN(new_n873));
  INV_X1    g672(.A(new_n847), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n849), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n804), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n875), .A2(new_n876), .A3(new_n852), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n588), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n836), .B1(new_n878), .B2(new_n785), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n634), .B(new_n869), .C1(new_n879), .C2(new_n856), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n867), .A2(KEYINPUT59), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n881), .B1(new_n880), .B2(new_n882), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n804), .B1(new_n851), .B2(new_n847), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n785), .B1(new_n887), .B2(new_n589), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT57), .B1(new_n888), .B2(new_n442), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n836), .B1(new_n785), .B2(new_n805), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n869), .B(new_n634), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT125), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n867), .B1(new_n891), .B2(new_n892), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n886), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n868), .B1(new_n885), .B2(new_n895), .ZN(G1345gat));
  INV_X1    g695(.A(G155gat), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n866), .A2(new_n897), .A3(new_n589), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n835), .B1(new_n854), .B2(new_n857), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n899), .A2(new_n589), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n898), .B1(new_n897), .B2(new_n900), .ZN(G1346gat));
  AOI21_X1  g700(.A(G162gat), .B1(new_n866), .B2(new_n650), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n650), .A2(G162gat), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n899), .B2(new_n903), .ZN(G1347gat));
  AOI21_X1  g703(.A(new_n480), .B1(new_n785), .B2(new_n805), .ZN(new_n905));
  INV_X1    g704(.A(new_n475), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n907), .A2(new_n689), .ZN(new_n908));
  AOI21_X1  g707(.A(G169gat), .B1(new_n908), .B2(new_n553), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n810), .A2(new_n480), .A3(new_n689), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n554), .A2(new_n211), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n909), .B1(new_n910), .B2(new_n911), .ZN(G1348gat));
  AOI21_X1  g711(.A(new_n212), .B1(new_n910), .B2(new_n634), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n907), .A2(G176gat), .A3(new_n750), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n913), .A2(new_n914), .ZN(G1349gat));
  AOI21_X1  g714(.A(new_n205), .B1(new_n910), .B2(new_n589), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT126), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(KEYINPUT60), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n908), .A2(new_n228), .A3(new_n589), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n917), .A2(KEYINPUT60), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n920), .B(new_n921), .ZN(G1350gat));
  AOI21_X1  g721(.A(new_n206), .B1(new_n910), .B2(new_n650), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n923), .B(KEYINPUT61), .Z(new_n924));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n223), .A3(new_n650), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1351gat));
  OR2_X1    g725(.A1(new_n889), .A2(new_n890), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n666), .A2(new_n351), .A3(new_n460), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n930), .A2(new_n363), .A3(new_n554), .ZN(new_n931));
  AND4_X1   g730(.A1(new_n460), .A2(new_n905), .A3(new_n442), .A4(new_n666), .ZN(new_n932));
  AOI21_X1  g731(.A(G197gat), .B1(new_n932), .B2(new_n553), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n931), .A2(new_n933), .ZN(G1352gat));
  NAND3_X1  g733(.A1(new_n932), .A2(new_n364), .A3(new_n634), .ZN(new_n935));
  XOR2_X1   g734(.A(new_n935), .B(KEYINPUT62), .Z(new_n936));
  AND3_X1   g735(.A1(new_n927), .A2(new_n634), .A3(new_n929), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n364), .B2(new_n937), .ZN(G1353gat));
  INV_X1    g737(.A(G211gat), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT63), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(KEYINPUT127), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n941), .B1(new_n930), .B2(new_n588), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(new_n943), .A3(KEYINPUT63), .ZN(new_n944));
  OAI221_X1 g743(.A(new_n941), .B1(KEYINPUT127), .B2(new_n940), .C1(new_n930), .C2(new_n588), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n932), .A2(new_n939), .A3(new_n589), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n944), .A2(new_n945), .A3(new_n946), .ZN(G1354gat));
  OAI21_X1  g746(.A(G218gat), .B1(new_n930), .B2(new_n651), .ZN(new_n948));
  INV_X1    g747(.A(G218gat), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n932), .A2(new_n949), .A3(new_n650), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1355gat));
endmodule


