//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 1 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n544, new_n546, new_n547, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n451), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n461), .A2(new_n462), .A3(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(KEYINPUT66), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n466));
  OAI211_X1 g041(.A(new_n460), .B(new_n463), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G137), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n462), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n464), .A2(G2105), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n469), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n483), .B1(new_n467), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n462), .A2(G2104), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n471), .B1(new_n486), .B2(KEYINPUT66), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n487), .A2(G2105), .A3(new_n463), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n485), .B1(G124), .B2(new_n489), .ZN(G162));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  OAI21_X1  g066(.A(KEYINPUT4), .B1(new_n467), .B2(new_n491), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n491), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n493), .A2(new_n471), .A3(new_n472), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G126), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n460), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  OAI22_X1  g073(.A1(new_n488), .A2(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n495), .A2(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  OAI21_X1  g076(.A(G543), .B1(new_n501), .B2(KEYINPUT67), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT5), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT6), .B(G651), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(G543), .ZN(new_n511));
  OAI22_X1  g086(.A1(new_n508), .A2(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  XOR2_X1   g088(.A(new_n513), .B(KEYINPUT69), .Z(new_n514));
  NAND2_X1  g089(.A1(new_n506), .A2(G62), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n514), .B1(new_n515), .B2(KEYINPUT68), .ZN(new_n516));
  OAI21_X1  g091(.A(new_n516), .B1(KEYINPUT68), .B2(new_n515), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n512), .B1(new_n517), .B2(G651), .ZN(G166));
  INV_X1    g093(.A(new_n511), .ZN(new_n519));
  XOR2_X1   g094(.A(KEYINPUT70), .B(G51), .Z(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n506), .A2(G89), .A3(new_n507), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n521), .A2(new_n522), .A3(new_n523), .A4(new_n525), .ZN(G286));
  INV_X1    g101(.A(G286), .ZN(G168));
  INV_X1    g102(.A(G90), .ZN(new_n528));
  INV_X1    g103(.A(G52), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n508), .A2(new_n528), .B1(new_n529), .B2(new_n511), .ZN(new_n530));
  INV_X1    g105(.A(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n506), .A2(G64), .ZN(new_n532));
  NAND2_X1  g107(.A1(G77), .A2(G543), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n530), .A2(new_n534), .ZN(G171));
  INV_X1    g110(.A(G81), .ZN(new_n536));
  INV_X1    g111(.A(G43), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n508), .A2(new_n536), .B1(new_n537), .B2(new_n511), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n506), .A2(G56), .ZN(new_n539));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n531), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  AND3_X1   g118(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G36), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n544), .A2(new_n547), .ZN(G188));
  INV_X1    g123(.A(KEYINPUT9), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(KEYINPUT71), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n549), .A2(KEYINPUT71), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n519), .A2(G53), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(G53), .ZN(new_n553));
  OAI211_X1 g128(.A(KEYINPUT71), .B(new_n549), .C1(new_n511), .C2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(KEYINPUT72), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n502), .A2(new_n505), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n531), .A2(KEYINPUT6), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT6), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G651), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT73), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT73), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n507), .A2(new_n563), .A3(new_n502), .A4(new_n505), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n557), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n565), .A2(G91), .B1(G651), .B2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT72), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n552), .A2(new_n554), .A3(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n556), .A2(new_n569), .A3(new_n571), .ZN(G299));
  INV_X1    g147(.A(G171), .ZN(G301));
  INV_X1    g148(.A(G166), .ZN(G303));
  NAND2_X1  g149(.A1(new_n565), .A2(G87), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT74), .ZN(new_n576));
  OAI211_X1 g151(.A(new_n576), .B(G651), .C1(new_n506), .C2(G74), .ZN(new_n577));
  AOI21_X1  g152(.A(G74), .B1(new_n502), .B2(new_n505), .ZN(new_n578));
  OAI21_X1  g153(.A(KEYINPUT74), .B1(new_n578), .B2(new_n531), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  AND3_X1   g155(.A1(new_n507), .A2(G49), .A3(G543), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n575), .A2(new_n580), .A3(new_n582), .ZN(G288));
  NAND2_X1  g158(.A1(new_n519), .A2(G48), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n585), .B2(new_n531), .ZN(new_n586));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n562), .B2(new_n564), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G305));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  XOR2_X1   g166(.A(KEYINPUT75), .B(G47), .Z(new_n592));
  OAI22_X1  g167(.A1(new_n508), .A2(new_n591), .B1(new_n511), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n506), .A2(G60), .ZN(new_n594));
  NAND2_X1  g169(.A1(G72), .A2(G543), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n531), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n557), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(new_n519), .B2(G54), .ZN(new_n603));
  AND3_X1   g178(.A1(new_n565), .A2(KEYINPUT10), .A3(G92), .ZN(new_n604));
  AOI21_X1  g179(.A(KEYINPUT10), .B1(new_n565), .B2(G92), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n599), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n599), .B1(new_n607), .B2(G868), .ZN(G321));
  NAND2_X1  g184(.A1(G286), .A2(G868), .ZN(new_n610));
  INV_X1    g185(.A(G299), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G297));
  OAI21_X1  g187(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND2_X1  g190(.A1(new_n607), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n542), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n468), .A2(G135), .ZN(new_n620));
  INV_X1    g195(.A(G123), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n460), .A2(G111), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  OAI221_X1 g198(.A(new_n620), .B1(new_n621), .B2(new_n488), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(G2096), .Z(new_n625));
  NAND3_X1  g200(.A1(new_n460), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT12), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT76), .B(KEYINPUT13), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n625), .A2(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  INV_X1    g210(.A(KEYINPUT79), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n634), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n639), .A2(G2438), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(G2438), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2430), .ZN(new_n643));
  OR2_X1    g218(.A1(new_n643), .A2(KEYINPUT78), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n643), .A2(KEYINPUT78), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g222(.A1(new_n640), .A2(new_n644), .A3(new_n641), .A4(new_n645), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(new_n648), .A3(KEYINPUT14), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n638), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n652), .A2(KEYINPUT80), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(KEYINPUT80), .ZN(new_n654));
  INV_X1    g229(.A(G14), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n650), .B2(new_n651), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n653), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(G401));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(G2084), .B(G2090), .Z(new_n662));
  OR3_X1    g237(.A1(new_n661), .A2(KEYINPUT81), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(KEYINPUT81), .B1(new_n661), .B2(new_n662), .ZN(new_n664));
  INV_X1    g239(.A(new_n659), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n660), .B(KEYINPUT17), .Z(new_n666));
  OAI211_X1 g241(.A(new_n663), .B(new_n664), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(new_n662), .A3(new_n665), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n662), .A2(new_n659), .A3(new_n660), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT18), .Z(new_n670));
  NAND3_X1  g245(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2096), .B(G2100), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  OR2_X1    g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n674), .A2(new_n675), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n676), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT82), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n678), .A2(new_n680), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n681), .A2(new_n683), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n684), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT83), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(G229));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G6), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n589), .B2(new_n700), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT32), .B(G1981), .Z(new_n703));
  XOR2_X1   g278(.A(new_n702), .B(new_n703), .Z(new_n704));
  NAND2_X1  g279(.A1(new_n700), .A2(G22), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G166), .B2(new_n700), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n704), .B1(G1971), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(G16), .A2(G23), .ZN(new_n708));
  NAND2_X1  g283(.A1(G288), .A2(KEYINPUT89), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n581), .B1(new_n565), .B2(G87), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT89), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n710), .A2(new_n711), .A3(new_n580), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n708), .B1(new_n713), .B2(G16), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT33), .B(G1976), .Z(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n706), .A2(G1971), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n707), .A2(new_n716), .A3(new_n717), .A4(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT34), .Z(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT84), .B(G29), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n722), .A2(G25), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n468), .A2(G131), .ZN(new_n724));
  INV_X1    g299(.A(G119), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n460), .A2(G107), .ZN(new_n726));
  OAI21_X1  g301(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n727));
  OAI221_X1 g302(.A(new_n724), .B1(new_n725), .B2(new_n488), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n723), .B1(new_n728), .B2(new_n721), .ZN(new_n729));
  MUX2_X1   g304(.A(new_n723), .B(new_n729), .S(KEYINPUT85), .Z(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT35), .B(G1991), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT86), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT87), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n730), .B(new_n733), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n700), .A2(G24), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT88), .Z(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n597), .B2(new_n700), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(G1986), .Z(new_n738));
  NAND3_X1  g313(.A1(new_n720), .A2(new_n734), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n607), .A2(G16), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G4), .B2(G16), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G2090), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n722), .A2(G35), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G162), .B2(new_n722), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT29), .Z(new_n748));
  AOI22_X1  g323(.A1(new_n744), .A2(G1348), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(new_n745), .B2(new_n748), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n722), .A2(G27), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G164), .B2(new_n722), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n752), .A2(G2078), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n700), .A2(G5), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G171), .B2(new_n700), .ZN(new_n755));
  INV_X1    g330(.A(G1961), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n700), .A2(G19), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(new_n542), .B2(new_n700), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT91), .B(G1341), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G139), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n467), .A2(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT93), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(G115), .A2(G2104), .ZN(new_n766));
  INV_X1    g341(.A(G127), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n473), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n477), .A2(G103), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT25), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n477), .A2(KEYINPUT25), .A3(G103), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n768), .A2(G2105), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n765), .A2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(G29), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n775), .B2(G33), .ZN(new_n777));
  INV_X1    g352(.A(G2072), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n757), .B(new_n761), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  AOI211_X1 g354(.A(new_n753), .B(new_n779), .C1(new_n778), .C2(new_n777), .ZN(new_n780));
  NOR2_X1   g355(.A1(G168), .A2(new_n700), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n700), .B2(G21), .ZN(new_n782));
  INV_X1    g357(.A(G1966), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G2084), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT24), .B(G34), .Z(new_n786));
  OAI22_X1  g361(.A1(new_n480), .A2(new_n775), .B1(new_n721), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n784), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(G28), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n789), .A2(KEYINPUT30), .ZN(new_n790));
  AOI21_X1  g365(.A(G29), .B1(new_n789), .B2(KEYINPUT30), .ZN(new_n791));
  OR2_X1    g366(.A1(KEYINPUT31), .A2(G11), .ZN(new_n792));
  NAND2_X1  g367(.A1(KEYINPUT31), .A2(G11), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n790), .A2(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI221_X1 g369(.A(new_n794), .B1(new_n624), .B2(new_n722), .C1(new_n782), .C2(new_n783), .ZN(new_n795));
  NOR2_X1   g370(.A1(G29), .A2(G32), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n489), .A2(G129), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n468), .A2(G141), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n477), .A2(G105), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT94), .B(KEYINPUT26), .ZN(new_n800));
  NAND3_X1  g375(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(new_n801), .B2(new_n800), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n797), .A2(new_n798), .A3(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n796), .B1(new_n805), .B2(G29), .ZN(new_n806));
  XOR2_X1   g381(.A(KEYINPUT27), .B(G1996), .Z(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT95), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n806), .B(new_n808), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n788), .A2(new_n795), .A3(new_n809), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n780), .B(new_n810), .C1(G1348), .C2(new_n744), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT23), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n700), .A2(G20), .ZN(new_n813));
  AOI211_X1 g388(.A(new_n812), .B(new_n813), .C1(G299), .C2(G16), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n812), .B2(new_n813), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT97), .B(G1956), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n787), .A2(new_n785), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT96), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n722), .A2(G26), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT92), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT28), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n468), .A2(G140), .ZN(new_n823));
  INV_X1    g398(.A(G128), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n460), .A2(G116), .ZN(new_n825));
  OAI21_X1  g400(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n826));
  OAI221_X1 g401(.A(new_n823), .B1(new_n824), .B2(new_n488), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(G29), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n822), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G2067), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(G2078), .B2(new_n752), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n817), .A2(new_n819), .A3(new_n831), .ZN(new_n832));
  NOR4_X1   g407(.A1(new_n741), .A2(new_n750), .A3(new_n811), .A4(new_n832), .ZN(G311));
  OR4_X1    g408(.A1(new_n741), .A2(new_n750), .A3(new_n811), .A4(new_n832), .ZN(G150));
  INV_X1    g409(.A(G93), .ZN(new_n835));
  INV_X1    g410(.A(G55), .ZN(new_n836));
  OAI22_X1  g411(.A1(new_n508), .A2(new_n835), .B1(new_n836), .B2(new_n511), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n506), .A2(G67), .ZN(new_n838));
  NAND2_X1  g413(.A1(G80), .A2(G543), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n531), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(G860), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT37), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n607), .A2(G559), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT38), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n841), .A2(new_n542), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n538), .A2(new_n541), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n837), .A2(new_n840), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n845), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT39), .ZN(new_n852));
  AOI21_X1  g427(.A(G860), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n851), .A2(new_n852), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n853), .B1(new_n854), .B2(KEYINPUT98), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n854), .A2(KEYINPUT98), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n843), .B1(new_n855), .B2(new_n856), .ZN(G145));
  XNOR2_X1  g432(.A(new_n624), .B(new_n480), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(G162), .Z(new_n859));
  INV_X1    g434(.A(G142), .ZN(new_n860));
  OAI21_X1  g435(.A(KEYINPUT101), .B1(new_n460), .B2(G118), .ZN(new_n861));
  OR2_X1    g436(.A1(G106), .A2(G2105), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n861), .A2(G2104), .A3(new_n862), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n460), .A2(KEYINPUT101), .A3(G118), .ZN(new_n864));
  OAI22_X1  g439(.A1(new_n467), .A2(new_n860), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(G130), .B2(new_n489), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n728), .B(new_n866), .Z(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT102), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n627), .ZN(new_n869));
  INV_X1    g444(.A(new_n499), .ZN(new_n870));
  AND3_X1   g445(.A1(new_n492), .A2(KEYINPUT99), .A3(new_n494), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT99), .B1(new_n492), .B2(new_n494), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n774), .A2(KEYINPUT100), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n827), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n804), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n875), .A2(new_n804), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n873), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n878), .ZN(new_n880));
  INV_X1    g455(.A(new_n873), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n880), .A2(new_n881), .A3(new_n876), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n869), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n869), .B1(new_n879), .B2(new_n882), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n859), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  INV_X1    g461(.A(new_n627), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n868), .B(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n881), .B1(new_n880), .B2(new_n876), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n877), .A2(new_n873), .A3(new_n878), .ZN(new_n890));
  OAI211_X1 g465(.A(KEYINPUT103), .B(new_n888), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n869), .A2(new_n879), .A3(new_n882), .ZN(new_n892));
  INV_X1    g467(.A(new_n859), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n884), .A2(KEYINPUT103), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n885), .B(new_n886), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g472(.A1(G303), .A2(new_n589), .ZN(new_n898));
  NAND2_X1  g473(.A1(G166), .A2(G305), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n898), .A2(new_n597), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n597), .B1(new_n898), .B2(new_n899), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n901), .A2(KEYINPUT106), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT106), .ZN(new_n904));
  XNOR2_X1  g479(.A(G166), .B(G305), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(G290), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n904), .B1(new_n906), .B2(new_n900), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n713), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT106), .B1(new_n901), .B2(new_n902), .ZN(new_n909));
  INV_X1    g484(.A(new_n713), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(new_n904), .A3(new_n900), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT42), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n850), .B(KEYINPUT104), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(new_n616), .ZN(new_n916));
  XNOR2_X1  g491(.A(G299), .B(new_n606), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(KEYINPUT41), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT105), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n611), .A2(new_n606), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n921), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n919), .B1(new_n923), .B2(KEYINPUT41), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n918), .B1(new_n916), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n914), .B(new_n925), .ZN(new_n926));
  MUX2_X1   g501(.A(new_n841), .B(new_n926), .S(G868), .Z(G295));
  MUX2_X1   g502(.A(new_n841), .B(new_n926), .S(G868), .Z(G331));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n929));
  NAND2_X1  g504(.A1(G301), .A2(G168), .ZN(new_n930));
  NAND2_X1  g505(.A1(G171), .A2(G286), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g507(.A(new_n932), .B(new_n850), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n929), .B1(new_n933), .B2(new_n917), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n932), .A2(new_n850), .ZN(new_n935));
  AOI22_X1  g510(.A1(new_n930), .A2(new_n931), .B1(new_n846), .B2(new_n849), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n917), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(KEYINPUT107), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n924), .B2(new_n933), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n886), .B1(new_n941), .B2(new_n913), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n943));
  AOI22_X1  g518(.A1(new_n942), .A2(new_n943), .B1(new_n913), .B2(new_n941), .ZN(new_n944));
  OAI211_X1 g519(.A(KEYINPUT108), .B(new_n886), .C1(new_n941), .C2(new_n913), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT43), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(G37), .B1(new_n941), .B2(new_n913), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n903), .A2(new_n907), .A3(new_n713), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n910), .B1(new_n909), .B2(new_n911), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT41), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n937), .B1(new_n951), .B2(new_n917), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n921), .B(KEYINPUT41), .C1(new_n920), .C2(new_n922), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(new_n953), .A3(KEYINPUT109), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT110), .B1(new_n933), .B2(new_n917), .ZN(new_n955));
  OR3_X1    g530(.A1(new_n933), .A2(KEYINPUT110), .A3(new_n917), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT109), .B1(new_n952), .B2(new_n953), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n950), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n947), .A2(new_n959), .A3(KEYINPUT43), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT44), .B1(new_n946), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n947), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n942), .A2(new_n943), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n941), .A2(new_n913), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n945), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n963), .B1(new_n966), .B2(KEYINPUT43), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n961), .B1(KEYINPUT44), .B2(new_n967), .ZN(G397));
  XOR2_X1   g543(.A(new_n827), .B(G2067), .Z(new_n969));
  INV_X1    g544(.A(G1996), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n804), .B(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g547(.A(new_n728), .B(new_n732), .Z(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(G290), .A2(G1986), .ZN(new_n975));
  AND2_X1   g550(.A1(G290), .A2(G1986), .ZN(new_n976));
  OR3_X1    g551(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(KEYINPUT111), .B(G1384), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n873), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  XOR2_X1   g556(.A(KEYINPUT112), .B(G40), .Z(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n469), .A2(new_n476), .A3(new_n479), .A4(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n977), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  XOR2_X1   g562(.A(KEYINPUT113), .B(G8), .Z(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n492), .A2(new_n494), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT99), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n492), .A2(KEYINPUT99), .A3(new_n494), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(G1384), .B1(new_n994), .B2(new_n870), .ZN(new_n995));
  INV_X1    g570(.A(new_n984), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n989), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OR3_X1    g572(.A1(new_n586), .A2(G1981), .A3(new_n588), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n508), .A2(new_n587), .ZN(new_n999));
  OAI21_X1  g574(.A(G1981), .B1(new_n586), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT49), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n998), .A2(KEYINPUT49), .A3(new_n1000), .ZN(new_n1004));
  AND2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI211_X1 g580(.A(G1976), .B(G288), .C1(new_n1005), .C2(new_n997), .ZN(new_n1006));
  XOR2_X1   g581(.A(new_n998), .B(KEYINPUT115), .Z(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n997), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  AND4_X1   g584(.A1(new_n711), .A2(new_n575), .A3(new_n580), .A4(new_n582), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n711), .B1(new_n710), .B2(new_n580), .ZN(new_n1011));
  OAI21_X1  g586(.A(G1976), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G1384), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n873), .A2(new_n1013), .A3(new_n996), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1012), .A2(KEYINPUT114), .A3(new_n1014), .A4(new_n988), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n1016));
  INV_X1    g591(.A(G288), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(G1976), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1014), .A2(new_n1018), .A3(new_n988), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1015), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT114), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(new_n713), .B2(G1976), .ZN(new_n1022));
  OAI211_X1 g597(.A(new_n1022), .B(new_n997), .C1(KEYINPUT52), .C2(new_n1018), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1020), .A2(new_n1023), .B1(new_n1005), .B2(new_n997), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n873), .A2(new_n1025), .A3(new_n1013), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1013), .B1(new_n495), .B2(new_n499), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n984), .B1(new_n1027), .B2(KEYINPUT50), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(G2090), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n873), .A2(KEYINPUT45), .A3(new_n978), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n984), .B1(new_n1027), .B2(new_n980), .ZN(new_n1032));
  AOI21_X1  g607(.A(G1971), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1030), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(G8), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(G166), .B2(new_n1035), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1024), .A2(new_n1036), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1009), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1025), .B1(new_n873), .B2(new_n1013), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n996), .B1(new_n1027), .B2(KEYINPUT50), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT116), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1384), .B1(new_n870), .B2(new_n990), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n984), .B1(new_n1047), .B2(new_n1025), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT116), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1048), .B(new_n1049), .C1(new_n995), .C2(new_n1025), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1046), .A2(new_n1050), .A3(new_n745), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1033), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1040), .B1(new_n1053), .B2(new_n988), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1055));
  OAI211_X1 g630(.A(G8), .B(new_n1040), .C1(new_n1030), .C2(new_n1033), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1005), .A2(new_n997), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1054), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT45), .B1(new_n873), .B2(new_n1013), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n996), .B1(new_n1027), .B2(new_n980), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n783), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1026), .A2(new_n1028), .A3(new_n785), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n988), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1065), .A2(G286), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT63), .B1(new_n1059), .B2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g642(.A(new_n1066), .B(KEYINPUT63), .C1(new_n1036), .C2(new_n1040), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1068), .A2(new_n1058), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1043), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT61), .ZN(new_n1071));
  INV_X1    g646(.A(G1956), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT56), .B(G2072), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1031), .A2(new_n1032), .A3(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n555), .A2(KEYINPUT57), .ZN(new_n1077));
  AOI22_X1  g652(.A1(G299), .A2(KEYINPUT57), .B1(new_n569), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1076), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT121), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1078), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT121), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1073), .A2(new_n1078), .A3(new_n1075), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n1087));
  XNOR2_X1  g662(.A(new_n1086), .B(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1071), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1031), .A2(new_n1032), .A3(new_n970), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  XOR2_X1   g667(.A(KEYINPUT58), .B(G1341), .Z(new_n1093));
  AOI22_X1  g668(.A1(new_n1090), .A2(new_n1091), .B1(new_n1014), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n847), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  XOR2_X1   g672(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(G1348), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1014), .A2(G2067), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n606), .B1(new_n1102), .B2(KEYINPUT60), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT60), .ZN(new_n1104));
  NOR4_X1   g679(.A1(new_n1100), .A2(new_n1101), .A3(new_n1104), .A4(new_n607), .ZN(new_n1105));
  OAI22_X1  g680(.A1(new_n1103), .A2(new_n1105), .B1(KEYINPUT60), .B2(new_n1102), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1083), .A2(KEYINPUT118), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT118), .ZN(new_n1108));
  AOI211_X1 g683(.A(new_n1108), .B(new_n1078), .C1(new_n1073), .C2(new_n1075), .ZN(new_n1109));
  OAI211_X1 g684(.A(KEYINPUT61), .B(new_n1086), .C1(new_n1107), .C2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1089), .A2(new_n1099), .A3(new_n1106), .A4(new_n1110), .ZN(new_n1111));
  OAI22_X1  g686(.A1(new_n1107), .A2(new_n1109), .B1(new_n606), .B2(new_n1102), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1086), .B(KEYINPUT117), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1111), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n1116));
  INV_X1    g691(.A(G2078), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1031), .A2(new_n1032), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1118), .A2(new_n1119), .B1(new_n1029), .B2(new_n756), .ZN(new_n1120));
  AND4_X1   g695(.A1(KEYINPUT53), .A2(G160), .A3(G40), .A4(new_n1117), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n981), .A2(new_n1031), .A3(new_n1121), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1120), .A2(G301), .A3(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1124), .A2(KEYINPUT53), .A3(new_n1117), .ZN(new_n1125));
  AOI21_X1  g700(.A(G301), .B1(new_n1120), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1116), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g704(.A(KEYINPUT122), .B(new_n1116), .C1(new_n1123), .C2(new_n1126), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1116), .B1(new_n1132), .B2(G171), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1120), .A2(new_n1125), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1133), .B1(G171), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(G168), .A2(new_n989), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1064), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT51), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1064), .A2(G8), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1136), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AOI211_X1 g716(.A(KEYINPUT51), .B(new_n1136), .C1(new_n1064), .C2(new_n988), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1137), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1135), .A2(new_n1059), .A3(new_n1143), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1131), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1070), .B1(new_n1115), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1148), .B(new_n1137), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1149), .A2(new_n1059), .A3(new_n1126), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1065), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1035), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1152));
  OAI21_X1  g727(.A(KEYINPUT51), .B1(new_n1152), .B2(new_n1136), .ZN(new_n1153));
  AOI22_X1  g728(.A1(new_n1151), .A2(new_n1153), .B1(new_n1136), .B2(new_n1064), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1154), .A2(new_n1148), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1147), .B1(new_n1150), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1143), .A2(KEYINPUT62), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n989), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1024), .B(new_n1056), .C1(new_n1158), .C2(new_n1040), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1126), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1157), .A2(new_n1161), .A3(KEYINPUT123), .A4(new_n1149), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n1156), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n987), .B1(new_n1146), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT46), .ZN(new_n1165));
  INV_X1    g740(.A(new_n985), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1165), .B1(new_n1166), .B2(G1996), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n985), .A2(KEYINPUT46), .A3(new_n970), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n969), .A2(new_n805), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1167), .B(new_n1168), .C1(new_n1166), .C2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g745(.A(new_n1170), .B(KEYINPUT47), .ZN(new_n1171));
  AOI21_X1  g746(.A(KEYINPUT48), .B1(new_n985), .B2(new_n975), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1172), .B1(new_n974), .B2(new_n985), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n985), .A2(KEYINPUT48), .A3(new_n975), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n728), .A2(new_n732), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n972), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1176), .B1(G2067), .B2(new_n827), .ZN(new_n1177));
  AOI22_X1  g752(.A1(new_n1173), .A2(new_n1174), .B1(new_n1177), .B2(new_n985), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1171), .A2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT124), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(KEYINPUT125), .B1(new_n1164), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1059), .A2(new_n1066), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT63), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1069), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1042), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1083), .B(new_n1081), .ZN(new_n1188));
  AOI21_X1  g763(.A(KEYINPUT61), .B1(new_n1188), .B2(new_n1113), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1110), .A2(new_n1106), .ZN(new_n1190));
  NOR2_X1   g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AOI22_X1  g766(.A1(new_n1191), .A2(new_n1099), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1154), .A2(new_n1159), .ZN(new_n1193));
  NAND4_X1  g768(.A1(new_n1193), .A2(new_n1135), .A3(new_n1129), .A4(new_n1130), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1187), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1156), .A2(new_n1162), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n986), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT125), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1197), .A2(new_n1198), .A3(new_n1180), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1182), .A2(new_n1199), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g775(.A1(G227), .A2(new_n458), .ZN(new_n1202));
  AND2_X1   g776(.A1(new_n657), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g777(.A1(new_n698), .A2(KEYINPUT126), .A3(new_n1203), .ZN(new_n1204));
  NOR2_X1   g778(.A1(new_n695), .A2(new_n697), .ZN(new_n1205));
  OR2_X1    g779(.A1(new_n692), .A2(new_n694), .ZN(new_n1206));
  NAND2_X1  g780(.A1(new_n692), .A2(new_n694), .ZN(new_n1207));
  AOI21_X1  g781(.A(new_n696), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g782(.A(new_n1203), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1209));
  INV_X1    g783(.A(KEYINPUT126), .ZN(new_n1210));
  NAND2_X1  g784(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  AND2_X1   g785(.A1(new_n1204), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g786(.A1(new_n896), .A2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g787(.A(KEYINPUT127), .B1(new_n967), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g788(.A1(new_n1204), .A2(new_n1211), .ZN(new_n1215));
  OAI21_X1  g789(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n1216));
  NAND2_X1  g790(.A1(new_n1216), .A2(new_n892), .ZN(new_n1217));
  AOI21_X1  g791(.A(G37), .B1(new_n1217), .B2(new_n859), .ZN(new_n1218));
  INV_X1    g792(.A(KEYINPUT103), .ZN(new_n1219));
  NAND2_X1  g793(.A1(new_n1216), .A2(new_n1219), .ZN(new_n1220));
  NAND4_X1  g794(.A1(new_n1220), .A2(new_n891), .A3(new_n892), .A4(new_n893), .ZN(new_n1221));
  AOI21_X1  g795(.A(new_n1215), .B1(new_n1218), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n1223));
  AOI21_X1  g797(.A(new_n962), .B1(new_n944), .B2(new_n945), .ZN(new_n1224));
  OAI211_X1 g798(.A(new_n1222), .B(new_n1223), .C1(new_n1224), .C2(new_n963), .ZN(new_n1225));
  AND2_X1   g799(.A1(new_n1214), .A2(new_n1225), .ZN(G308));
  NAND2_X1  g800(.A1(new_n1214), .A2(new_n1225), .ZN(G225));
endmodule


