//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n764, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT24), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  OR2_X1    g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212));
  INV_X1    g011(.A(G169gat), .ZN(new_n213));
  INV_X1    g012(.A(G176gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT64), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n220), .A2(G169gat), .A3(G176gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n211), .A2(new_n217), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT25), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n223), .A2(KEYINPUT65), .A3(new_n224), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n208), .A2(KEYINPUT66), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n206), .A2(new_n230), .A3(new_n207), .ZN(new_n231));
  NAND4_X1  g030(.A1(new_n229), .A2(new_n209), .A3(new_n210), .A4(new_n231), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n232), .A2(KEYINPUT25), .A3(new_n222), .A4(new_n217), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n227), .A2(new_n228), .A3(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT28), .ZN(new_n235));
  INV_X1    g034(.A(G190gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(KEYINPUT67), .A2(G183gat), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n236), .B1(new_n237), .B2(KEYINPUT27), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT27), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n239), .B1(KEYINPUT67), .B2(G183gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n235), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT68), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n243), .B(new_n235), .C1(new_n238), .C2(new_n240), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT27), .B(G183gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n245), .A2(KEYINPUT28), .A3(new_n236), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n242), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n248));
  OR3_X1    g047(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n222), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n247), .A2(new_n250), .A3(new_n206), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT29), .ZN(new_n253));
  NAND2_X1  g052(.A1(G226gat), .A2(G233gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G197gat), .B(G204gat), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT22), .ZN(new_n257));
  INV_X1    g056(.A(G211gat), .ZN(new_n258));
  INV_X1    g057(.A(G218gat), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(G211gat), .B(G218gat), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n262), .A2(new_n256), .A3(new_n260), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n254), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n234), .A2(new_n251), .A3(new_n267), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n255), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n266), .B1(new_n255), .B2(new_n268), .ZN(new_n270));
  OAI211_X1 g069(.A(KEYINPUT30), .B(new_n205), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n266), .ZN(new_n272));
  AOI211_X1 g071(.A(KEYINPUT29), .B(new_n267), .C1(new_n234), .C2(new_n251), .ZN(new_n273));
  INV_X1    g072(.A(new_n268), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n255), .A2(new_n266), .A3(new_n268), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n276), .A3(new_n204), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n280));
  XNOR2_X1  g079(.A(G1gat), .B(G29gat), .ZN(new_n281));
  INV_X1    g080(.A(G85gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT0), .B(G57gat), .ZN(new_n284));
  XOR2_X1   g083(.A(new_n283), .B(new_n284), .Z(new_n285));
  NAND2_X1  g084(.A1(G225gat), .A2(G233gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(G127gat), .B(G134gat), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT1), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT69), .ZN(new_n289));
  INV_X1    g088(.A(G113gat), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n289), .A2(new_n290), .A3(G120gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n287), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G120gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G113gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n290), .A2(G120gat), .ZN(new_n295));
  AND3_X1   g094(.A1(new_n294), .A2(new_n295), .A3(KEYINPUT69), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT70), .B1(new_n292), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G127gat), .ZN(new_n298));
  INV_X1    g097(.A(G134gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G127gat), .A2(G134gat), .ZN(new_n301));
  AOI21_X1  g100(.A(KEYINPUT1), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n294), .A2(new_n295), .A3(KEYINPUT69), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n302), .A2(new_n303), .A3(new_n304), .A4(new_n291), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n297), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n294), .A2(new_n295), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n287), .B1(new_n288), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311));
  OR2_X1    g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n311), .B1(new_n312), .B2(KEYINPUT2), .ZN(new_n313));
  INV_X1    g112(.A(G148gat), .ZN(new_n314));
  INV_X1    g113(.A(G141gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT73), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G141gat), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n314), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n314), .A2(KEYINPUT74), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G148gat), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n315), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n313), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT3), .ZN(new_n325));
  NOR2_X1   g124(.A1(G141gat), .A2(G148gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT2), .ZN(new_n328));
  NAND2_X1  g127(.A1(G141gat), .A2(G148gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n330), .A2(new_n311), .A3(new_n312), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n324), .A2(new_n325), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n324), .A2(new_n331), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT3), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n310), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n308), .B1(new_n297), .B2(new_n305), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT4), .ZN(new_n337));
  XNOR2_X1  g136(.A(KEYINPUT74), .B(G148gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(KEYINPUT73), .B(G141gat), .ZN(new_n339));
  OAI22_X1  g138(.A1(new_n315), .A2(new_n338), .B1(new_n339), .B2(new_n314), .ZN(new_n340));
  INV_X1    g139(.A(new_n311), .ZN(new_n341));
  AND2_X1   g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n342), .A2(new_n326), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n341), .B1(new_n343), .B2(new_n328), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n340), .A2(new_n313), .B1(new_n344), .B2(new_n312), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n336), .A2(new_n337), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n337), .B1(new_n336), .B2(new_n345), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n286), .B(new_n335), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT5), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n310), .A2(new_n333), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n306), .A2(new_n345), .A3(new_n309), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n286), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(KEYINPUT4), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n337), .A3(new_n345), .ZN(new_n355));
  AOI22_X1  g154(.A1(new_n306), .A2(new_n309), .B1(new_n333), .B2(KEYINPUT3), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n354), .A2(new_n355), .B1(new_n356), .B2(new_n332), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n353), .B1(new_n357), .B2(new_n286), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n285), .B(new_n350), .C1(new_n358), .C2(new_n349), .ZN(new_n359));
  INV_X1    g158(.A(new_n285), .ZN(new_n360));
  INV_X1    g159(.A(new_n286), .ZN(new_n361));
  INV_X1    g160(.A(new_n352), .ZN(new_n362));
  NOR2_X1   g161(.A1(new_n336), .A2(new_n345), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n349), .B1(new_n348), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT5), .B1(new_n357), .B2(new_n286), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n360), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT6), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n359), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n365), .A2(new_n366), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n370), .A2(KEYINPUT6), .A3(new_n285), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n279), .A2(new_n280), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT75), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n275), .A2(new_n276), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT30), .B1(new_n374), .B2(new_n205), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n278), .A2(KEYINPUT72), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n372), .A2(new_n373), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n369), .A2(new_n371), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n271), .A2(new_n280), .A3(new_n277), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n379), .A2(new_n380), .A3(new_n376), .A4(new_n377), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(KEYINPUT75), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n332), .A2(new_n253), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT77), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n332), .A2(KEYINPUT77), .A3(new_n253), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n386), .A2(new_n272), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT78), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n386), .A2(KEYINPUT78), .A3(new_n272), .A4(new_n387), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT29), .B1(new_n264), .B2(new_n265), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n333), .B1(new_n392), .B2(KEYINPUT3), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n390), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(G228gat), .A2(G233gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT76), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n392), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT3), .B1(new_n392), .B2(new_n397), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n345), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n266), .B1(new_n332), .B2(new_n253), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n400), .A2(new_n401), .A3(new_n395), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n396), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT31), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT31), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n396), .A2(new_n406), .A3(new_n403), .ZN(new_n407));
  XOR2_X1   g206(.A(G22gat), .B(G50gat), .Z(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n405), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n406), .B1(new_n396), .B2(new_n403), .ZN(new_n411));
  AOI211_X1 g210(.A(KEYINPUT31), .B(new_n402), .C1(new_n394), .C2(new_n395), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(G78gat), .B(G106gat), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n410), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n414), .B1(new_n410), .B2(new_n413), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n383), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n234), .A2(new_n251), .A3(new_n336), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT71), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n252), .A2(new_n310), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n234), .A2(new_n251), .A3(KEYINPUT71), .A4(new_n336), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(G227gat), .A2(G233gat), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT33), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G15gat), .B(G43gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(G71gat), .B(G99gat), .ZN(new_n431));
  XOR2_X1   g230(.A(new_n430), .B(new_n431), .Z(new_n432));
  NAND4_X1  g231(.A1(new_n421), .A2(new_n422), .A3(new_n425), .A4(new_n423), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n433), .A2(KEYINPUT34), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n433), .A2(KEYINPUT34), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n429), .B(new_n432), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n427), .A2(KEYINPUT32), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n421), .A2(new_n423), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT34), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n439), .A2(new_n440), .A3(new_n425), .A4(new_n422), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n433), .A2(KEYINPUT34), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT33), .B1(new_n424), .B2(new_n426), .ZN(new_n443));
  INV_X1    g242(.A(new_n432), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n441), .B(new_n442), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n436), .A2(new_n438), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n438), .B1(new_n436), .B2(new_n445), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(KEYINPUT36), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n436), .A2(new_n445), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n437), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n436), .A2(new_n445), .A3(new_n438), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT36), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n449), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n410), .A2(new_n413), .ZN(new_n457));
  INV_X1    g256(.A(new_n414), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n410), .A2(new_n413), .A3(new_n414), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OR2_X1    g260(.A1(new_n357), .A2(new_n286), .ZN(new_n462));
  OR2_X1    g261(.A1(new_n462), .A2(KEYINPUT39), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n351), .A2(new_n286), .A3(new_n352), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(KEYINPUT39), .A3(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n360), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT40), .ZN(new_n467));
  OR2_X1    g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n278), .A2(new_n375), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n466), .A2(new_n467), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n468), .A2(new_n470), .A3(new_n359), .A4(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT37), .B1(new_n275), .B2(new_n276), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n473), .A2(new_n205), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n275), .A2(KEYINPUT37), .A3(new_n276), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT79), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n473), .A2(new_n477), .A3(new_n205), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n476), .B1(KEYINPUT38), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n379), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n374), .A2(new_n205), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT38), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n474), .A2(new_n477), .A3(new_n482), .A4(new_n475), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n479), .A2(new_n480), .A3(new_n481), .A4(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n461), .A2(new_n472), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n418), .A2(new_n456), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT35), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n378), .A2(new_n382), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n453), .B1(new_n460), .B2(new_n459), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT80), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n491), .B1(new_n446), .B2(new_n447), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n451), .A2(KEYINPUT80), .A3(new_n452), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n492), .A2(new_n493), .A3(new_n469), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n480), .A2(KEYINPUT35), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NOR3_X1   g295(.A1(new_n494), .A2(new_n417), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n486), .B1(new_n490), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT82), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  OR3_X1    g300(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G43gat), .B(G50gat), .ZN(new_n504));
  OR3_X1    g303(.A1(new_n504), .A2(KEYINPUT86), .A3(KEYINPUT15), .ZN(new_n505));
  XNOR2_X1  g304(.A(KEYINPUT85), .B(G36gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(G29gat), .ZN(new_n507));
  OAI21_X1  g306(.A(KEYINPUT15), .B1(new_n504), .B2(KEYINPUT86), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n503), .A2(new_n505), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n501), .A2(KEYINPUT83), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n499), .B(KEYINPUT82), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT83), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n502), .B(KEYINPUT84), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n510), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n515), .A2(new_n507), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n504), .A2(KEYINPUT15), .ZN(new_n517));
  OAI211_X1 g316(.A(KEYINPUT17), .B(new_n509), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G15gat), .B(G22gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT87), .B(G1gat), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT16), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n522), .B(KEYINPUT88), .C1(G1gat), .C2(new_n519), .ZN(new_n523));
  INV_X1    g322(.A(G8gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n523), .B(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT17), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n517), .B1(new_n515), .B2(new_n507), .ZN(new_n527));
  INV_X1    g326(.A(new_n509), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n518), .A2(new_n525), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n509), .B1(new_n516), .B2(new_n517), .ZN(new_n531));
  INV_X1    g330(.A(new_n525), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(KEYINPUT89), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n530), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT18), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n535), .B(KEYINPUT13), .Z(new_n539));
  INV_X1    g338(.A(new_n533), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n531), .A2(new_n532), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n530), .A2(KEYINPUT18), .A3(new_n533), .A4(new_n535), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n538), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(KEYINPUT81), .B(KEYINPUT11), .Z(new_n545));
  XNOR2_X1  g344(.A(G113gat), .B(G141gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G169gat), .B(G197gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT12), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n544), .A2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT90), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n538), .A2(new_n550), .A3(new_n542), .A4(new_n543), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n552), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n544), .A2(KEYINPUT90), .A3(new_n551), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n498), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(G71gat), .A2(G78gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT91), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT9), .ZN(new_n561));
  XNOR2_X1  g360(.A(G57gat), .B(G64gat), .ZN(new_n562));
  INV_X1    g361(.A(G71gat), .ZN(new_n563));
  INV_X1    g362(.A(G78gat), .ZN(new_n564));
  OAI221_X1 g363(.A(new_n560), .B1(new_n561), .B2(new_n562), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n563), .A2(new_n564), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n566), .B1(KEYINPUT9), .B2(new_n559), .ZN(new_n567));
  OR2_X1    g366(.A1(new_n567), .A2(new_n562), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n565), .A2(KEYINPUT21), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n525), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT92), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n565), .A2(new_n568), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT21), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(G183gat), .B(G211gat), .Z(new_n577));
  XOR2_X1   g376(.A(new_n576), .B(new_n577), .Z(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n572), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n571), .B(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(new_n578), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G127gat), .B(G155gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n585), .B(new_n586), .Z(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n580), .A2(new_n583), .A3(new_n587), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G99gat), .A2(G106gat), .ZN(new_n592));
  INV_X1    g391(.A(G92gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(KEYINPUT8), .A2(new_n592), .B1(new_n282), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT7), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n595), .B1(new_n282), .B2(new_n593), .ZN(new_n596));
  NAND3_X1  g395(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n594), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G99gat), .B(G106gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  AND2_X1   g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601));
  AOI22_X1  g400(.A1(new_n531), .A2(new_n600), .B1(KEYINPUT41), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n600), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n518), .A2(new_n529), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G190gat), .B(G218gat), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n602), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n605), .B1(new_n602), .B2(new_n604), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT94), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT94), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n610), .B1(new_n606), .B2(new_n607), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n601), .A2(KEYINPUT41), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT93), .ZN(new_n613));
  XNOR2_X1  g412(.A(G134gat), .B(G162gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n609), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n615), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n608), .A2(KEYINPUT94), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n591), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT95), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n591), .A2(KEYINPUT95), .A3(new_n619), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n603), .A2(new_n574), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT10), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n600), .A2(new_n568), .A3(new_n565), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n626), .A2(new_n625), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(G230gat), .A2(G233gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(new_n624), .A2(new_n626), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(new_n630), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n631), .B1(new_n634), .B2(KEYINPUT96), .ZN(new_n635));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(G176gat), .B(G204gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT96), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n639), .B1(new_n633), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n630), .B(KEYINPUT97), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n645), .B1(new_n627), .B2(new_n628), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n638), .B1(new_n646), .B2(new_n633), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n622), .A2(new_n623), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n558), .A2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n379), .B(KEYINPUT98), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g455(.A1(new_n652), .A2(new_n469), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT42), .B1(new_n657), .B2(new_n524), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT99), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G8gat), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  MUX2_X1   g460(.A(KEYINPUT42), .B(new_n658), .S(new_n661), .Z(G1325gat));
  INV_X1    g461(.A(G15gat), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n652), .A2(new_n663), .A3(new_n456), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n492), .A2(new_n493), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n653), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n664), .B1(new_n663), .B2(new_n666), .ZN(G1326gat));
  NAND2_X1  g466(.A1(new_n653), .A2(new_n417), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(G22gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT100), .B(KEYINPUT43), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(G1327gat));
  NOR2_X1   g470(.A1(new_n619), .A2(KEYINPUT107), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n673), .B1(new_n616), .B2(new_n618), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(KEYINPUT44), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n486), .A2(new_n677), .ZN(new_n678));
  AOI22_X1  g477(.A1(new_n383), .A2(new_n417), .B1(new_n449), .B2(new_n455), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(KEYINPUT104), .A3(new_n485), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n490), .B2(new_n497), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n665), .A2(new_n461), .A3(new_n495), .A4(new_n469), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n448), .B1(new_n415), .B2(new_n416), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT35), .B1(new_n383), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(KEYINPUT105), .A3(new_n686), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n681), .A2(KEYINPUT106), .A3(new_n683), .A4(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  AND3_X1   g488(.A1(new_n684), .A2(KEYINPUT105), .A3(new_n686), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT105), .B1(new_n684), .B2(new_n686), .ZN(new_n691));
  NOR2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(KEYINPUT106), .B1(new_n692), .B2(new_n681), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n676), .B1(new_n689), .B2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n619), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n498), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n696), .A2(KEYINPUT44), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n591), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n557), .A2(KEYINPUT102), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n555), .A2(new_n556), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT102), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n648), .B(KEYINPUT103), .Z(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n699), .A2(new_n700), .A3(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(new_n654), .ZN(new_n710));
  OAI21_X1  g509(.A(G29gat), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n700), .A2(new_n695), .A3(new_n649), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n558), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n716), .A2(G29gat), .A3(new_n710), .ZN(new_n717));
  XOR2_X1   g516(.A(new_n717), .B(KEYINPUT45), .Z(new_n718));
  NAND2_X1  g517(.A1(new_n711), .A2(new_n718), .ZN(G1328gat));
  OAI21_X1  g518(.A(new_n506), .B1(new_n709), .B2(new_n469), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n716), .A2(new_n469), .A3(new_n506), .ZN(new_n721));
  XNOR2_X1  g520(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(G1329gat));
  INV_X1    g523(.A(new_n709), .ZN(new_n725));
  INV_X1    g524(.A(new_n456), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n725), .A2(G43gat), .A3(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(G43gat), .ZN(new_n728));
  INV_X1    g527(.A(new_n665), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n716), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n731));
  AND3_X1   g530(.A1(new_n727), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n731), .B1(new_n727), .B2(new_n730), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(G1330gat));
  NAND3_X1  g533(.A1(new_n725), .A2(G50gat), .A3(new_n417), .ZN(new_n735));
  INV_X1    g534(.A(new_n716), .ZN(new_n736));
  AOI21_X1  g535(.A(G50gat), .B1(new_n736), .B2(new_n417), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT48), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT48), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n735), .A2(new_n741), .A3(new_n738), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(G1331gat));
  AND4_X1   g542(.A1(KEYINPUT104), .A2(new_n418), .A3(new_n456), .A4(new_n485), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT104), .B1(new_n679), .B2(new_n485), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n683), .B(new_n687), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n688), .ZN(new_n749));
  AND4_X1   g548(.A1(new_n622), .A2(new_n706), .A3(new_n623), .A4(new_n707), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(new_n710), .ZN(new_n752));
  XNOR2_X1  g551(.A(KEYINPUT110), .B(G57gat), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1332gat));
  NOR2_X1   g553(.A1(new_n751), .A2(new_n469), .ZN(new_n755));
  NOR2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  AND2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(new_n755), .B2(new_n756), .ZN(G1333gat));
  OAI21_X1  g558(.A(new_n563), .B1(new_n751), .B2(new_n729), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n749), .A2(G71gat), .A3(new_n726), .A4(new_n750), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g562(.A1(new_n751), .A2(new_n461), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(new_n564), .ZN(G1335gat));
  INV_X1    g564(.A(KEYINPUT111), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n706), .A2(new_n700), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n699), .A2(new_n766), .A3(new_n648), .A4(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n676), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n748), .B2(new_n688), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n648), .B(new_n768), .C1(new_n771), .C2(new_n697), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT111), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n282), .B1(new_n774), .B2(new_n654), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n746), .A2(new_n695), .A3(new_n768), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(KEYINPUT51), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n777), .A2(new_n649), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n778), .A2(new_n282), .A3(new_n654), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT112), .B1(new_n775), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n710), .B1(new_n769), .B2(new_n773), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n782), .B(new_n779), .C1(new_n783), .C2(new_n282), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n781), .A2(new_n784), .ZN(G1336gat));
  INV_X1    g584(.A(new_n707), .ZN(new_n786));
  NOR4_X1   g585(.A1(new_n777), .A2(G92gat), .A3(new_n469), .A4(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(G92gat), .B1(new_n772), .B2(new_n469), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT52), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n769), .A2(new_n773), .ZN(new_n792));
  OAI211_X1 g591(.A(KEYINPUT52), .B(G92gat), .C1(new_n792), .C2(new_n469), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT52), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n787), .B1(new_n788), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n791), .B1(new_n793), .B2(new_n795), .ZN(G1337gat));
  OAI21_X1  g595(.A(G99gat), .B1(new_n792), .B2(new_n456), .ZN(new_n797));
  INV_X1    g596(.A(G99gat), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n778), .A2(new_n798), .A3(new_n665), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1338gat));
  NOR4_X1   g599(.A1(new_n777), .A2(G106gat), .A3(new_n461), .A4(new_n786), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n801), .A2(KEYINPUT53), .ZN(new_n802));
  OAI21_X1  g601(.A(G106gat), .B1(new_n772), .B2(new_n461), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n774), .A2(new_n417), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n801), .B1(new_n805), .B2(G106gat), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n804), .B1(new_n806), .B2(new_n807), .ZN(G1339gat));
  NAND3_X1  g607(.A1(new_n627), .A2(new_n628), .A3(new_n645), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n631), .A2(KEYINPUT54), .A3(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT54), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n639), .B1(new_n646), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(KEYINPUT55), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n810), .A2(new_n815), .A3(new_n812), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n642), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n540), .A2(new_n541), .A3(new_n539), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n535), .B1(new_n530), .B2(new_n533), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n549), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n817), .A2(new_n554), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n821), .B1(new_n672), .B2(new_n674), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n648), .A2(new_n554), .A3(new_n820), .ZN(new_n823));
  INV_X1    g622(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n824), .B1(new_n705), .B2(new_n817), .ZN(new_n825));
  INV_X1    g624(.A(new_n675), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n822), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  AOI22_X1  g626(.A1(new_n827), .A2(new_n700), .B1(new_n651), .B2(new_n706), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(new_n710), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n665), .A2(new_n461), .A3(new_n469), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(G113gat), .B1(new_n832), .B2(new_n702), .ZN(new_n833));
  NOR4_X1   g632(.A1(new_n828), .A2(new_n685), .A3(new_n470), .A4(new_n710), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n290), .A3(new_n705), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(G1340gat));
  NOR3_X1   g635(.A1(new_n832), .A2(new_n293), .A3(new_n786), .ZN(new_n837));
  AOI21_X1  g636(.A(G120gat), .B1(new_n834), .B2(new_n648), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT114), .ZN(G1341gat));
  NOR3_X1   g639(.A1(new_n832), .A2(new_n298), .A3(new_n700), .ZN(new_n841));
  AOI21_X1  g640(.A(G127gat), .B1(new_n834), .B2(new_n591), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(G1342gat));
  NAND3_X1  g642(.A1(new_n834), .A2(new_n299), .A3(new_n695), .ZN(new_n844));
  XOR2_X1   g643(.A(new_n844), .B(KEYINPUT56), .Z(new_n845));
  OAI21_X1  g644(.A(G134gat), .B1(new_n832), .B2(new_n619), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1343gat));
  NAND3_X1  g646(.A1(new_n555), .A2(new_n556), .A3(new_n817), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n823), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(KEYINPUT115), .A3(new_n619), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n822), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT115), .B1(new_n849), .B2(new_n619), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n700), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT116), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n651), .A2(new_n706), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n856), .B(new_n700), .C1(new_n851), .C2(new_n852), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n854), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n461), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n859), .B1(new_n828), .B2(new_n461), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n858), .A2(KEYINPUT117), .A3(new_n860), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n726), .A2(new_n470), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n868), .A2(new_n710), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n866), .A2(new_n557), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n339), .ZN(new_n871));
  NOR4_X1   g670(.A1(new_n828), .A2(new_n461), .A3(new_n710), .A4(new_n868), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n702), .A2(G141gat), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(KEYINPUT58), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n866), .A2(new_n705), .A3(new_n869), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n874), .B1(new_n878), .B2(new_n339), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n876), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT118), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n876), .B(KEYINPUT118), .C1(new_n877), .C2(new_n879), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(G1344gat));
  INV_X1    g683(.A(new_n338), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n872), .A2(new_n885), .A3(new_n648), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n886), .B(KEYINPUT119), .Z(new_n887));
  NAND2_X1  g686(.A1(new_n827), .A2(new_n700), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n855), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n889), .A2(KEYINPUT57), .A3(new_n417), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n695), .B1(new_n823), .B2(new_n848), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n821), .A2(new_n695), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n700), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n893), .B1(new_n650), .B2(new_n557), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT57), .B1(new_n894), .B2(new_n417), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n895), .A2(KEYINPUT121), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(KEYINPUT121), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n890), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n649), .B1(new_n869), .B2(KEYINPUT120), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n898), .B(new_n899), .C1(KEYINPUT120), .C2(new_n869), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n866), .A2(new_n869), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n885), .B1(new_n902), .B2(new_n648), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n887), .B(new_n901), .C1(new_n903), .C2(KEYINPUT59), .ZN(G1345gat));
  NAND2_X1  g703(.A1(new_n872), .A2(new_n591), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT122), .ZN(new_n906));
  INV_X1    g705(.A(G155gat), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n700), .A2(new_n907), .ZN(new_n908));
  AOI22_X1  g707(.A1(new_n906), .A2(new_n907), .B1(new_n902), .B2(new_n908), .ZN(G1346gat));
  AOI21_X1  g708(.A(G162gat), .B1(new_n872), .B2(new_n695), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n902), .A2(new_n826), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n911), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g711(.A1(new_n654), .A2(new_n469), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n889), .A2(new_n489), .A3(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(new_n213), .A3(new_n705), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n889), .A2(new_n461), .A3(new_n665), .A4(new_n913), .ZN(new_n917));
  OAI21_X1  g716(.A(G169gat), .B1(new_n917), .B2(new_n702), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(G1348gat));
  AOI21_X1  g718(.A(G176gat), .B1(new_n915), .B2(new_n648), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n917), .A2(new_n214), .A3(new_n786), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n920), .A2(new_n921), .ZN(G1349gat));
  NAND3_X1  g721(.A1(new_n915), .A2(new_n245), .A3(new_n591), .ZN(new_n923));
  OAI21_X1  g722(.A(G183gat), .B1(new_n917), .B2(new_n700), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g724(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n925), .B(new_n926), .ZN(G1350gat));
  OAI21_X1  g726(.A(G190gat), .B1(new_n917), .B2(new_n619), .ZN(new_n928));
  XOR2_X1   g727(.A(KEYINPUT124), .B(KEYINPUT61), .Z(new_n929));
  XNOR2_X1  g728(.A(new_n928), .B(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n915), .A2(new_n236), .A3(new_n826), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1351gat));
  NAND2_X1  g731(.A1(new_n898), .A2(KEYINPUT125), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n456), .A2(new_n913), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n890), .A2(new_n896), .A3(new_n936), .A4(new_n897), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n933), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g737(.A(G197gat), .B1(new_n938), .B2(new_n702), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n828), .A2(new_n461), .A3(new_n934), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n706), .A2(G197gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(G1352gat));
  OAI21_X1  g742(.A(G204gat), .B1(new_n938), .B2(new_n786), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n941), .A2(G204gat), .A3(new_n649), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT62), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT126), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT126), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n944), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1353gat));
  NAND3_X1  g750(.A1(new_n940), .A2(new_n258), .A3(new_n591), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n898), .A2(new_n591), .A3(new_n935), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n953), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n954));
  AOI21_X1  g753(.A(KEYINPUT63), .B1(new_n953), .B2(G211gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(G1354gat));
  NAND3_X1  g755(.A1(new_n940), .A2(new_n259), .A3(new_n826), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT127), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n938), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n933), .A2(KEYINPUT127), .A3(new_n935), .A4(new_n937), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n959), .A2(new_n695), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n957), .B1(new_n961), .B2(new_n259), .ZN(G1355gat));
endmodule


