

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U562 ( .A(KEYINPUT27), .ZN(n718) );
  XNOR2_X1 U563 ( .A(n719), .B(n718), .ZN(n722) );
  OR2_X1 U564 ( .A1(n712), .A2(n711), .ZN(n760) );
  NOR2_X1 U565 ( .A1(G651), .A2(n635), .ZN(n657) );
  INV_X1 U566 ( .A(G2105), .ZN(n528) );
  AND2_X1 U567 ( .A1(n528), .A2(G2104), .ZN(n898) );
  NAND2_X1 U568 ( .A1(G101), .A2(n898), .ZN(n527) );
  XNOR2_X1 U569 ( .A(n527), .B(KEYINPUT23), .ZN(n531) );
  NOR2_X4 U570 ( .A1(G2104), .A2(n528), .ZN(n894) );
  NAND2_X1 U571 ( .A1(G125), .A2(n894), .ZN(n529) );
  XOR2_X1 U572 ( .A(KEYINPUT64), .B(n529), .Z(n530) );
  NOR2_X1 U573 ( .A1(n531), .A2(n530), .ZN(n534) );
  NOR2_X1 U574 ( .A1(G2104), .A2(G2105), .ZN(n532) );
  XOR2_X2 U575 ( .A(KEYINPUT17), .B(n532), .Z(n897) );
  NAND2_X1 U576 ( .A1(n897), .A2(G137), .ZN(n533) );
  NAND2_X1 U577 ( .A1(n534), .A2(n533), .ZN(n537) );
  AND2_X1 U578 ( .A1(G2104), .A2(G2105), .ZN(n893) );
  NAND2_X1 U579 ( .A1(G113), .A2(n893), .ZN(n535) );
  XNOR2_X1 U580 ( .A(KEYINPUT65), .B(n535), .ZN(n536) );
  NOR2_X2 U581 ( .A1(n537), .A2(n536), .ZN(G160) );
  NOR2_X1 U582 ( .A1(G651), .A2(G543), .ZN(n650) );
  NAND2_X1 U583 ( .A1(n650), .A2(G89), .ZN(n538) );
  XNOR2_X1 U584 ( .A(n538), .B(KEYINPUT4), .ZN(n541) );
  XNOR2_X1 U585 ( .A(G543), .B(KEYINPUT0), .ZN(n539) );
  XNOR2_X1 U586 ( .A(n539), .B(KEYINPUT67), .ZN(n635) );
  XOR2_X1 U587 ( .A(G651), .B(KEYINPUT68), .Z(n543) );
  NOR2_X1 U588 ( .A1(n635), .A2(n543), .ZN(n652) );
  NAND2_X1 U589 ( .A1(G76), .A2(n652), .ZN(n540) );
  NAND2_X1 U590 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U591 ( .A(n542), .B(KEYINPUT5), .ZN(n549) );
  NAND2_X1 U592 ( .A1(n657), .A2(G51), .ZN(n546) );
  NOR2_X1 U593 ( .A1(G543), .A2(n543), .ZN(n544) );
  XOR2_X1 U594 ( .A(KEYINPUT1), .B(n544), .Z(n656) );
  NAND2_X1 U595 ( .A1(G63), .A2(n656), .ZN(n545) );
  NAND2_X1 U596 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U597 ( .A(KEYINPUT6), .B(n547), .Z(n548) );
  NAND2_X1 U598 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U599 ( .A(n550), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U600 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U601 ( .A(G2438), .B(G2454), .Z(n552) );
  XNOR2_X1 U602 ( .A(G2435), .B(G2430), .ZN(n551) );
  XNOR2_X1 U603 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U604 ( .A(n553), .B(KEYINPUT106), .Z(n555) );
  XNOR2_X1 U605 ( .A(G1341), .B(G1348), .ZN(n554) );
  XNOR2_X1 U606 ( .A(n555), .B(n554), .ZN(n559) );
  XOR2_X1 U607 ( .A(G2446), .B(G2451), .Z(n557) );
  XNOR2_X1 U608 ( .A(G2443), .B(G2427), .ZN(n556) );
  XNOR2_X1 U609 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U610 ( .A(n559), .B(n558), .Z(n560) );
  AND2_X1 U611 ( .A1(G14), .A2(n560), .ZN(G401) );
  AND2_X1 U612 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U613 ( .A(G132), .ZN(G219) );
  INV_X1 U614 ( .A(G82), .ZN(G220) );
  NAND2_X1 U615 ( .A1(n657), .A2(G52), .ZN(n562) );
  NAND2_X1 U616 ( .A1(G64), .A2(n656), .ZN(n561) );
  NAND2_X1 U617 ( .A1(n562), .A2(n561), .ZN(n567) );
  NAND2_X1 U618 ( .A1(n650), .A2(G90), .ZN(n564) );
  NAND2_X1 U619 ( .A1(G77), .A2(n652), .ZN(n563) );
  NAND2_X1 U620 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U621 ( .A(KEYINPUT9), .B(n565), .Z(n566) );
  NOR2_X1 U622 ( .A1(n567), .A2(n566), .ZN(G171) );
  INV_X1 U623 ( .A(G171), .ZN(G301) );
  NAND2_X1 U624 ( .A1(G7), .A2(G661), .ZN(n568) );
  XOR2_X1 U625 ( .A(n568), .B(KEYINPUT10), .Z(n918) );
  NAND2_X1 U626 ( .A1(n918), .A2(G567), .ZN(n569) );
  XOR2_X1 U627 ( .A(KEYINPUT11), .B(n569), .Z(G234) );
  XOR2_X1 U628 ( .A(KEYINPUT14), .B(KEYINPUT72), .Z(n571) );
  NAND2_X1 U629 ( .A1(G56), .A2(n656), .ZN(n570) );
  XNOR2_X1 U630 ( .A(n571), .B(n570), .ZN(n578) );
  NAND2_X1 U631 ( .A1(n650), .A2(G81), .ZN(n572) );
  XNOR2_X1 U632 ( .A(n572), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U633 ( .A1(G68), .A2(n652), .ZN(n573) );
  NAND2_X1 U634 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U635 ( .A(n575), .B(KEYINPUT73), .ZN(n576) );
  XNOR2_X1 U636 ( .A(KEYINPUT13), .B(n576), .ZN(n577) );
  NOR2_X1 U637 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U638 ( .A(n579), .B(KEYINPUT74), .ZN(n581) );
  NAND2_X1 U639 ( .A1(G43), .A2(n657), .ZN(n580) );
  NAND2_X1 U640 ( .A1(n581), .A2(n580), .ZN(n985) );
  INV_X1 U641 ( .A(G860), .ZN(n601) );
  OR2_X1 U642 ( .A1(n985), .A2(n601), .ZN(G153) );
  NAND2_X1 U643 ( .A1(G868), .A2(G301), .ZN(n591) );
  NAND2_X1 U644 ( .A1(G54), .A2(n657), .ZN(n588) );
  NAND2_X1 U645 ( .A1(G79), .A2(n652), .ZN(n583) );
  NAND2_X1 U646 ( .A1(G66), .A2(n656), .ZN(n582) );
  NAND2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U648 ( .A1(G92), .A2(n650), .ZN(n584) );
  XNOR2_X1 U649 ( .A(KEYINPUT75), .B(n584), .ZN(n585) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U651 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U652 ( .A(n589), .B(KEYINPUT15), .ZN(n974) );
  OR2_X1 U653 ( .A1(n974), .A2(G868), .ZN(n590) );
  NAND2_X1 U654 ( .A1(n591), .A2(n590), .ZN(G284) );
  NAND2_X1 U655 ( .A1(G91), .A2(n650), .ZN(n593) );
  NAND2_X1 U656 ( .A1(G53), .A2(n657), .ZN(n592) );
  NAND2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n596) );
  NAND2_X1 U658 ( .A1(n652), .A2(G78), .ZN(n594) );
  XOR2_X1 U659 ( .A(KEYINPUT70), .B(n594), .Z(n595) );
  NOR2_X1 U660 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U661 ( .A1(G65), .A2(n656), .ZN(n597) );
  NAND2_X1 U662 ( .A1(n598), .A2(n597), .ZN(G299) );
  NOR2_X1 U663 ( .A1(G868), .A2(G299), .ZN(n600) );
  INV_X1 U664 ( .A(G868), .ZN(n671) );
  NOR2_X1 U665 ( .A1(G286), .A2(n671), .ZN(n599) );
  NOR2_X1 U666 ( .A1(n600), .A2(n599), .ZN(G297) );
  NAND2_X1 U667 ( .A1(n601), .A2(G559), .ZN(n602) );
  NAND2_X1 U668 ( .A1(n602), .A2(n974), .ZN(n603) );
  XNOR2_X1 U669 ( .A(n603), .B(KEYINPUT76), .ZN(n604) );
  XNOR2_X1 U670 ( .A(KEYINPUT16), .B(n604), .ZN(G148) );
  NAND2_X1 U671 ( .A1(n974), .A2(G868), .ZN(n605) );
  XOR2_X1 U672 ( .A(KEYINPUT77), .B(n605), .Z(n606) );
  NOR2_X1 U673 ( .A1(G559), .A2(n606), .ZN(n608) );
  NOR2_X1 U674 ( .A1(G868), .A2(n985), .ZN(n607) );
  NOR2_X1 U675 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U676 ( .A1(G123), .A2(n894), .ZN(n609) );
  XNOR2_X1 U677 ( .A(n609), .B(KEYINPUT18), .ZN(n611) );
  NAND2_X1 U678 ( .A1(n893), .A2(G111), .ZN(n610) );
  NAND2_X1 U679 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U680 ( .A1(G135), .A2(n897), .ZN(n613) );
  NAND2_X1 U681 ( .A1(G99), .A2(n898), .ZN(n612) );
  NAND2_X1 U682 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U683 ( .A1(n615), .A2(n614), .ZN(n942) );
  XNOR2_X1 U684 ( .A(G2096), .B(n942), .ZN(n616) );
  INV_X1 U685 ( .A(G2100), .ZN(n854) );
  NAND2_X1 U686 ( .A1(n616), .A2(n854), .ZN(G156) );
  NAND2_X1 U687 ( .A1(n974), .A2(G559), .ZN(n668) );
  XNOR2_X1 U688 ( .A(n985), .B(n668), .ZN(n617) );
  NOR2_X1 U689 ( .A1(n617), .A2(G860), .ZN(n625) );
  NAND2_X1 U690 ( .A1(G67), .A2(n656), .ZN(n618) );
  XNOR2_X1 U691 ( .A(n618), .B(KEYINPUT78), .ZN(n620) );
  NAND2_X1 U692 ( .A1(G93), .A2(n650), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n624) );
  NAND2_X1 U694 ( .A1(n657), .A2(G55), .ZN(n622) );
  NAND2_X1 U695 ( .A1(G80), .A2(n652), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n622), .A2(n621), .ZN(n623) );
  OR2_X1 U697 ( .A1(n624), .A2(n623), .ZN(n670) );
  XOR2_X1 U698 ( .A(n625), .B(n670), .Z(G145) );
  NAND2_X1 U699 ( .A1(n657), .A2(G48), .ZN(n626) );
  XNOR2_X1 U700 ( .A(KEYINPUT82), .B(n626), .ZN(n634) );
  NAND2_X1 U701 ( .A1(n650), .A2(G86), .ZN(n628) );
  NAND2_X1 U702 ( .A1(G61), .A2(n656), .ZN(n627) );
  NAND2_X1 U703 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U704 ( .A1(G73), .A2(n652), .ZN(n629) );
  XOR2_X1 U705 ( .A(KEYINPUT2), .B(n629), .Z(n630) );
  NOR2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U707 ( .A(KEYINPUT81), .B(n632), .Z(n633) );
  NAND2_X1 U708 ( .A1(n634), .A2(n633), .ZN(G305) );
  NAND2_X1 U709 ( .A1(G87), .A2(n635), .ZN(n641) );
  NAND2_X1 U710 ( .A1(G49), .A2(n657), .ZN(n637) );
  NAND2_X1 U711 ( .A1(G74), .A2(G651), .ZN(n636) );
  NAND2_X1 U712 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U713 ( .A1(n656), .A2(n638), .ZN(n639) );
  XOR2_X1 U714 ( .A(KEYINPUT79), .B(n639), .Z(n640) );
  NAND2_X1 U715 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U716 ( .A(n642), .B(KEYINPUT80), .ZN(G288) );
  NAND2_X1 U717 ( .A1(G88), .A2(n650), .ZN(n644) );
  NAND2_X1 U718 ( .A1(G50), .A2(n657), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U720 ( .A1(G75), .A2(n652), .ZN(n645) );
  XNOR2_X1 U721 ( .A(KEYINPUT83), .B(n645), .ZN(n646) );
  NOR2_X1 U722 ( .A1(n647), .A2(n646), .ZN(n649) );
  NAND2_X1 U723 ( .A1(G62), .A2(n656), .ZN(n648) );
  NAND2_X1 U724 ( .A1(n649), .A2(n648), .ZN(G303) );
  NAND2_X1 U725 ( .A1(n650), .A2(G85), .ZN(n651) );
  XNOR2_X1 U726 ( .A(n651), .B(KEYINPUT66), .ZN(n654) );
  NAND2_X1 U727 ( .A1(G72), .A2(n652), .ZN(n653) );
  NAND2_X1 U728 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U729 ( .A(KEYINPUT69), .B(n655), .ZN(n661) );
  NAND2_X1 U730 ( .A1(n656), .A2(G60), .ZN(n659) );
  NAND2_X1 U731 ( .A1(n657), .A2(G47), .ZN(n658) );
  AND2_X1 U732 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U733 ( .A1(n661), .A2(n660), .ZN(G290) );
  XNOR2_X1 U734 ( .A(G305), .B(G288), .ZN(n663) );
  INV_X1 U735 ( .A(G299), .ZN(n980) );
  XOR2_X1 U736 ( .A(G303), .B(n980), .Z(n662) );
  XNOR2_X1 U737 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U738 ( .A(n664), .B(n985), .ZN(n667) );
  XOR2_X1 U739 ( .A(n670), .B(KEYINPUT19), .Z(n665) );
  XNOR2_X1 U740 ( .A(n665), .B(G290), .ZN(n666) );
  XNOR2_X1 U741 ( .A(n667), .B(n666), .ZN(n845) );
  XNOR2_X1 U742 ( .A(n668), .B(n845), .ZN(n669) );
  NAND2_X1 U743 ( .A1(n669), .A2(G868), .ZN(n673) );
  NAND2_X1 U744 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U745 ( .A1(n673), .A2(n672), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n675) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n674) );
  XNOR2_X1 U748 ( .A(n675), .B(n674), .ZN(n676) );
  NAND2_X1 U749 ( .A1(n676), .A2(G2090), .ZN(n677) );
  XOR2_X1 U750 ( .A(KEYINPUT21), .B(n677), .Z(n678) );
  XNOR2_X1 U751 ( .A(KEYINPUT85), .B(n678), .ZN(n679) );
  NAND2_X1 U752 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U753 ( .A(KEYINPUT71), .B(G57), .ZN(G237) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U755 ( .A1(G69), .A2(G120), .ZN(n680) );
  NOR2_X1 U756 ( .A1(G237), .A2(n680), .ZN(n681) );
  XNOR2_X1 U757 ( .A(KEYINPUT86), .B(n681), .ZN(n682) );
  NAND2_X1 U758 ( .A1(n682), .A2(G108), .ZN(n843) );
  NAND2_X1 U759 ( .A1(n843), .A2(G567), .ZN(n687) );
  NOR2_X1 U760 ( .A1(G220), .A2(G219), .ZN(n683) );
  XOR2_X1 U761 ( .A(KEYINPUT22), .B(n683), .Z(n684) );
  NOR2_X1 U762 ( .A1(G218), .A2(n684), .ZN(n685) );
  NAND2_X1 U763 ( .A1(G96), .A2(n685), .ZN(n844) );
  NAND2_X1 U764 ( .A1(n844), .A2(G2106), .ZN(n686) );
  NAND2_X1 U765 ( .A1(n687), .A2(n686), .ZN(n917) );
  NAND2_X1 U766 ( .A1(G661), .A2(G483), .ZN(n688) );
  NOR2_X1 U767 ( .A1(n917), .A2(n688), .ZN(n842) );
  NAND2_X1 U768 ( .A1(n842), .A2(G36), .ZN(G176) );
  NAND2_X1 U769 ( .A1(n897), .A2(G138), .ZN(n691) );
  NAND2_X1 U770 ( .A1(G114), .A2(n893), .ZN(n689) );
  XOR2_X1 U771 ( .A(KEYINPUT87), .B(n689), .Z(n690) );
  NAND2_X1 U772 ( .A1(n691), .A2(n690), .ZN(n695) );
  NAND2_X1 U773 ( .A1(G102), .A2(n898), .ZN(n693) );
  NAND2_X1 U774 ( .A1(G126), .A2(n894), .ZN(n692) );
  NAND2_X1 U775 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U776 ( .A1(n695), .A2(n694), .ZN(G164) );
  XNOR2_X1 U777 ( .A(G1986), .B(G290), .ZN(n977) );
  NOR2_X1 U778 ( .A1(G164), .A2(G1384), .ZN(n710) );
  NAND2_X1 U779 ( .A1(G160), .A2(G40), .ZN(n711) );
  NOR2_X1 U780 ( .A1(n710), .A2(n711), .ZN(n834) );
  NAND2_X1 U781 ( .A1(n977), .A2(n834), .ZN(n696) );
  XNOR2_X1 U782 ( .A(n696), .B(KEYINPUT88), .ZN(n709) );
  NAND2_X1 U783 ( .A1(G140), .A2(n897), .ZN(n698) );
  NAND2_X1 U784 ( .A1(G104), .A2(n898), .ZN(n697) );
  NAND2_X1 U785 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U786 ( .A(KEYINPUT34), .B(n699), .ZN(n705) );
  NAND2_X1 U787 ( .A1(n893), .A2(G116), .ZN(n700) );
  XNOR2_X1 U788 ( .A(n700), .B(KEYINPUT90), .ZN(n702) );
  NAND2_X1 U789 ( .A1(G128), .A2(n894), .ZN(n701) );
  NAND2_X1 U790 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U791 ( .A(n703), .B(KEYINPUT35), .Z(n704) );
  NOR2_X1 U792 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U793 ( .A(KEYINPUT36), .B(n706), .Z(n707) );
  XNOR2_X1 U794 ( .A(KEYINPUT91), .B(n707), .ZN(n890) );
  XOR2_X1 U795 ( .A(G2067), .B(KEYINPUT37), .Z(n708) );
  XNOR2_X1 U796 ( .A(KEYINPUT89), .B(n708), .ZN(n832) );
  NOR2_X1 U797 ( .A1(n890), .A2(n832), .ZN(n960) );
  NAND2_X1 U798 ( .A1(n834), .A2(n960), .ZN(n830) );
  NAND2_X1 U799 ( .A1(n709), .A2(n830), .ZN(n806) );
  INV_X1 U800 ( .A(n710), .ZN(n712) );
  NAND2_X1 U801 ( .A1(G8), .A2(n760), .ZN(n799) );
  NOR2_X1 U802 ( .A1(G1981), .A2(G305), .ZN(n713) );
  XOR2_X1 U803 ( .A(n713), .B(KEYINPUT24), .Z(n714) );
  NOR2_X1 U804 ( .A1(n799), .A2(n714), .ZN(n804) );
  XOR2_X1 U805 ( .A(KEYINPUT32), .B(KEYINPUT103), .Z(n768) );
  XOR2_X1 U806 ( .A(G2078), .B(KEYINPUT25), .Z(n922) );
  XOR2_X1 U807 ( .A(n760), .B(KEYINPUT95), .Z(n720) );
  NOR2_X1 U808 ( .A1(n922), .A2(n720), .ZN(n716) );
  INV_X1 U809 ( .A(n760), .ZN(n727) );
  NOR2_X1 U810 ( .A1(n727), .A2(G1961), .ZN(n715) );
  NOR2_X1 U811 ( .A1(n716), .A2(n715), .ZN(n749) );
  NOR2_X1 U812 ( .A1(n749), .A2(G301), .ZN(n717) );
  XOR2_X1 U813 ( .A(KEYINPUT96), .B(n717), .Z(n748) );
  INV_X1 U814 ( .A(n720), .ZN(n735) );
  NAND2_X1 U815 ( .A1(n735), .A2(G2072), .ZN(n719) );
  NAND2_X1 U816 ( .A1(n720), .A2(G1956), .ZN(n721) );
  NAND2_X1 U817 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U818 ( .A(n723), .B(KEYINPUT97), .ZN(n726) );
  NOR2_X1 U819 ( .A1(n726), .A2(n980), .ZN(n725) );
  XOR2_X1 U820 ( .A(KEYINPUT98), .B(KEYINPUT28), .Z(n724) );
  XNOR2_X1 U821 ( .A(n725), .B(n724), .ZN(n745) );
  NAND2_X1 U822 ( .A1(n726), .A2(n980), .ZN(n743) );
  AND2_X1 U823 ( .A1(n727), .A2(G1996), .ZN(n729) );
  XNOR2_X1 U824 ( .A(KEYINPUT26), .B(KEYINPUT99), .ZN(n728) );
  XNOR2_X1 U825 ( .A(n729), .B(n728), .ZN(n731) );
  NAND2_X1 U826 ( .A1(n760), .A2(G1341), .ZN(n730) );
  NAND2_X1 U827 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U828 ( .A1(n985), .A2(n732), .ZN(n734) );
  NOR2_X1 U829 ( .A1(n974), .A2(n734), .ZN(n733) );
  XOR2_X1 U830 ( .A(n733), .B(KEYINPUT100), .Z(n741) );
  NAND2_X1 U831 ( .A1(n974), .A2(n734), .ZN(n739) );
  NAND2_X1 U832 ( .A1(G2067), .A2(n735), .ZN(n737) );
  NAND2_X1 U833 ( .A1(G1348), .A2(n760), .ZN(n736) );
  NAND2_X1 U834 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U835 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U836 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U837 ( .A1(n743), .A2(n742), .ZN(n744) );
  NAND2_X1 U838 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U839 ( .A(KEYINPUT29), .B(n746), .Z(n747) );
  NAND2_X1 U840 ( .A1(n748), .A2(n747), .ZN(n759) );
  NAND2_X1 U841 ( .A1(n749), .A2(G301), .ZN(n750) );
  XNOR2_X1 U842 ( .A(n750), .B(KEYINPUT101), .ZN(n756) );
  NOR2_X1 U843 ( .A1(G2084), .A2(n760), .ZN(n772) );
  NOR2_X1 U844 ( .A1(G1966), .A2(n799), .ZN(n751) );
  XNOR2_X1 U845 ( .A(KEYINPUT94), .B(n751), .ZN(n770) );
  NOR2_X1 U846 ( .A1(n772), .A2(n770), .ZN(n752) );
  NAND2_X1 U847 ( .A1(G8), .A2(n752), .ZN(n753) );
  XNOR2_X1 U848 ( .A(KEYINPUT30), .B(n753), .ZN(n754) );
  NOR2_X1 U849 ( .A1(n754), .A2(G168), .ZN(n755) );
  NOR2_X1 U850 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U851 ( .A(KEYINPUT31), .B(n757), .Z(n758) );
  NAND2_X1 U852 ( .A1(n759), .A2(n758), .ZN(n769) );
  NAND2_X1 U853 ( .A1(n769), .A2(G286), .ZN(n765) );
  NOR2_X1 U854 ( .A1(G1971), .A2(n799), .ZN(n762) );
  NOR2_X1 U855 ( .A1(G2090), .A2(n760), .ZN(n761) );
  NOR2_X1 U856 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U857 ( .A1(n763), .A2(G303), .ZN(n764) );
  NAND2_X1 U858 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U859 ( .A1(n766), .A2(G8), .ZN(n767) );
  XNOR2_X1 U860 ( .A(n768), .B(n767), .ZN(n777) );
  INV_X1 U861 ( .A(n769), .ZN(n771) );
  NOR2_X1 U862 ( .A1(n771), .A2(n770), .ZN(n774) );
  NAND2_X1 U863 ( .A1(G8), .A2(n772), .ZN(n773) );
  NAND2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U865 ( .A(KEYINPUT102), .B(n775), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n798) );
  NOR2_X1 U867 ( .A1(G1971), .A2(G303), .ZN(n778) );
  XNOR2_X1 U868 ( .A(KEYINPUT104), .B(n778), .ZN(n779) );
  NOR2_X1 U869 ( .A1(KEYINPUT33), .A2(n779), .ZN(n780) );
  NAND2_X1 U870 ( .A1(n798), .A2(n780), .ZN(n783) );
  INV_X1 U871 ( .A(n799), .ZN(n781) );
  NAND2_X1 U872 ( .A1(n781), .A2(KEYINPUT105), .ZN(n782) );
  NAND2_X1 U873 ( .A1(n783), .A2(n782), .ZN(n784) );
  OR2_X1 U874 ( .A1(G288), .A2(G1976), .ZN(n787) );
  NAND2_X1 U875 ( .A1(n784), .A2(n787), .ZN(n795) );
  XNOR2_X1 U876 ( .A(G1981), .B(G305), .ZN(n971) );
  NAND2_X1 U877 ( .A1(G288), .A2(G1976), .ZN(n785) );
  NOR2_X1 U878 ( .A1(KEYINPUT105), .A2(n799), .ZN(n789) );
  NAND2_X1 U879 ( .A1(n785), .A2(n789), .ZN(n786) );
  INV_X1 U880 ( .A(KEYINPUT33), .ZN(n788) );
  NAND2_X1 U881 ( .A1(n786), .A2(n788), .ZN(n792) );
  NOR2_X1 U882 ( .A1(n788), .A2(n787), .ZN(n790) );
  NAND2_X1 U883 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U884 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U885 ( .A1(n971), .A2(n793), .ZN(n794) );
  NAND2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n802) );
  NOR2_X1 U887 ( .A1(G2090), .A2(G303), .ZN(n796) );
  NAND2_X1 U888 ( .A1(G8), .A2(n796), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n800) );
  NAND2_X1 U890 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n803) );
  NOR2_X1 U892 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U893 ( .A1(n806), .A2(n805), .ZN(n824) );
  NAND2_X1 U894 ( .A1(G131), .A2(n897), .ZN(n808) );
  NAND2_X1 U895 ( .A1(G119), .A2(n894), .ZN(n807) );
  NAND2_X1 U896 ( .A1(n808), .A2(n807), .ZN(n812) );
  NAND2_X1 U897 ( .A1(G107), .A2(n893), .ZN(n810) );
  NAND2_X1 U898 ( .A1(G95), .A2(n898), .ZN(n809) );
  NAND2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n811) );
  OR2_X1 U900 ( .A1(n812), .A2(n811), .ZN(n878) );
  NAND2_X1 U901 ( .A1(G1991), .A2(n878), .ZN(n821) );
  NAND2_X1 U902 ( .A1(G141), .A2(n897), .ZN(n814) );
  NAND2_X1 U903 ( .A1(G129), .A2(n894), .ZN(n813) );
  NAND2_X1 U904 ( .A1(n814), .A2(n813), .ZN(n817) );
  NAND2_X1 U905 ( .A1(n898), .A2(G105), .ZN(n815) );
  XOR2_X1 U906 ( .A(KEYINPUT38), .B(n815), .Z(n816) );
  NOR2_X1 U907 ( .A1(n817), .A2(n816), .ZN(n819) );
  NAND2_X1 U908 ( .A1(n893), .A2(G117), .ZN(n818) );
  NAND2_X1 U909 ( .A1(n819), .A2(n818), .ZN(n904) );
  NAND2_X1 U910 ( .A1(G1996), .A2(n904), .ZN(n820) );
  NAND2_X1 U911 ( .A1(n821), .A2(n820), .ZN(n947) );
  NAND2_X1 U912 ( .A1(n947), .A2(n834), .ZN(n822) );
  XOR2_X1 U913 ( .A(KEYINPUT92), .B(n822), .Z(n827) );
  XNOR2_X1 U914 ( .A(KEYINPUT93), .B(n827), .ZN(n823) );
  NAND2_X1 U915 ( .A1(n824), .A2(n823), .ZN(n837) );
  NOR2_X1 U916 ( .A1(G1996), .A2(n904), .ZN(n940) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n825) );
  NOR2_X1 U918 ( .A1(G1991), .A2(n878), .ZN(n943) );
  NOR2_X1 U919 ( .A1(n825), .A2(n943), .ZN(n826) );
  NOR2_X1 U920 ( .A1(n827), .A2(n826), .ZN(n828) );
  NOR2_X1 U921 ( .A1(n940), .A2(n828), .ZN(n829) );
  XNOR2_X1 U922 ( .A(n829), .B(KEYINPUT39), .ZN(n831) );
  NAND2_X1 U923 ( .A1(n831), .A2(n830), .ZN(n833) );
  NAND2_X1 U924 ( .A1(n890), .A2(n832), .ZN(n957) );
  NAND2_X1 U925 ( .A1(n833), .A2(n957), .ZN(n835) );
  NAND2_X1 U926 ( .A1(n835), .A2(n834), .ZN(n836) );
  NAND2_X1 U927 ( .A1(n837), .A2(n836), .ZN(n838) );
  XNOR2_X1 U928 ( .A(n838), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n918), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n839) );
  NAND2_X1 U931 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n840) );
  XOR2_X1 U933 ( .A(KEYINPUT107), .B(n840), .Z(n841) );
  NAND2_X1 U934 ( .A1(n842), .A2(n841), .ZN(G188) );
  XOR2_X1 U935 ( .A(G108), .B(KEYINPUT114), .Z(G238) );
  INV_X1 U937 ( .A(G120), .ZN(G236) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  INV_X1 U939 ( .A(G69), .ZN(G235) );
  NOR2_X1 U940 ( .A1(n844), .A2(n843), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U942 ( .A(n845), .B(G301), .ZN(n847) );
  XNOR2_X1 U943 ( .A(G286), .B(n974), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n848) );
  NOR2_X1 U945 ( .A1(G37), .A2(n848), .ZN(G397) );
  XOR2_X1 U946 ( .A(G2096), .B(KEYINPUT43), .Z(n850) );
  XNOR2_X1 U947 ( .A(G2090), .B(KEYINPUT108), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U949 ( .A(n851), .B(G2678), .Z(n853) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2072), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n858) );
  XNOR2_X1 U952 ( .A(KEYINPUT42), .B(n854), .ZN(n856) );
  XNOR2_X1 U953 ( .A(G2078), .B(G2084), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n857) );
  XNOR2_X1 U955 ( .A(n858), .B(n857), .ZN(G227) );
  XOR2_X1 U956 ( .A(G1961), .B(G1956), .Z(n860) );
  XNOR2_X1 U957 ( .A(G1986), .B(G1971), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U959 ( .A(n861), .B(G2474), .Z(n863) );
  XNOR2_X1 U960 ( .A(G1966), .B(G1981), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n867) );
  XOR2_X1 U962 ( .A(KEYINPUT41), .B(G1976), .Z(n865) );
  XNOR2_X1 U963 ( .A(G1996), .B(G1991), .ZN(n864) );
  XNOR2_X1 U964 ( .A(n865), .B(n864), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n867), .B(n866), .ZN(G229) );
  NAND2_X1 U966 ( .A1(G112), .A2(n893), .ZN(n868) );
  XNOR2_X1 U967 ( .A(n868), .B(KEYINPUT110), .ZN(n872) );
  XOR2_X1 U968 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n870) );
  NAND2_X1 U969 ( .A1(G124), .A2(n894), .ZN(n869) );
  XNOR2_X1 U970 ( .A(n870), .B(n869), .ZN(n871) );
  NAND2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n876) );
  NAND2_X1 U972 ( .A1(G136), .A2(n897), .ZN(n874) );
  NAND2_X1 U973 ( .A1(G100), .A2(n898), .ZN(n873) );
  NAND2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n875) );
  NOR2_X1 U975 ( .A1(n876), .A2(n875), .ZN(G162) );
  XOR2_X1 U976 ( .A(G164), .B(n942), .Z(n877) );
  XNOR2_X1 U977 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U978 ( .A(n879), .B(KEYINPUT48), .Z(n881) );
  XNOR2_X1 U979 ( .A(KEYINPUT111), .B(KEYINPUT46), .ZN(n880) );
  XNOR2_X1 U980 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U981 ( .A(G162), .B(n882), .ZN(n892) );
  NAND2_X1 U982 ( .A1(G139), .A2(n897), .ZN(n884) );
  NAND2_X1 U983 ( .A1(G103), .A2(n898), .ZN(n883) );
  NAND2_X1 U984 ( .A1(n884), .A2(n883), .ZN(n889) );
  NAND2_X1 U985 ( .A1(G115), .A2(n893), .ZN(n886) );
  NAND2_X1 U986 ( .A1(G127), .A2(n894), .ZN(n885) );
  NAND2_X1 U987 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n887), .Z(n888) );
  NOR2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n950) );
  XNOR2_X1 U990 ( .A(n890), .B(n950), .ZN(n891) );
  XNOR2_X1 U991 ( .A(n892), .B(n891), .ZN(n908) );
  NAND2_X1 U992 ( .A1(G118), .A2(n893), .ZN(n896) );
  NAND2_X1 U993 ( .A1(G130), .A2(n894), .ZN(n895) );
  NAND2_X1 U994 ( .A1(n896), .A2(n895), .ZN(n903) );
  NAND2_X1 U995 ( .A1(G142), .A2(n897), .ZN(n900) );
  NAND2_X1 U996 ( .A1(G106), .A2(n898), .ZN(n899) );
  NAND2_X1 U997 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U998 ( .A(n901), .B(KEYINPUT45), .Z(n902) );
  NOR2_X1 U999 ( .A1(n903), .A2(n902), .ZN(n905) );
  XNOR2_X1 U1000 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1001 ( .A(G160), .B(n906), .Z(n907) );
  XNOR2_X1 U1002 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n909), .ZN(G395) );
  NOR2_X1 U1004 ( .A1(G227), .A2(G229), .ZN(n910) );
  XOR2_X1 U1005 ( .A(KEYINPUT49), .B(n910), .Z(n911) );
  XNOR2_X1 U1006 ( .A(n911), .B(KEYINPUT113), .ZN(n912) );
  NOR2_X1 U1007 ( .A1(G397), .A2(n912), .ZN(n916) );
  NOR2_X1 U1008 ( .A1(n917), .A2(G401), .ZN(n913) );
  XOR2_X1 U1009 ( .A(KEYINPUT112), .B(n913), .Z(n914) );
  NOR2_X1 U1010 ( .A1(G395), .A2(n914), .ZN(n915) );
  NAND2_X1 U1011 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(n917), .ZN(G319) );
  INV_X1 U1014 ( .A(n918), .ZN(G223) );
  INV_X1 U1015 ( .A(G303), .ZN(G166) );
  XOR2_X1 U1016 ( .A(G29), .B(KEYINPUT118), .Z(n938) );
  XOR2_X1 U1017 ( .A(G2067), .B(G26), .Z(n919) );
  NAND2_X1 U1018 ( .A1(n919), .A2(G28), .ZN(n928) );
  XNOR2_X1 U1019 ( .A(G1996), .B(G32), .ZN(n921) );
  XNOR2_X1 U1020 ( .A(G33), .B(G2072), .ZN(n920) );
  NOR2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(G1991), .B(G25), .ZN(n924) );
  XNOR2_X1 U1023 ( .A(G27), .B(n922), .ZN(n923) );
  NOR2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1027 ( .A(KEYINPUT53), .B(n929), .Z(n932) );
  XOR2_X1 U1028 ( .A(G34), .B(KEYINPUT54), .Z(n930) );
  XNOR2_X1 U1029 ( .A(G2084), .B(n930), .ZN(n931) );
  NAND2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n935) );
  XOR2_X1 U1031 ( .A(KEYINPUT117), .B(G2090), .Z(n933) );
  XNOR2_X1 U1032 ( .A(G35), .B(n933), .ZN(n934) );
  NOR2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  INV_X1 U1034 ( .A(KEYINPUT55), .ZN(n964) );
  XOR2_X1 U1035 ( .A(n936), .B(n964), .Z(n937) );
  NAND2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n1023) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(KEYINPUT116), .ZN(n962) );
  XOR2_X1 U1038 ( .A(G2090), .B(G162), .Z(n939) );
  NOR2_X1 U1039 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1040 ( .A(KEYINPUT51), .B(n941), .Z(n949) );
  XNOR2_X1 U1041 ( .A(G160), .B(G2084), .ZN(n945) );
  NOR2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1043 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1045 ( .A1(n949), .A2(n948), .ZN(n956) );
  XNOR2_X1 U1046 ( .A(G2072), .B(n950), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(G164), .B(G2078), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1049 ( .A(KEYINPUT115), .B(n953), .Z(n954) );
  XNOR2_X1 U1050 ( .A(KEYINPUT50), .B(n954), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n958) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(n962), .B(n961), .ZN(n963) );
  NAND2_X1 U1055 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1056 ( .A1(n965), .A2(G29), .ZN(n966) );
  NAND2_X1 U1057 ( .A1(n966), .A2(G11), .ZN(n1021) );
  INV_X1 U1058 ( .A(G16), .ZN(n1016) );
  XOR2_X1 U1059 ( .A(n1016), .B(KEYINPUT56), .Z(n991) );
  XNOR2_X1 U1060 ( .A(G288), .B(KEYINPUT121), .ZN(n967) );
  XOR2_X1 U1061 ( .A(n967), .B(G1976), .Z(n969) );
  XOR2_X1 U1062 ( .A(G1961), .B(G171), .Z(n968) );
  NOR2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n989) );
  XOR2_X1 U1064 ( .A(G168), .B(G1966), .Z(n970) );
  NOR2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1066 ( .A(KEYINPUT57), .B(n972), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(n973), .B(KEYINPUT119), .ZN(n984) );
  XNOR2_X1 U1068 ( .A(G1348), .B(n974), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(n975), .B(KEYINPUT120), .ZN(n979) );
  XOR2_X1 U1070 ( .A(G1971), .B(G166), .Z(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n982) );
  XOR2_X1 U1073 ( .A(G1956), .B(n980), .Z(n981) );
  NOR2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(G1341), .B(n985), .ZN(n986) );
  NOR2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1078 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n1018) );
  XNOR2_X1 U1080 ( .A(G1961), .B(G5), .ZN(n1002) );
  XOR2_X1 U1081 ( .A(G1348), .B(KEYINPUT59), .Z(n992) );
  XNOR2_X1 U1082 ( .A(G4), .B(n992), .ZN(n994) );
  XNOR2_X1 U1083 ( .A(G20), .B(G1956), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n998) );
  XNOR2_X1 U1085 ( .A(G1341), .B(G19), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(G1981), .B(G6), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(n999), .B(KEYINPUT122), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(KEYINPUT60), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1010) );
  XOR2_X1 U1092 ( .A(G1986), .B(KEYINPUT123), .Z(n1003) );
  XNOR2_X1 U1093 ( .A(G24), .B(n1003), .ZN(n1007) );
  XOR2_X1 U1094 ( .A(G1971), .B(G22), .Z(n1005) );
  XOR2_X1 U1095 ( .A(G1976), .B(G23), .Z(n1004) );
  NAND2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(n1008), .B(KEYINPUT58), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(G21), .B(G1966), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(n1013), .B(KEYINPUT61), .ZN(n1014) );
  XNOR2_X1 U1103 ( .A(n1014), .B(KEYINPUT124), .ZN(n1015) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1106 ( .A(KEYINPUT125), .B(n1019), .Z(n1020) );
  NOR2_X1 U1107 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1109 ( .A(n1024), .B(KEYINPUT126), .ZN(n1025) );
  XOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1025), .Z(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

