//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 0 1 0 1 0 1 1 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT3), .B1(new_n190), .B2(G107), .ZN(new_n191));
  AOI21_X1  g005(.A(G101), .B1(new_n190), .B2(G107), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G104), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n192), .A3(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT82), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT82), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n191), .A2(new_n192), .A3(new_n195), .A4(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n194), .A2(G104), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n190), .A2(G107), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G101), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT1), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n210), .B1(G143), .B2(new_n205), .ZN(new_n211));
  INV_X1    g025(.A(G128), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n209), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(G143), .B(G146), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(new_n210), .A3(G128), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n200), .A2(new_n204), .A3(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT68), .B(G128), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n209), .B1(new_n218), .B2(new_n211), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n215), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n197), .A2(new_n199), .B1(G101), .B2(new_n203), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n217), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n223));
  INV_X1    g037(.A(G137), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G134), .ZN(new_n225));
  NOR2_X1   g039(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n223), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G131), .ZN(new_n228));
  INV_X1    g042(.A(G134), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G137), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n224), .A2(KEYINPUT64), .A3(KEYINPUT11), .A4(G134), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n227), .A2(new_n228), .A3(new_n230), .A4(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(KEYINPUT65), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n231), .A2(new_n230), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n234), .A2(new_n235), .A3(new_n228), .A4(new_n227), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(new_n227), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G131), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n222), .A2(KEYINPUT84), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT12), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT12), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n222), .A2(KEYINPUT84), .A3(new_n243), .A4(new_n240), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  XOR2_X1   g059(.A(KEYINPUT71), .B(G953), .Z(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G227), .ZN(new_n247));
  XOR2_X1   g061(.A(G110), .B(G140), .Z(new_n248));
  XNOR2_X1  g062(.A(new_n247), .B(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT10), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n217), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n191), .A2(new_n195), .A3(new_n202), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(G101), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n200), .A2(new_n254), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n253), .A2(new_n252), .A3(G101), .ZN(new_n256));
  NAND2_X1  g070(.A1(KEYINPUT0), .A2(G128), .ZN(new_n257));
  OR2_X1    g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n209), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n214), .A2(KEYINPUT0), .A3(G128), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n233), .A2(new_n236), .B1(G131), .B2(new_n238), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n250), .B1(new_n219), .B2(new_n215), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n221), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n251), .A2(new_n263), .A3(new_n264), .A4(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT83), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n255), .A2(new_n262), .B1(new_n221), .B2(new_n265), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n270), .A2(KEYINPUT83), .A3(new_n264), .A4(new_n251), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n249), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT86), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n245), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI211_X1 g088(.A(KEYINPUT86), .B(new_n249), .C1(new_n269), .C2(new_n271), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT87), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n269), .A2(new_n271), .ZN(new_n277));
  INV_X1    g091(.A(new_n249), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT86), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT87), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n272), .A2(new_n273), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n280), .A2(new_n281), .A3(new_n282), .A4(new_n245), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n251), .A2(new_n263), .A3(new_n266), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n240), .ZN(new_n285));
  XOR2_X1   g099(.A(new_n285), .B(KEYINPUT85), .Z(new_n286));
  INV_X1    g100(.A(new_n277), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n249), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n276), .A2(new_n283), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G469), .ZN(new_n290));
  INV_X1    g104(.A(G902), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n290), .A2(new_n291), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n278), .B1(new_n245), .B2(new_n277), .ZN(new_n294));
  XNOR2_X1  g108(.A(new_n285), .B(KEYINPUT85), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n294), .B1(new_n272), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n293), .B1(new_n296), .B2(G469), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n189), .B1(new_n292), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT88), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n298), .B(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G214), .B1(G237), .B2(G902), .ZN(new_n301));
  INV_X1    g115(.A(G952), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n302), .A2(G953), .ZN(new_n303));
  INV_X1    g117(.A(G234), .ZN(new_n304));
  INV_X1    g118(.A(G237), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  AOI211_X1 g121(.A(new_n291), .B(new_n246), .C1(G234), .C2(G237), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT21), .B(G898), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT6), .ZN(new_n312));
  INV_X1    g126(.A(G116), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(G119), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT69), .B(G116), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n314), .B1(new_n315), .B2(G119), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT2), .B(G113), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n313), .A2(KEYINPUT69), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT69), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G116), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(new_n322), .A3(G119), .ZN(new_n323));
  INV_X1    g137(.A(new_n314), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(new_n317), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n319), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n256), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n255), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n323), .A2(KEYINPUT5), .A3(new_n324), .ZN(new_n330));
  INV_X1    g144(.A(G113), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT5), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n331), .B1(new_n314), .B2(new_n332), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n330), .A2(new_n333), .B1(new_n316), .B2(new_n318), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(new_n221), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G110), .B(G122), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(KEYINPUT89), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n312), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n256), .B1(new_n326), .B2(new_n319), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n340), .A2(new_n255), .B1(new_n221), .B2(new_n334), .ZN(new_n341));
  AOI21_X1  g155(.A(KEYINPUT90), .B1(new_n341), .B2(new_n337), .ZN(new_n342));
  AND4_X1   g156(.A1(KEYINPUT90), .A2(new_n329), .A3(new_n337), .A4(new_n335), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n339), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT91), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT74), .B(G125), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n220), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n347), .B1(new_n261), .B2(new_n346), .ZN(new_n348));
  INV_X1    g162(.A(G224), .ZN(new_n349));
  OR2_X1    g163(.A1(new_n349), .A2(G953), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n348), .B(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n338), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n341), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n312), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n329), .A2(new_n337), .A3(new_n335), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT90), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n341), .A2(KEYINPUT90), .A3(new_n337), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT91), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(new_n339), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n345), .A2(new_n351), .A3(new_n354), .A4(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT92), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(KEYINPUT6), .B1(new_n341), .B2(new_n352), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(new_n357), .B2(new_n358), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n366), .A2(new_n360), .B1(new_n312), .B2(new_n353), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n367), .A2(KEYINPUT92), .A3(new_n351), .A4(new_n345), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n337), .B(KEYINPUT8), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n330), .A2(KEYINPUT93), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(new_n333), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n330), .A2(KEYINPUT93), .ZN(new_n373));
  OAI211_X1 g187(.A(new_n319), .B(new_n221), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT94), .ZN(new_n375));
  OAI22_X1  g189(.A1(new_n374), .A2(new_n375), .B1(new_n221), .B2(new_n334), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n374), .A2(new_n375), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n370), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n350), .A2(KEYINPUT7), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n348), .B(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n359), .A3(new_n380), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n381), .A2(KEYINPUT95), .A3(new_n291), .ZN(new_n382));
  AOI21_X1  g196(.A(KEYINPUT95), .B1(new_n381), .B2(new_n291), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(G210), .B1(G237), .B2(G902), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n369), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n385), .B1(new_n369), .B2(new_n384), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n301), .B(new_n311), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT20), .ZN(new_n389));
  NOR2_X1   g203(.A1(G475), .A2(G902), .ZN(new_n390));
  XNOR2_X1  g204(.A(G113), .B(G122), .ZN(new_n391));
  XNOR2_X1  g205(.A(KEYINPUT96), .B(G104), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n391), .B(new_n392), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n246), .A2(G143), .A3(G214), .A4(new_n305), .ZN(new_n394));
  OR2_X1    g208(.A1(KEYINPUT71), .A2(G953), .ZN(new_n395));
  NAND2_X1  g209(.A1(KEYINPUT71), .A2(G953), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n395), .A2(G214), .A3(new_n305), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n207), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(KEYINPUT18), .A3(G131), .ZN(new_n400));
  NOR2_X1   g214(.A1(G125), .A2(G140), .ZN(new_n401));
  XOR2_X1   g215(.A(KEYINPUT74), .B(G125), .Z(new_n402));
  AOI21_X1  g216(.A(new_n401), .B1(new_n402), .B2(G140), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G146), .ZN(new_n404));
  XOR2_X1   g218(.A(G125), .B(G140), .Z(new_n405));
  OR2_X1    g219(.A1(new_n405), .A2(G146), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(KEYINPUT18), .A2(G131), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n394), .A2(new_n398), .A3(new_n408), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n400), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT17), .ZN(new_n411));
  AOI211_X1 g225(.A(new_n411), .B(new_n228), .C1(new_n394), .C2(new_n398), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n394), .A2(new_n228), .A3(new_n398), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n228), .B1(new_n394), .B2(new_n398), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n412), .B1(new_n415), .B2(new_n411), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT16), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT74), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(G125), .ZN(new_n419));
  INV_X1    g233(.A(G125), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n420), .A2(KEYINPUT74), .ZN(new_n421));
  OAI21_X1  g235(.A(G140), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n401), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n417), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n346), .A2(KEYINPUT16), .A3(G140), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n205), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(G140), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n402), .A2(new_n417), .A3(new_n427), .ZN(new_n428));
  OAI211_X1 g242(.A(G146), .B(new_n428), .C1(new_n403), .C2(new_n417), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n429), .A3(KEYINPUT75), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT75), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n431), .B(new_n205), .C1(new_n424), .C2(new_n425), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  AOI211_X1 g247(.A(new_n393), .B(new_n410), .C1(new_n416), .C2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n393), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n405), .A2(KEYINPUT19), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(new_n403), .B2(KEYINPUT19), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  OAI221_X1 g252(.A(new_n429), .B1(new_n413), .B2(new_n414), .C1(new_n438), .C2(G146), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n400), .A2(new_n407), .A3(new_n409), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n435), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n389), .B(new_n390), .C1(new_n434), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT97), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n410), .B1(new_n416), .B2(new_n433), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n441), .B1(new_n435), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n390), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT20), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n435), .ZN(new_n448));
  INV_X1    g262(.A(new_n441), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT97), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n450), .A2(new_n451), .A3(new_n389), .A4(new_n390), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n443), .A2(new_n447), .A3(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n444), .A2(new_n435), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n291), .B1(new_n454), .B2(new_n434), .ZN(new_n455));
  XOR2_X1   g269(.A(KEYINPUT98), .B(G475), .Z(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AND2_X1   g271(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G217), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n187), .A2(new_n459), .A3(G953), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n315), .A2(G122), .ZN(new_n462));
  OR2_X1    g276(.A1(new_n313), .A2(G122), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n462), .A2(new_n194), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n218), .A2(G143), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT99), .B1(new_n212), .B2(G143), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT99), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(new_n207), .A3(G128), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n465), .A2(new_n229), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n229), .B1(new_n465), .B2(new_n469), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n315), .A2(KEYINPUT14), .A3(G122), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G107), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n462), .A2(new_n463), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT14), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(KEYINPUT101), .B1(new_n472), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n471), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n465), .A2(new_n229), .A3(new_n469), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n462), .A2(new_n463), .ZN(new_n482));
  OAI211_X1 g296(.A(G107), .B(new_n473), .C1(new_n482), .C2(KEYINPUT14), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT101), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n481), .A2(new_n483), .A3(new_n484), .A4(new_n464), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n478), .A2(new_n485), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n462), .A2(new_n194), .A3(new_n463), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n194), .B1(new_n462), .B2(new_n463), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT13), .ZN(new_n490));
  AOI22_X1  g304(.A1(new_n469), .A2(new_n490), .B1(new_n218), .B2(G143), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n466), .A2(new_n468), .A3(KEYINPUT13), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n229), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT100), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n489), .A2(new_n494), .A3(new_n495), .A4(new_n480), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n480), .B1(new_n487), .B2(new_n488), .ZN(new_n497));
  OAI21_X1  g311(.A(KEYINPUT100), .B1(new_n497), .B2(new_n493), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n461), .B1(new_n486), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n478), .A2(new_n485), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n501), .A2(new_n498), .A3(new_n496), .A4(new_n460), .ZN(new_n502));
  AOI21_X1  g316(.A(G902), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(G478), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(KEYINPUT15), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n503), .B(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n458), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n388), .A2(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n300), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n246), .A2(G221), .A3(G234), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT22), .B(G137), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n512), .B(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n218), .A2(KEYINPUT23), .A3(G119), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT23), .B1(new_n212), .B2(G119), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n212), .A2(G119), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n517), .B1(new_n218), .B2(G119), .ZN(new_n520));
  XOR2_X1   g334(.A(KEYINPUT24), .B(G110), .Z(new_n521));
  AOI22_X1  g335(.A1(new_n519), .A2(G110), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n430), .A2(new_n432), .A3(new_n522), .ZN(new_n523));
  OAI22_X1  g337(.A1(new_n519), .A2(G110), .B1(new_n520), .B2(new_n521), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(new_n429), .A3(new_n406), .ZN(new_n525));
  AND3_X1   g339(.A1(new_n523), .A2(KEYINPUT78), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(KEYINPUT78), .B1(new_n523), .B2(new_n525), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n514), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n514), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n523), .A2(new_n525), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT78), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n528), .A2(new_n291), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT25), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT25), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n528), .A2(new_n535), .A3(new_n532), .A4(new_n291), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n459), .B1(G234), .B2(new_n291), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n537), .B(KEYINPUT73), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n534), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT79), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT79), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n534), .A2(new_n541), .A3(new_n536), .A4(new_n538), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n537), .A2(G902), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n528), .A2(new_n532), .A3(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(KEYINPUT80), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n540), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT81), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n540), .A2(KEYINPUT81), .A3(new_n542), .A4(new_n545), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(G472), .ZN(new_n551));
  INV_X1    g365(.A(new_n261), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n240), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n327), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT67), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(new_n224), .B2(G134), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n225), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n230), .A2(new_n555), .ZN(new_n558));
  OAI21_X1  g372(.A(G131), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n206), .A2(KEYINPUT1), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n212), .A2(KEYINPUT68), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT68), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(G128), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n214), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  AND4_X1   g379(.A1(new_n210), .A2(new_n206), .A3(new_n208), .A4(G128), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n559), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(new_n237), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n553), .A2(new_n554), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT28), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n240), .A2(new_n552), .B1(new_n237), .B2(new_n568), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(KEYINPUT28), .A3(new_n554), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n567), .B1(new_n236), .B2(new_n233), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n240), .A2(KEYINPUT66), .A3(new_n552), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT66), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n264), .B2(new_n261), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n575), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n572), .B(new_n574), .C1(new_n554), .C2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n246), .A2(G210), .A3(new_n305), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(KEYINPUT27), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT26), .B(G101), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n580), .A2(new_n585), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(KEYINPUT29), .ZN(new_n587));
  INV_X1    g401(.A(new_n570), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT70), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n589), .B1(new_n573), .B2(KEYINPUT30), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n261), .B1(new_n237), .B2(new_n239), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT30), .ZN(new_n592));
  NOR4_X1   g406(.A1(new_n591), .A2(new_n575), .A3(KEYINPUT70), .A4(new_n592), .ZN(new_n593));
  OAI22_X1  g407(.A1(new_n590), .A2(new_n593), .B1(new_n579), .B2(KEYINPUT30), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n588), .B1(new_n595), .B2(new_n327), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n587), .B1(new_n584), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n327), .B1(new_n591), .B2(new_n575), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n570), .A2(KEYINPUT72), .A3(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT72), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n600), .B(new_n327), .C1(new_n591), .C2(new_n575), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(KEYINPUT28), .A3(new_n601), .ZN(new_n602));
  AND4_X1   g416(.A1(KEYINPUT29), .A2(new_n602), .A3(new_n584), .A4(new_n572), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(G902), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n551), .B1(new_n597), .B2(new_n604), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n584), .B(new_n570), .C1(new_n594), .C2(new_n554), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(KEYINPUT31), .ZN(new_n607));
  OAI221_X1 g421(.A(new_n327), .B1(new_n579), .B2(KEYINPUT30), .C1(new_n590), .C2(new_n593), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT31), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n608), .A2(new_n609), .A3(new_n584), .A4(new_n570), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n580), .A2(new_n585), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n607), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(G472), .A2(G902), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT32), .ZN(new_n615));
  INV_X1    g429(.A(new_n613), .ZN(new_n616));
  AOI22_X1  g430(.A1(new_n606), .A2(KEYINPUT31), .B1(new_n585), .B2(new_n580), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n616), .B1(new_n617), .B2(new_n610), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT32), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n605), .B1(new_n615), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n550), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n509), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G101), .ZN(G3));
  INV_X1    g438(.A(new_n550), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n551), .B1(new_n612), .B2(new_n291), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(new_n618), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n300), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT33), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n500), .A2(new_n629), .A3(new_n502), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n629), .B1(new_n500), .B2(new_n502), .ZN(new_n631));
  OAI211_X1 g445(.A(G478), .B(new_n291), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n500), .A2(new_n502), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n291), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n633), .B1(new_n635), .B2(new_n504), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n503), .A2(KEYINPUT102), .A3(G478), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n632), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n458), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n388), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n628), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(new_n190), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT103), .B(KEYINPUT34), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G6));
  INV_X1    g460(.A(new_n457), .ZN(new_n647));
  INV_X1    g461(.A(new_n506), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n447), .A2(KEYINPUT104), .A3(new_n442), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n447), .A2(new_n442), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT104), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n648), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n388), .A2(new_n647), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n628), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT105), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT35), .B(G107), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G9));
  INV_X1    g472(.A(new_n627), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n529), .A2(KEYINPUT36), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(new_n530), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(new_n543), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n540), .A2(new_n542), .A3(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n509), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT37), .B(G110), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(G12));
  INV_X1    g481(.A(new_n301), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n369), .A2(new_n384), .ZN(new_n669));
  INV_X1    g483(.A(new_n385), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n369), .A2(new_n385), .A3(new_n384), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n668), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n540), .A2(new_n542), .A3(new_n662), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT106), .B(G900), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n307), .B1(new_n308), .B2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n457), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n653), .A2(new_n678), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n673), .A2(new_n674), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n597), .A2(new_n604), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(G472), .ZN(new_n682));
  AOI211_X1 g496(.A(KEYINPUT32), .B(new_n616), .C1(new_n617), .C2(new_n610), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n619), .B1(new_n612), .B2(new_n613), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n682), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n680), .A2(new_n300), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  XOR2_X1   g501(.A(new_n676), .B(KEYINPUT39), .Z(new_n688));
  NAND2_X1  g502(.A1(new_n300), .A2(new_n688), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n689), .A2(KEYINPUT40), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n671), .A2(new_n672), .ZN(new_n691));
  XNOR2_X1  g505(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n691), .B(new_n692), .Z(new_n693));
  NOR3_X1   g507(.A1(new_n693), .A2(new_n668), .A3(new_n674), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n689), .A2(KEYINPUT40), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n458), .A2(new_n506), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n615), .A2(new_n620), .ZN(new_n698));
  INV_X1    g512(.A(new_n606), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n599), .A2(new_n601), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n699), .B1(new_n585), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g515(.A(G472), .B1(new_n701), .B2(G902), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n697), .B1(new_n698), .B2(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n690), .A2(new_n694), .A3(new_n695), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G143), .ZN(G45));
  OAI211_X1 g519(.A(new_n301), .B(new_n677), .C1(new_n386), .C2(new_n387), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n640), .A2(new_n674), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n300), .A2(new_n685), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G146), .ZN(G48));
  AND3_X1   g524(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n290), .B1(new_n289), .B2(new_n291), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n711), .A2(new_n712), .A3(new_n189), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n622), .A2(new_n642), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  NAND3_X1  g530(.A1(new_n654), .A2(new_n622), .A3(new_n713), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G116), .ZN(G18));
  INV_X1    g532(.A(new_n507), .ZN(new_n719));
  AND4_X1   g533(.A1(new_n685), .A2(new_n311), .A3(new_n719), .A4(new_n674), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n301), .B1(new_n386), .B2(new_n387), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n289), .A2(new_n291), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(G469), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n188), .A3(new_n292), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n721), .A2(new_n724), .A3(KEYINPUT108), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n726), .B1(new_n673), .B2(new_n713), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n720), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G119), .ZN(G21));
  NAND2_X1  g543(.A1(new_n602), .A2(new_n572), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n584), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n602), .A2(KEYINPUT109), .A3(new_n572), .ZN(new_n733));
  AOI22_X1  g547(.A1(new_n732), .A2(new_n733), .B1(KEYINPUT31), .B2(new_n606), .ZN(new_n734));
  AOI22_X1  g548(.A1(new_n734), .A2(KEYINPUT110), .B1(new_n609), .B2(new_n699), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n732), .A2(new_n733), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n607), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n616), .B1(new_n735), .B2(new_n739), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n740), .A2(new_n546), .A3(new_n626), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n724), .A2(new_n310), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n741), .A2(new_n673), .A3(new_n696), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  OAI21_X1  g558(.A(KEYINPUT108), .B1(new_n721), .B2(new_n724), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n673), .A2(new_n713), .A3(new_n726), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n453), .A2(new_n457), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n638), .A3(new_n677), .ZN(new_n749));
  NOR4_X1   g563(.A1(new_n740), .A2(new_n626), .A3(new_n663), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G125), .ZN(G27));
  INV_X1    g566(.A(KEYINPUT42), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n754), .B1(new_n621), .B2(new_n546), .ZN(new_n755));
  INV_X1    g569(.A(new_n546), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n685), .A2(KEYINPUT113), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n242), .A2(new_n244), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n759), .B(new_n249), .C1(new_n287), .C2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n295), .A2(new_n272), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n294), .A2(new_n759), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n293), .B1(new_n765), .B2(G469), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n189), .B1(new_n766), .B2(new_n292), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI211_X1 g583(.A(KEYINPUT112), .B(new_n189), .C1(new_n766), .C2(new_n292), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n748), .A2(new_n638), .A3(new_n677), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(new_n671), .A3(new_n301), .A4(new_n672), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n769), .A2(new_n770), .A3(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n753), .B1(new_n758), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n766), .A2(new_n292), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n188), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT112), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n671), .A2(new_n301), .A3(new_n672), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n767), .A2(new_n768), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n778), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n685), .A2(new_n548), .A3(new_n549), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n771), .A2(new_n753), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n775), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(new_n228), .ZN(G33));
  NOR2_X1   g602(.A1(new_n769), .A2(new_n770), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n789), .A2(new_n622), .A3(new_n679), .A4(new_n780), .ZN(new_n790));
  XOR2_X1   g604(.A(KEYINPUT114), .B(G134), .Z(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(G36));
  NOR3_X1   g606(.A1(new_n639), .A2(KEYINPUT43), .A3(new_n748), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n748), .A2(KEYINPUT117), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n748), .A2(KEYINPUT117), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n795), .A2(new_n796), .A3(new_n639), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT43), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n794), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT44), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n659), .A2(new_n674), .ZN(new_n801));
  OR3_X1    g615(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n800), .B1(new_n799), .B2(new_n801), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n803), .A3(new_n780), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(G469), .B1(new_n296), .B2(KEYINPUT45), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n807), .B1(KEYINPUT45), .B2(new_n765), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n293), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT115), .B1(new_n809), .B2(KEYINPUT46), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n711), .B1(new_n809), .B2(KEYINPUT46), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT46), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n812), .B(new_n813), .C1(new_n808), .C2(new_n293), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n810), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n815), .A2(new_n188), .A3(new_n688), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT116), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT116), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n815), .A2(new_n818), .A3(new_n188), .A4(new_n688), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n802), .A2(new_n803), .A3(KEYINPUT118), .A4(new_n780), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n806), .A2(new_n820), .A3(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G137), .ZN(G39));
  NAND2_X1  g637(.A1(new_n815), .A2(new_n188), .ZN(new_n824));
  AND2_X1   g638(.A1(KEYINPUT119), .A2(KEYINPUT47), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(KEYINPUT119), .A2(KEYINPUT47), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n828), .B1(new_n815), .B2(new_n188), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n780), .A2(new_n550), .A3(new_n621), .A4(new_n771), .ZN(new_n830));
  OR3_X1    g644(.A1(new_n826), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(G140), .ZN(G42));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n750), .A2(new_n789), .A3(new_n780), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n790), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n298), .A2(new_n299), .ZN(new_n836));
  AOI211_X1 g650(.A(KEYINPUT88), .B(new_n189), .C1(new_n292), .C2(new_n297), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n685), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n648), .A2(new_n678), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n674), .A2(new_n649), .A3(new_n652), .A4(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n779), .ZN(new_n841));
  INV_X1    g655(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(KEYINPUT120), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n300), .A2(new_n844), .A3(new_n685), .A4(new_n841), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n835), .A2(new_n775), .A3(new_n786), .A4(new_n846), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n717), .A2(new_n743), .A3(new_n714), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n507), .B1(new_n458), .B2(new_n638), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n388), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n300), .A2(new_n625), .A3(new_n627), .A4(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n728), .A2(new_n851), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n300), .B(new_n508), .C1(new_n622), .C2(new_n664), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n848), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n706), .A2(new_n777), .A3(new_n674), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n747), .A2(new_n750), .B1(new_n703), .B2(new_n856), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n685), .B(new_n300), .C1(new_n680), .C2(new_n708), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT52), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n857), .A2(new_n858), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n857), .A2(KEYINPUT52), .A3(new_n858), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(KEYINPUT121), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n855), .A2(new_n861), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n790), .A2(new_n834), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n870), .A2(new_n774), .A3(new_n785), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n853), .A2(new_n728), .A3(new_n851), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n717), .A2(new_n743), .A3(new_n714), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n871), .A2(new_n874), .A3(new_n846), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n856), .A2(new_n703), .ZN(new_n876));
  AND4_X1   g690(.A1(KEYINPUT52), .A2(new_n858), .A3(new_n751), .A4(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(new_n859), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n875), .A2(new_n878), .A3(new_n868), .ZN(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n833), .B1(new_n869), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT51), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n711), .A2(new_n712), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n189), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n884), .B1(new_n826), .B2(new_n829), .ZN(new_n885));
  INV_X1    g699(.A(new_n799), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n886), .A2(new_n307), .A3(new_n741), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n780), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n693), .A2(new_n668), .A3(new_n713), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(new_n887), .ZN(new_n891));
  XOR2_X1   g705(.A(KEYINPUT122), .B(KEYINPUT50), .Z(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(KEYINPUT122), .A2(KEYINPUT50), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n890), .A2(new_n887), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n780), .A2(new_n713), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n799), .A2(new_n896), .A3(new_n306), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n740), .A2(new_n626), .A3(new_n663), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n896), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n698), .A2(new_n702), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n900), .A2(new_n625), .A3(new_n307), .A4(new_n901), .ZN(new_n902));
  OR3_X1    g716(.A1(new_n902), .A2(new_n748), .A3(new_n638), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n893), .A2(new_n895), .A3(new_n899), .A4(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n882), .B1(new_n889), .B2(new_n904), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n893), .A2(new_n899), .A3(new_n903), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n906), .A2(new_n888), .A3(KEYINPUT51), .A4(new_n895), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n897), .A2(new_n758), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT123), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n909), .A3(KEYINPUT48), .ZN(new_n910));
  XOR2_X1   g724(.A(KEYINPUT123), .B(KEYINPUT48), .Z(new_n911));
  OAI21_X1  g725(.A(new_n910), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n887), .A2(new_n747), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n913), .B(new_n303), .C1(new_n641), .C2(new_n902), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n905), .A2(new_n907), .A3(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n855), .A2(KEYINPUT53), .A3(new_n861), .A4(new_n866), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n868), .B1(new_n875), .B2(new_n878), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n917), .A2(new_n833), .A3(new_n918), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n881), .A2(new_n916), .A3(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(G952), .A2(G953), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n797), .A2(new_n756), .A3(new_n188), .A4(new_n301), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n883), .B(KEYINPUT49), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n693), .A2(new_n923), .A3(new_n901), .ZN(new_n924));
  OAI22_X1  g738(.A1(new_n920), .A2(new_n921), .B1(new_n922), .B2(new_n924), .ZN(G75));
  NAND2_X1  g739(.A1(new_n917), .A2(new_n918), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n926), .A2(G210), .A3(G902), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT56), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n367), .A2(new_n345), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(new_n351), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT55), .Z(new_n931));
  AND3_X1   g745(.A1(new_n927), .A2(new_n928), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n931), .B1(new_n927), .B2(new_n928), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n246), .A2(G952), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(G51));
  XNOR2_X1  g749(.A(new_n293), .B(KEYINPUT57), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n833), .B1(new_n917), .B2(new_n918), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n936), .B1(new_n919), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n289), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n926), .A2(G902), .A3(new_n808), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n934), .B1(new_n939), .B2(new_n940), .ZN(G54));
  INV_X1    g755(.A(new_n934), .ZN(new_n942));
  NAND2_X1  g756(.A1(KEYINPUT58), .A2(G475), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n926), .A2(G902), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n942), .B1(new_n945), .B2(new_n445), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n445), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(KEYINPUT124), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT124), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n945), .A2(new_n949), .A3(new_n445), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n946), .B1(new_n948), .B2(new_n950), .ZN(G60));
  OR2_X1    g765(.A1(new_n630), .A2(new_n631), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n917), .A2(new_n833), .A3(new_n918), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n879), .B1(new_n868), .B2(new_n867), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n953), .B1(new_n954), .B2(new_n833), .ZN(new_n955));
  NAND2_X1  g769(.A1(G478), .A2(G902), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT59), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n952), .B1(new_n955), .B2(new_n957), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n952), .A2(new_n957), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n919), .B2(new_n937), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n942), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n958), .A2(new_n961), .ZN(G63));
  XNOR2_X1  g776(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  XNOR2_X1  g778(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n459), .A2(new_n291), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n917), .B2(new_n918), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n661), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n528), .A2(new_n532), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n942), .B1(new_n969), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n964), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n926), .A2(new_n967), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n972), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n977), .A2(new_n942), .A3(new_n970), .A4(new_n963), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n975), .A2(new_n978), .ZN(G66));
  OAI21_X1  g793(.A(G953), .B1(new_n309), .B2(new_n349), .ZN(new_n980));
  INV_X1    g794(.A(new_n246), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n980), .B1(new_n874), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(G898), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n929), .B1(new_n983), .B2(new_n981), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n982), .B(new_n984), .Z(G69));
  XNOR2_X1  g799(.A(new_n594), .B(new_n438), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n981), .A2(G900), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n822), .A2(new_n831), .ZN(new_n989));
  AOI211_X1 g803(.A(new_n721), .B(new_n697), .C1(new_n755), .C2(new_n757), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n820), .A2(new_n990), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n858), .A2(new_n751), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n775), .A2(new_n786), .A3(new_n790), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n991), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n989), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n988), .B1(new_n995), .B2(new_n246), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n246), .B1(G227), .B2(G900), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  NOR4_X1   g813(.A1(new_n689), .A2(new_n783), .A3(new_n779), .A4(new_n849), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n704), .A2(new_n992), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT62), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n704), .A2(KEYINPUT62), .A3(new_n992), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1000), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n989), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n981), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n997), .B(new_n999), .C1(new_n1007), .C2(new_n986), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1007), .A2(new_n986), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n998), .B1(new_n1009), .B2(new_n996), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1008), .A2(new_n1010), .ZN(G72));
  NAND2_X1  g825(.A1(G472), .A2(G902), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(KEYINPUT63), .Z(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1014), .B1(new_n995), .B2(new_n874), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n596), .B(KEYINPUT127), .ZN(new_n1016));
  OR2_X1    g830(.A1(new_n1016), .A2(new_n584), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n942), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g832(.A1(new_n596), .A2(new_n584), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1013), .B1(new_n1019), .B2(new_n699), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n954), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1016), .A2(new_n584), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1005), .A2(new_n1006), .A3(new_n874), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1022), .B1(new_n1023), .B2(new_n1013), .ZN(new_n1024));
  NOR3_X1   g838(.A1(new_n1018), .A2(new_n1021), .A3(new_n1024), .ZN(G57));
endmodule


