

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U545 ( .A1(n717), .A2(n716), .ZN(n718) );
  OR2_X1 U546 ( .A1(n734), .A2(n511), .ZN(n735) );
  NOR2_X2 U547 ( .A1(n526), .A2(n525), .ZN(G160) );
  BUF_X1 U548 ( .A(n544), .Z(n545) );
  NAND2_X1 U549 ( .A1(n513), .A2(n512), .ZN(n795) );
  XNOR2_X1 U550 ( .A(n519), .B(KEYINPUT23), .ZN(n520) );
  AND2_X1 U551 ( .A1(n510), .A2(n794), .ZN(n509) );
  AND2_X1 U552 ( .A1(n803), .A2(n793), .ZN(n510) );
  AND2_X1 U553 ( .A1(G8), .A2(n733), .ZN(n511) );
  OR2_X1 U554 ( .A1(n759), .A2(n758), .ZN(n512) );
  AND2_X1 U555 ( .A1(n756), .A2(n755), .ZN(n513) );
  INV_X1 U556 ( .A(KEYINPUT93), .ZN(n707) );
  AND2_X1 U557 ( .A1(n772), .A2(n670), .ZN(n686) );
  NOR2_X1 U558 ( .A1(n706), .A2(n705), .ZN(n717) );
  XNOR2_X1 U559 ( .A(n718), .B(KEYINPUT94), .ZN(n731) );
  NAND2_X1 U560 ( .A1(G8), .A2(n720), .ZN(n759) );
  INV_X1 U561 ( .A(KEYINPUT64), .ZN(n519) );
  XOR2_X1 U562 ( .A(KEYINPUT15), .B(n579), .Z(n925) );
  XNOR2_X1 U563 ( .A(KEYINPUT67), .B(n531), .ZN(n631) );
  NOR2_X1 U564 ( .A1(G2104), .A2(n522), .ZN(n879) );
  XNOR2_X1 U565 ( .A(n521), .B(n520), .ZN(n524) );
  XNOR2_X1 U566 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n515) );
  NOR2_X1 U567 ( .A1(G2105), .A2(G2104), .ZN(n514) );
  XNOR2_X1 U568 ( .A(n515), .B(n514), .ZN(n544) );
  NAND2_X1 U569 ( .A1(n544), .A2(G137), .ZN(n517) );
  AND2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n876) );
  NAND2_X1 U571 ( .A1(G113), .A2(n876), .ZN(n516) );
  NAND2_X1 U572 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U573 ( .A(n518), .B(KEYINPUT66), .ZN(n526) );
  INV_X1 U574 ( .A(G2105), .ZN(n522) );
  AND2_X1 U575 ( .A1(n522), .A2(G2104), .ZN(n663) );
  NAND2_X1 U576 ( .A1(G101), .A2(n663), .ZN(n521) );
  NAND2_X1 U577 ( .A1(G125), .A2(n879), .ZN(n523) );
  NAND2_X1 U578 ( .A1(n524), .A2(n523), .ZN(n525) );
  NOR2_X1 U579 ( .A1(G651), .A2(G543), .ZN(n626) );
  NAND2_X1 U580 ( .A1(G91), .A2(n626), .ZN(n529) );
  INV_X1 U581 ( .A(G651), .ZN(n530) );
  NOR2_X1 U582 ( .A1(G543), .A2(n530), .ZN(n527) );
  XOR2_X1 U583 ( .A(KEYINPUT1), .B(n527), .Z(n627) );
  NAND2_X1 U584 ( .A1(G65), .A2(n627), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n529), .A2(n528), .ZN(n536) );
  XOR2_X1 U586 ( .A(G543), .B(KEYINPUT0), .Z(n532) );
  OR2_X1 U587 ( .A1(n530), .A2(n532), .ZN(n531) );
  NAND2_X1 U588 ( .A1(G78), .A2(n631), .ZN(n534) );
  NOR2_X2 U589 ( .A1(G651), .A2(n532), .ZN(n635) );
  NAND2_X1 U590 ( .A1(G53), .A2(n635), .ZN(n533) );
  NAND2_X1 U591 ( .A1(n534), .A2(n533), .ZN(n535) );
  OR2_X1 U592 ( .A1(n536), .A2(n535), .ZN(G299) );
  NAND2_X1 U593 ( .A1(G85), .A2(n626), .ZN(n538) );
  NAND2_X1 U594 ( .A1(G60), .A2(n627), .ZN(n537) );
  NAND2_X1 U595 ( .A1(n538), .A2(n537), .ZN(n542) );
  NAND2_X1 U596 ( .A1(G72), .A2(n631), .ZN(n540) );
  NAND2_X1 U597 ( .A1(G47), .A2(n635), .ZN(n539) );
  NAND2_X1 U598 ( .A1(n540), .A2(n539), .ZN(n541) );
  OR2_X1 U599 ( .A1(n542), .A2(n541), .ZN(G290) );
  AND2_X1 U600 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U601 ( .A1(n879), .A2(G123), .ZN(n543) );
  XNOR2_X1 U602 ( .A(n543), .B(KEYINPUT18), .ZN(n547) );
  NAND2_X1 U603 ( .A1(G135), .A2(n545), .ZN(n546) );
  NAND2_X1 U604 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U605 ( .A(KEYINPUT71), .B(n548), .ZN(n552) );
  NAND2_X1 U606 ( .A1(n663), .A2(G99), .ZN(n550) );
  NAND2_X1 U607 ( .A1(G111), .A2(n876), .ZN(n549) );
  AND2_X1 U608 ( .A1(n550), .A2(n549), .ZN(n551) );
  NAND2_X1 U609 ( .A1(n552), .A2(n551), .ZN(n990) );
  XNOR2_X1 U610 ( .A(G2096), .B(n990), .ZN(n553) );
  OR2_X1 U611 ( .A1(G2100), .A2(n553), .ZN(G156) );
  NAND2_X1 U612 ( .A1(G52), .A2(n635), .ZN(n555) );
  NAND2_X1 U613 ( .A1(G64), .A2(n627), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n560) );
  NAND2_X1 U615 ( .A1(G90), .A2(n626), .ZN(n557) );
  NAND2_X1 U616 ( .A1(G77), .A2(n631), .ZN(n556) );
  NAND2_X1 U617 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U618 ( .A(KEYINPUT9), .B(n558), .Z(n559) );
  NOR2_X1 U619 ( .A1(n560), .A2(n559), .ZN(G171) );
  NAND2_X1 U620 ( .A1(G7), .A2(G661), .ZN(n561) );
  XNOR2_X1 U621 ( .A(n561), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U622 ( .A(G223), .ZN(n822) );
  NAND2_X1 U623 ( .A1(n822), .A2(G567), .ZN(n562) );
  XOR2_X1 U624 ( .A(KEYINPUT11), .B(n562), .Z(G234) );
  NAND2_X1 U625 ( .A1(n626), .A2(G81), .ZN(n563) );
  XNOR2_X1 U626 ( .A(n563), .B(KEYINPUT12), .ZN(n565) );
  NAND2_X1 U627 ( .A1(G68), .A2(n631), .ZN(n564) );
  NAND2_X1 U628 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U629 ( .A(n566), .B(KEYINPUT13), .ZN(n568) );
  NAND2_X1 U630 ( .A1(G43), .A2(n635), .ZN(n567) );
  NAND2_X1 U631 ( .A1(n568), .A2(n567), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n627), .A2(G56), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT14), .B(n569), .Z(n570) );
  NOR2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n684) );
  BUF_X1 U635 ( .A(n684), .Z(n915) );
  NAND2_X1 U636 ( .A1(n915), .A2(G860), .ZN(G153) );
  INV_X1 U637 ( .A(G171), .ZN(G301) );
  INV_X1 U638 ( .A(G868), .ZN(n647) );
  NOR2_X1 U639 ( .A1(G301), .A2(n647), .ZN(n581) );
  NAND2_X1 U640 ( .A1(n631), .A2(G79), .ZN(n578) );
  NAND2_X1 U641 ( .A1(G92), .A2(n626), .ZN(n573) );
  NAND2_X1 U642 ( .A1(G66), .A2(n627), .ZN(n572) );
  NAND2_X1 U643 ( .A1(n573), .A2(n572), .ZN(n576) );
  NAND2_X1 U644 ( .A1(G54), .A2(n635), .ZN(n574) );
  XNOR2_X1 U645 ( .A(KEYINPUT69), .B(n574), .ZN(n575) );
  NOR2_X1 U646 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U647 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U648 ( .A1(G868), .A2(n925), .ZN(n580) );
  NOR2_X1 U649 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U650 ( .A(KEYINPUT70), .B(n582), .ZN(G284) );
  NAND2_X1 U651 ( .A1(n626), .A2(G89), .ZN(n583) );
  XNOR2_X1 U652 ( .A(n583), .B(KEYINPUT4), .ZN(n585) );
  NAND2_X1 U653 ( .A1(G76), .A2(n631), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U655 ( .A(n586), .B(KEYINPUT5), .ZN(n591) );
  NAND2_X1 U656 ( .A1(G51), .A2(n635), .ZN(n588) );
  NAND2_X1 U657 ( .A1(G63), .A2(n627), .ZN(n587) );
  NAND2_X1 U658 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U659 ( .A(KEYINPUT6), .B(n589), .Z(n590) );
  NAND2_X1 U660 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U661 ( .A(n592), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U662 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U663 ( .A1(G286), .A2(n647), .ZN(n594) );
  NOR2_X1 U664 ( .A1(G868), .A2(G299), .ZN(n593) );
  NOR2_X1 U665 ( .A1(n594), .A2(n593), .ZN(G297) );
  INV_X1 U666 ( .A(G860), .ZN(n595) );
  NAND2_X1 U667 ( .A1(n595), .A2(G559), .ZN(n596) );
  INV_X1 U668 ( .A(n925), .ZN(n601) );
  NAND2_X1 U669 ( .A1(n596), .A2(n601), .ZN(n597) );
  XNOR2_X1 U670 ( .A(n597), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U671 ( .A1(n601), .A2(G868), .ZN(n598) );
  NOR2_X1 U672 ( .A1(G559), .A2(n598), .ZN(n600) );
  AND2_X1 U673 ( .A1(n647), .A2(n915), .ZN(n599) );
  NOR2_X1 U674 ( .A1(n600), .A2(n599), .ZN(G282) );
  XOR2_X1 U675 ( .A(n915), .B(KEYINPUT72), .Z(n603) );
  NAND2_X1 U676 ( .A1(G559), .A2(n601), .ZN(n602) );
  XNOR2_X1 U677 ( .A(n603), .B(n602), .ZN(n644) );
  XOR2_X1 U678 ( .A(n644), .B(KEYINPUT73), .Z(n604) );
  NOR2_X1 U679 ( .A1(G860), .A2(n604), .ZN(n613) );
  NAND2_X1 U680 ( .A1(G80), .A2(n631), .ZN(n605) );
  XNOR2_X1 U681 ( .A(n605), .B(KEYINPUT74), .ZN(n612) );
  NAND2_X1 U682 ( .A1(G93), .A2(n626), .ZN(n607) );
  NAND2_X1 U683 ( .A1(G67), .A2(n627), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U685 ( .A1(G55), .A2(n635), .ZN(n608) );
  XNOR2_X1 U686 ( .A(KEYINPUT75), .B(n608), .ZN(n609) );
  NOR2_X1 U687 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n612), .A2(n611), .ZN(n646) );
  XOR2_X1 U689 ( .A(n613), .B(n646), .Z(G145) );
  NAND2_X1 U690 ( .A1(G49), .A2(n635), .ZN(n615) );
  NAND2_X1 U691 ( .A1(G74), .A2(G651), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U693 ( .A1(n627), .A2(n616), .ZN(n618) );
  NAND2_X1 U694 ( .A1(n532), .A2(G87), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n618), .A2(n617), .ZN(G288) );
  NAND2_X1 U696 ( .A1(n631), .A2(G75), .ZN(n621) );
  NAND2_X1 U697 ( .A1(n626), .A2(G88), .ZN(n619) );
  XOR2_X1 U698 ( .A(KEYINPUT77), .B(n619), .Z(n620) );
  NAND2_X1 U699 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G50), .A2(n635), .ZN(n623) );
  NAND2_X1 U701 ( .A1(G62), .A2(n627), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U703 ( .A1(n625), .A2(n624), .ZN(G166) );
  NAND2_X1 U704 ( .A1(G86), .A2(n626), .ZN(n629) );
  NAND2_X1 U705 ( .A1(G61), .A2(n627), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U707 ( .A(KEYINPUT76), .B(n630), .ZN(n634) );
  NAND2_X1 U708 ( .A1(n631), .A2(G73), .ZN(n632) );
  XOR2_X1 U709 ( .A(KEYINPUT2), .B(n632), .Z(n633) );
  NOR2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U711 ( .A1(n635), .A2(G48), .ZN(n636) );
  NAND2_X1 U712 ( .A1(n637), .A2(n636), .ZN(G305) );
  XNOR2_X1 U713 ( .A(KEYINPUT19), .B(G299), .ZN(n638) );
  XNOR2_X1 U714 ( .A(n638), .B(G288), .ZN(n641) );
  XNOR2_X1 U715 ( .A(G166), .B(G305), .ZN(n639) );
  XNOR2_X1 U716 ( .A(n639), .B(G290), .ZN(n640) );
  XNOR2_X1 U717 ( .A(n641), .B(n640), .ZN(n643) );
  XNOR2_X1 U718 ( .A(n646), .B(KEYINPUT78), .ZN(n642) );
  XNOR2_X1 U719 ( .A(n643), .B(n642), .ZN(n892) );
  XNOR2_X1 U720 ( .A(n892), .B(n644), .ZN(n645) );
  NAND2_X1 U721 ( .A1(n645), .A2(G868), .ZN(n649) );
  NAND2_X1 U722 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U723 ( .A1(n649), .A2(n648), .ZN(G295) );
  NAND2_X1 U724 ( .A1(G2084), .A2(G2078), .ZN(n650) );
  XOR2_X1 U725 ( .A(KEYINPUT20), .B(n650), .Z(n651) );
  NAND2_X1 U726 ( .A1(G2090), .A2(n651), .ZN(n652) );
  XNOR2_X1 U727 ( .A(KEYINPUT21), .B(n652), .ZN(n653) );
  NAND2_X1 U728 ( .A1(n653), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U729 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U730 ( .A(KEYINPUT68), .B(G57), .Z(G237) );
  XOR2_X1 U731 ( .A(KEYINPUT22), .B(KEYINPUT79), .Z(n655) );
  NAND2_X1 U732 ( .A1(G132), .A2(G82), .ZN(n654) );
  XNOR2_X1 U733 ( .A(n655), .B(n654), .ZN(n656) );
  NOR2_X1 U734 ( .A1(n656), .A2(G218), .ZN(n657) );
  NAND2_X1 U735 ( .A1(G96), .A2(n657), .ZN(n828) );
  NAND2_X1 U736 ( .A1(n828), .A2(G2106), .ZN(n661) );
  NAND2_X1 U737 ( .A1(G108), .A2(G120), .ZN(n658) );
  NOR2_X1 U738 ( .A1(G237), .A2(n658), .ZN(n659) );
  NAND2_X1 U739 ( .A1(G69), .A2(n659), .ZN(n829) );
  NAND2_X1 U740 ( .A1(G567), .A2(n829), .ZN(n660) );
  NAND2_X1 U741 ( .A1(n661), .A2(n660), .ZN(n831) );
  NAND2_X1 U742 ( .A1(G661), .A2(G483), .ZN(n662) );
  NOR2_X1 U743 ( .A1(n831), .A2(n662), .ZN(n825) );
  NAND2_X1 U744 ( .A1(n825), .A2(G36), .ZN(G176) );
  NAND2_X1 U745 ( .A1(G102), .A2(n663), .ZN(n665) );
  NAND2_X1 U746 ( .A1(G138), .A2(n545), .ZN(n664) );
  NAND2_X1 U747 ( .A1(n665), .A2(n664), .ZN(n669) );
  NAND2_X1 U748 ( .A1(G114), .A2(n876), .ZN(n667) );
  NAND2_X1 U749 ( .A1(G126), .A2(n879), .ZN(n666) );
  NAND2_X1 U750 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U751 ( .A1(n669), .A2(n668), .ZN(G164) );
  XOR2_X1 U752 ( .A(KEYINPUT80), .B(G166), .Z(G303) );
  NOR2_X1 U753 ( .A1(G164), .A2(G1384), .ZN(n772) );
  NAND2_X1 U754 ( .A1(G160), .A2(G40), .ZN(n771) );
  XOR2_X1 U755 ( .A(KEYINPUT88), .B(n771), .Z(n670) );
  NOR2_X1 U756 ( .A1(n686), .A2(G1961), .ZN(n672) );
  XOR2_X1 U757 ( .A(G2078), .B(KEYINPUT25), .Z(n964) );
  NAND2_X1 U758 ( .A1(n772), .A2(n670), .ZN(n720) );
  NOR2_X1 U759 ( .A1(n964), .A2(n720), .ZN(n671) );
  NOR2_X1 U760 ( .A1(n672), .A2(n671), .ZN(n712) );
  NOR2_X1 U761 ( .A1(n712), .A2(G301), .ZN(n673) );
  XOR2_X1 U762 ( .A(KEYINPUT89), .B(n673), .Z(n706) );
  NAND2_X1 U763 ( .A1(n686), .A2(G2072), .ZN(n675) );
  INV_X1 U764 ( .A(KEYINPUT27), .ZN(n674) );
  XNOR2_X1 U765 ( .A(n675), .B(n674), .ZN(n677) );
  NAND2_X1 U766 ( .A1(G1956), .A2(n720), .ZN(n676) );
  NAND2_X1 U767 ( .A1(n677), .A2(n676), .ZN(n698) );
  NOR2_X1 U768 ( .A1(n698), .A2(G299), .ZN(n681) );
  NAND2_X1 U769 ( .A1(G1348), .A2(n720), .ZN(n679) );
  NAND2_X1 U770 ( .A1(n686), .A2(G2067), .ZN(n678) );
  NAND2_X1 U771 ( .A1(n679), .A2(n678), .ZN(n682) );
  NOR2_X1 U772 ( .A1(n925), .A2(n682), .ZN(n680) );
  NOR2_X1 U773 ( .A1(n681), .A2(n680), .ZN(n696) );
  NAND2_X1 U774 ( .A1(n682), .A2(n925), .ZN(n694) );
  XOR2_X1 U775 ( .A(KEYINPUT26), .B(KEYINPUT91), .Z(n687) );
  OR2_X1 U776 ( .A1(n687), .A2(G1996), .ZN(n683) );
  NAND2_X1 U777 ( .A1(n684), .A2(n683), .ZN(n692) );
  INV_X1 U778 ( .A(G1341), .ZN(n938) );
  NAND2_X1 U779 ( .A1(n938), .A2(n687), .ZN(n685) );
  NAND2_X1 U780 ( .A1(n685), .A2(n720), .ZN(n690) );
  AND2_X1 U781 ( .A1(n686), .A2(G1996), .ZN(n688) );
  NAND2_X1 U782 ( .A1(n688), .A2(n687), .ZN(n689) );
  NAND2_X1 U783 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U784 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U785 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U786 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U787 ( .A(n697), .B(KEYINPUT92), .Z(n703) );
  INV_X1 U788 ( .A(KEYINPUT28), .ZN(n701) );
  NAND2_X1 U789 ( .A1(n698), .A2(G299), .ZN(n699) );
  XNOR2_X1 U790 ( .A(n699), .B(KEYINPUT90), .ZN(n700) );
  XNOR2_X1 U791 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U792 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U793 ( .A(KEYINPUT29), .B(n704), .Z(n705) );
  NOR2_X1 U794 ( .A1(G2084), .A2(n720), .ZN(n733) );
  NOR2_X1 U795 ( .A1(G1966), .A2(n759), .ZN(n730) );
  NOR2_X1 U796 ( .A1(n733), .A2(n730), .ZN(n708) );
  XNOR2_X1 U797 ( .A(n708), .B(n707), .ZN(n709) );
  NAND2_X1 U798 ( .A1(n709), .A2(G8), .ZN(n710) );
  XNOR2_X1 U799 ( .A(KEYINPUT30), .B(n710), .ZN(n711) );
  NOR2_X1 U800 ( .A1(G168), .A2(n711), .ZN(n714) );
  AND2_X1 U801 ( .A1(G301), .A2(n712), .ZN(n713) );
  NOR2_X1 U802 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U803 ( .A(n715), .B(KEYINPUT31), .ZN(n716) );
  INV_X1 U804 ( .A(n731), .ZN(n719) );
  NAND2_X1 U805 ( .A1(n719), .A2(G286), .ZN(n726) );
  NOR2_X1 U806 ( .A1(G1971), .A2(n759), .ZN(n722) );
  NOR2_X1 U807 ( .A1(G2090), .A2(n720), .ZN(n721) );
  NOR2_X1 U808 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U809 ( .A(KEYINPUT96), .B(n723), .ZN(n724) );
  NAND2_X1 U810 ( .A1(n724), .A2(G303), .ZN(n725) );
  NAND2_X1 U811 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U812 ( .A1(n727), .A2(G8), .ZN(n729) );
  XOR2_X1 U813 ( .A(KEYINPUT32), .B(KEYINPUT97), .Z(n728) );
  XNOR2_X1 U814 ( .A(n729), .B(n728), .ZN(n736) );
  NOR2_X1 U815 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U816 ( .A(n732), .B(KEYINPUT95), .ZN(n734) );
  NAND2_X1 U817 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U818 ( .A(n737), .B(KEYINPUT98), .ZN(n753) );
  NOR2_X1 U819 ( .A1(G303), .A2(G1971), .ZN(n738) );
  NOR2_X1 U820 ( .A1(G1976), .A2(G288), .ZN(n906) );
  NOR2_X1 U821 ( .A1(n738), .A2(n906), .ZN(n739) );
  INV_X1 U822 ( .A(KEYINPUT33), .ZN(n743) );
  AND2_X1 U823 ( .A1(n739), .A2(n743), .ZN(n740) );
  NAND2_X1 U824 ( .A1(n753), .A2(n740), .ZN(n750) );
  NAND2_X1 U825 ( .A1(G1976), .A2(G288), .ZN(n905) );
  INV_X1 U826 ( .A(n759), .ZN(n741) );
  NAND2_X1 U827 ( .A1(n905), .A2(n741), .ZN(n742) );
  NAND2_X1 U828 ( .A1(n743), .A2(n742), .ZN(n746) );
  NAND2_X1 U829 ( .A1(n906), .A2(KEYINPUT33), .ZN(n744) );
  OR2_X1 U830 ( .A1(n744), .A2(n759), .ZN(n745) );
  NAND2_X1 U831 ( .A1(n746), .A2(n745), .ZN(n748) );
  XOR2_X1 U832 ( .A(G1981), .B(G305), .Z(n920) );
  INV_X1 U833 ( .A(n920), .ZN(n747) );
  NOR2_X1 U834 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U835 ( .A1(n750), .A2(n749), .ZN(n756) );
  NOR2_X1 U836 ( .A1(G2090), .A2(G303), .ZN(n751) );
  NAND2_X1 U837 ( .A1(G8), .A2(n751), .ZN(n752) );
  NAND2_X1 U838 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U839 ( .A1(n754), .A2(n759), .ZN(n755) );
  NOR2_X1 U840 ( .A1(G1981), .A2(G305), .ZN(n757) );
  XOR2_X1 U841 ( .A(n757), .B(KEYINPUT24), .Z(n758) );
  NAND2_X1 U842 ( .A1(n663), .A2(G104), .ZN(n760) );
  XOR2_X1 U843 ( .A(KEYINPUT81), .B(n760), .Z(n762) );
  NAND2_X1 U844 ( .A1(n545), .A2(G140), .ZN(n761) );
  NAND2_X1 U845 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U846 ( .A(KEYINPUT34), .B(n763), .ZN(n768) );
  NAND2_X1 U847 ( .A1(G116), .A2(n876), .ZN(n765) );
  NAND2_X1 U848 ( .A1(G128), .A2(n879), .ZN(n764) );
  NAND2_X1 U849 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U850 ( .A(n766), .B(KEYINPUT35), .Z(n767) );
  NOR2_X1 U851 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U852 ( .A(KEYINPUT36), .B(n769), .Z(n770) );
  XOR2_X1 U853 ( .A(KEYINPUT82), .B(n770), .Z(n869) );
  XNOR2_X1 U854 ( .A(G2067), .B(KEYINPUT37), .ZN(n805) );
  NOR2_X1 U855 ( .A1(n869), .A2(n805), .ZN(n995) );
  NOR2_X1 U856 ( .A1(n772), .A2(n771), .ZN(n807) );
  NAND2_X1 U857 ( .A1(n995), .A2(n807), .ZN(n803) );
  NAND2_X1 U858 ( .A1(G95), .A2(n663), .ZN(n774) );
  NAND2_X1 U859 ( .A1(G131), .A2(n545), .ZN(n773) );
  NAND2_X1 U860 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U861 ( .A(KEYINPUT83), .B(n775), .ZN(n779) );
  NAND2_X1 U862 ( .A1(G107), .A2(n876), .ZN(n777) );
  NAND2_X1 U863 ( .A1(G119), .A2(n879), .ZN(n776) );
  AND2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U865 ( .A1(n779), .A2(n778), .ZN(n888) );
  NAND2_X1 U866 ( .A1(G1991), .A2(n888), .ZN(n780) );
  XOR2_X1 U867 ( .A(KEYINPUT84), .B(n780), .Z(n791) );
  NAND2_X1 U868 ( .A1(n663), .A2(G105), .ZN(n781) );
  XNOR2_X1 U869 ( .A(n781), .B(KEYINPUT38), .ZN(n783) );
  NAND2_X1 U870 ( .A1(G129), .A2(n879), .ZN(n782) );
  NAND2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n786) );
  NAND2_X1 U872 ( .A1(G117), .A2(n876), .ZN(n784) );
  XNOR2_X1 U873 ( .A(KEYINPUT85), .B(n784), .ZN(n785) );
  NOR2_X1 U874 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U875 ( .A(n787), .B(KEYINPUT86), .ZN(n789) );
  NAND2_X1 U876 ( .A1(G141), .A2(n545), .ZN(n788) );
  NAND2_X1 U877 ( .A1(n789), .A2(n788), .ZN(n885) );
  AND2_X1 U878 ( .A1(n885), .A2(G1996), .ZN(n790) );
  NOR2_X1 U879 ( .A1(n791), .A2(n790), .ZN(n994) );
  INV_X1 U880 ( .A(n807), .ZN(n792) );
  NOR2_X1 U881 ( .A1(n994), .A2(n792), .ZN(n800) );
  XNOR2_X1 U882 ( .A(KEYINPUT87), .B(n800), .ZN(n793) );
  XNOR2_X1 U883 ( .A(G1986), .B(G290), .ZN(n913) );
  NAND2_X1 U884 ( .A1(n913), .A2(n807), .ZN(n794) );
  NAND2_X1 U885 ( .A1(n795), .A2(n509), .ZN(n810) );
  NOR2_X1 U886 ( .A1(G1996), .A2(n885), .ZN(n984) );
  NOR2_X1 U887 ( .A1(n888), .A2(G1991), .ZN(n796) );
  XNOR2_X1 U888 ( .A(n796), .B(KEYINPUT100), .ZN(n992) );
  NOR2_X1 U889 ( .A1(G1986), .A2(G290), .ZN(n797) );
  XOR2_X1 U890 ( .A(n797), .B(KEYINPUT99), .Z(n798) );
  NOR2_X1 U891 ( .A1(n992), .A2(n798), .ZN(n799) );
  NOR2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U893 ( .A1(n984), .A2(n801), .ZN(n802) );
  XNOR2_X1 U894 ( .A(n802), .B(KEYINPUT39), .ZN(n804) );
  NAND2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n806) );
  NAND2_X1 U896 ( .A1(n869), .A2(n805), .ZN(n1000) );
  NAND2_X1 U897 ( .A1(n806), .A2(n1000), .ZN(n808) );
  NAND2_X1 U898 ( .A1(n808), .A2(n807), .ZN(n809) );
  NAND2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U900 ( .A(n811), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U901 ( .A(G2430), .B(G2451), .Z(n813) );
  XNOR2_X1 U902 ( .A(G2446), .B(G2427), .ZN(n812) );
  XNOR2_X1 U903 ( .A(n813), .B(n812), .ZN(n820) );
  XOR2_X1 U904 ( .A(G2438), .B(G2435), .Z(n815) );
  XNOR2_X1 U905 ( .A(G2443), .B(KEYINPUT101), .ZN(n814) );
  XNOR2_X1 U906 ( .A(n815), .B(n814), .ZN(n816) );
  XOR2_X1 U907 ( .A(n816), .B(G2454), .Z(n818) );
  XNOR2_X1 U908 ( .A(G1348), .B(G1341), .ZN(n817) );
  XNOR2_X1 U909 ( .A(n818), .B(n817), .ZN(n819) );
  XNOR2_X1 U910 ( .A(n820), .B(n819), .ZN(n821) );
  NAND2_X1 U911 ( .A1(n821), .A2(G14), .ZN(n897) );
  XOR2_X1 U912 ( .A(KEYINPUT102), .B(n897), .Z(G401) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n822), .ZN(G217) );
  NAND2_X1 U914 ( .A1(G15), .A2(G2), .ZN(n823) );
  XNOR2_X1 U915 ( .A(KEYINPUT103), .B(n823), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n824), .A2(G661), .ZN(G259) );
  NAND2_X1 U917 ( .A1(G1), .A2(G3), .ZN(n826) );
  NAND2_X1 U918 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U919 ( .A(n827), .B(KEYINPUT104), .ZN(G188) );
  INV_X1 U921 ( .A(G132), .ZN(G219) );
  INV_X1 U922 ( .A(G120), .ZN(G236) );
  INV_X1 U923 ( .A(G108), .ZN(G238) );
  INV_X1 U924 ( .A(G96), .ZN(G221) );
  INV_X1 U925 ( .A(G82), .ZN(G220) );
  INV_X1 U926 ( .A(G69), .ZN(G235) );
  NOR2_X1 U927 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U928 ( .A(n830), .B(KEYINPUT105), .ZN(G261) );
  INV_X1 U929 ( .A(G261), .ZN(G325) );
  INV_X1 U930 ( .A(n831), .ZN(G319) );
  XOR2_X1 U931 ( .A(G2096), .B(KEYINPUT43), .Z(n833) );
  XNOR2_X1 U932 ( .A(G2090), .B(KEYINPUT42), .ZN(n832) );
  XNOR2_X1 U933 ( .A(n833), .B(n832), .ZN(n834) );
  XOR2_X1 U934 ( .A(n834), .B(G2678), .Z(n836) );
  XNOR2_X1 U935 ( .A(G2072), .B(G2067), .ZN(n835) );
  XNOR2_X1 U936 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U937 ( .A(KEYINPUT106), .B(G2100), .Z(n838) );
  XNOR2_X1 U938 ( .A(G2084), .B(G2078), .ZN(n837) );
  XNOR2_X1 U939 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U940 ( .A(n840), .B(n839), .ZN(G227) );
  XOR2_X1 U941 ( .A(G1986), .B(G1976), .Z(n842) );
  XNOR2_X1 U942 ( .A(G1961), .B(G1971), .ZN(n841) );
  XNOR2_X1 U943 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U944 ( .A(n843), .B(G2474), .Z(n845) );
  XNOR2_X1 U945 ( .A(G1996), .B(G1991), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U947 ( .A(KEYINPUT41), .B(G1981), .Z(n847) );
  XNOR2_X1 U948 ( .A(G1966), .B(G1956), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(G229) );
  XOR2_X1 U951 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n851) );
  NAND2_X1 U952 ( .A1(G124), .A2(n879), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n852), .B(KEYINPUT107), .ZN(n854) );
  NAND2_X1 U955 ( .A1(n876), .A2(G112), .ZN(n853) );
  NAND2_X1 U956 ( .A1(n854), .A2(n853), .ZN(n858) );
  NAND2_X1 U957 ( .A1(G100), .A2(n663), .ZN(n856) );
  NAND2_X1 U958 ( .A1(G136), .A2(n545), .ZN(n855) );
  NAND2_X1 U959 ( .A1(n856), .A2(n855), .ZN(n857) );
  NOR2_X1 U960 ( .A1(n858), .A2(n857), .ZN(G162) );
  XOR2_X1 U961 ( .A(KEYINPUT48), .B(KEYINPUT111), .Z(n860) );
  XNOR2_X1 U962 ( .A(G164), .B(KEYINPUT46), .ZN(n859) );
  XNOR2_X1 U963 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U964 ( .A(n861), .B(G162), .Z(n871) );
  NAND2_X1 U965 ( .A1(G103), .A2(n663), .ZN(n863) );
  NAND2_X1 U966 ( .A1(G139), .A2(n545), .ZN(n862) );
  NAND2_X1 U967 ( .A1(n863), .A2(n862), .ZN(n868) );
  NAND2_X1 U968 ( .A1(G115), .A2(n876), .ZN(n865) );
  NAND2_X1 U969 ( .A1(G127), .A2(n879), .ZN(n864) );
  NAND2_X1 U970 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U971 ( .A(KEYINPUT47), .B(n866), .Z(n867) );
  NOR2_X1 U972 ( .A1(n868), .A2(n867), .ZN(n979) );
  XNOR2_X1 U973 ( .A(n869), .B(n979), .ZN(n870) );
  XNOR2_X1 U974 ( .A(n871), .B(n870), .ZN(n884) );
  NAND2_X1 U975 ( .A1(n545), .A2(G142), .ZN(n872) );
  XNOR2_X1 U976 ( .A(n872), .B(KEYINPUT110), .ZN(n874) );
  NAND2_X1 U977 ( .A1(G106), .A2(n663), .ZN(n873) );
  NAND2_X1 U978 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U979 ( .A(n875), .B(KEYINPUT45), .ZN(n878) );
  NAND2_X1 U980 ( .A1(G118), .A2(n876), .ZN(n877) );
  NAND2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n882) );
  NAND2_X1 U982 ( .A1(G130), .A2(n879), .ZN(n880) );
  XNOR2_X1 U983 ( .A(KEYINPUT109), .B(n880), .ZN(n881) );
  NOR2_X1 U984 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U985 ( .A(n884), .B(n883), .Z(n887) );
  XOR2_X1 U986 ( .A(G160), .B(n885), .Z(n886) );
  XNOR2_X1 U987 ( .A(n887), .B(n886), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n890), .B(n990), .ZN(n891) );
  NOR2_X1 U990 ( .A1(G37), .A2(n891), .ZN(G395) );
  XNOR2_X1 U991 ( .A(G286), .B(n892), .ZN(n894) );
  XNOR2_X1 U992 ( .A(n925), .B(G171), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U994 ( .A(n915), .B(n895), .Z(n896) );
  NOR2_X1 U995 ( .A1(G37), .A2(n896), .ZN(G397) );
  NAND2_X1 U996 ( .A1(G319), .A2(n897), .ZN(n900) );
  NOR2_X1 U997 ( .A1(G227), .A2(G229), .ZN(n898) );
  XNOR2_X1 U998 ( .A(n898), .B(KEYINPUT49), .ZN(n899) );
  NOR2_X1 U999 ( .A1(n900), .A2(n899), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(KEYINPUT112), .B(n901), .ZN(n903) );
  NOR2_X1 U1001 ( .A1(G395), .A2(G397), .ZN(n902) );
  NAND2_X1 U1002 ( .A1(n903), .A2(n902), .ZN(G225) );
  INV_X1 U1003 ( .A(G225), .ZN(G308) );
  XNOR2_X1 U1004 ( .A(KEYINPUT56), .B(G16), .ZN(n931) );
  XOR2_X1 U1005 ( .A(G1956), .B(G299), .Z(n904) );
  NAND2_X1 U1006 ( .A1(n905), .A2(n904), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(KEYINPUT120), .B(n906), .ZN(n907) );
  NOR2_X1 U1008 ( .A1(n908), .A2(n907), .ZN(n910) );
  XOR2_X1 U1009 ( .A(G303), .B(G1971), .Z(n909) );
  NAND2_X1 U1010 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1011 ( .A(KEYINPUT121), .B(n911), .Z(n912) );
  NOR2_X1 U1012 ( .A1(n913), .A2(n912), .ZN(n914) );
  XNOR2_X1 U1013 ( .A(KEYINPUT122), .B(n914), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(G1341), .B(n915), .ZN(n916) );
  NAND2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(n924) );
  XOR2_X1 U1016 ( .A(KEYINPUT119), .B(KEYINPUT57), .Z(n922) );
  XNOR2_X1 U1017 ( .A(G1966), .B(G168), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(n918), .B(KEYINPUT118), .ZN(n919) );
  NAND2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1020 ( .A(n922), .B(n921), .Z(n923) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n929) );
  XNOR2_X1 U1022 ( .A(n925), .B(G1348), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(G301), .B(G1961), .ZN(n926) );
  NOR2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1026 ( .A1(n931), .A2(n930), .ZN(n1010) );
  XOR2_X1 U1027 ( .A(G4), .B(KEYINPUT125), .Z(n933) );
  XNOR2_X1 U1028 ( .A(G1348), .B(KEYINPUT59), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(n933), .B(n932), .ZN(n937) );
  XNOR2_X1 U1030 ( .A(G1956), .B(G20), .ZN(n935) );
  XNOR2_X1 U1031 ( .A(G1981), .B(G6), .ZN(n934) );
  NOR2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n941) );
  XOR2_X1 U1034 ( .A(KEYINPUT124), .B(n938), .Z(n939) );
  XNOR2_X1 U1035 ( .A(G19), .B(n939), .ZN(n940) );
  NOR2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1037 ( .A(KEYINPUT60), .B(n942), .ZN(n952) );
  XNOR2_X1 U1038 ( .A(G1966), .B(KEYINPUT126), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(n943), .B(G21), .ZN(n950) );
  XNOR2_X1 U1040 ( .A(G1971), .B(G22), .ZN(n945) );
  XNOR2_X1 U1041 ( .A(G24), .B(G1986), .ZN(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n947) );
  XOR2_X1 U1043 ( .A(G1976), .B(G23), .Z(n946) );
  NAND2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(KEYINPUT58), .B(n948), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n954) );
  XNOR2_X1 U1048 ( .A(G5), .B(G1961), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(n955), .B(KEYINPUT61), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(G16), .B(KEYINPUT123), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(G11), .A2(n958), .ZN(n1008) );
  XOR2_X1 U1054 ( .A(KEYINPUT116), .B(G34), .Z(n960) );
  XNOR2_X1 U1055 ( .A(G2084), .B(KEYINPUT54), .ZN(n959) );
  XNOR2_X1 U1056 ( .A(n960), .B(n959), .ZN(n975) );
  XNOR2_X1 U1057 ( .A(G2090), .B(G35), .ZN(n973) );
  XOR2_X1 U1058 ( .A(G1991), .B(G25), .Z(n961) );
  NAND2_X1 U1059 ( .A1(n961), .A2(G28), .ZN(n970) );
  XNOR2_X1 U1060 ( .A(G2072), .B(G33), .ZN(n963) );
  XNOR2_X1 U1061 ( .A(G1996), .B(G32), .ZN(n962) );
  NOR2_X1 U1062 ( .A1(n963), .A2(n962), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(G2067), .B(G26), .ZN(n966) );
  XNOR2_X1 U1064 ( .A(G27), .B(n964), .ZN(n965) );
  NOR2_X1 U1065 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1066 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1068 ( .A(KEYINPUT53), .B(n971), .ZN(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1071 ( .A(KEYINPUT117), .B(n976), .ZN(n977) );
  NOR2_X1 U1072 ( .A1(G29), .A2(n977), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(n978), .B(KEYINPUT55), .ZN(n1006) );
  XOR2_X1 U1074 ( .A(KEYINPUT52), .B(KEYINPUT115), .Z(n1003) );
  XOR2_X1 U1075 ( .A(G2072), .B(n979), .Z(n981) );
  XOR2_X1 U1076 ( .A(G164), .B(G2078), .Z(n980) );
  NOR2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1078 ( .A(KEYINPUT50), .B(n982), .ZN(n987) );
  XOR2_X1 U1079 ( .A(G2090), .B(G162), .Z(n983) );
  NOR2_X1 U1080 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1081 ( .A(KEYINPUT51), .B(n985), .Z(n986) );
  NAND2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n999) );
  XOR2_X1 U1083 ( .A(G160), .B(G2084), .Z(n988) );
  XNOR2_X1 U1084 ( .A(KEYINPUT113), .B(n988), .ZN(n989) );
  NAND2_X1 U1085 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1089 ( .A(KEYINPUT114), .B(n997), .Z(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(n1003), .B(n1002), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(G29), .A2(n1004), .ZN(n1005) );
  NAND2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1096 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(n1011), .B(KEYINPUT127), .ZN(n1012) );
  XNOR2_X1 U1098 ( .A(KEYINPUT62), .B(n1012), .ZN(G311) );
  INV_X1 U1099 ( .A(G311), .ZN(G150) );
endmodule

