//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 1 0 0 0 1 0 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  XOR2_X1   g001(.A(KEYINPUT27), .B(G183gat), .Z(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT71), .B(G190gat), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT28), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT71), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT71), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT28), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT73), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT27), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(new_n214), .A3(G183gat), .ZN(new_n215));
  INV_X1    g014(.A(G183gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT27), .B1(new_n216), .B2(KEYINPUT73), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n211), .A2(new_n212), .A3(new_n215), .A4(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(KEYINPUT74), .A2(KEYINPUT26), .ZN(new_n219));
  INV_X1    g018(.A(G169gat), .ZN(new_n220));
  INV_X1    g019(.A(G176gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(KEYINPUT74), .A2(KEYINPUT26), .ZN(new_n224));
  OAI22_X1  g023(.A1(KEYINPUT74), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .A4(new_n225), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n205), .A2(new_n206), .A3(new_n218), .A4(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n227), .B(KEYINPUT75), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT67), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n221), .A2(KEYINPUT23), .ZN(new_n230));
  OR2_X1    g029(.A1(KEYINPUT66), .A2(G169gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(KEYINPUT66), .A2(G169gat), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(G169gat), .B2(G176gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n223), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n229), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT24), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n206), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n239), .B(new_n240), .C1(G183gat), .C2(G190gat), .ZN(new_n241));
  AND2_X1   g040(.A1(G169gat), .A2(G176gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n220), .A2(new_n221), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n242), .B1(new_n243), .B2(new_n234), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n234), .A2(G176gat), .ZN(new_n245));
  AND2_X1   g044(.A1(KEYINPUT66), .A2(G169gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(KEYINPUT66), .A2(G169gat), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n244), .A2(new_n248), .A3(KEYINPUT67), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n237), .A2(new_n241), .A3(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n223), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT23), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n254), .A2(new_n255), .A3(new_n235), .A4(KEYINPUT25), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n256), .B1(KEYINPUT68), .B2(new_n242), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n206), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(KEYINPUT69), .A2(G183gat), .A3(G190gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(new_n238), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n259), .A2(KEYINPUT70), .A3(new_n238), .A4(new_n260), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n240), .B1(new_n204), .B2(G183gat), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n257), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n252), .A2(KEYINPUT72), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT72), .B1(new_n252), .B2(new_n267), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n228), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(G120gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(G113gat), .ZN(new_n272));
  INV_X1    g071(.A(G113gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(G120gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT78), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT1), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT78), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n272), .A2(new_n274), .A3(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n276), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  AND2_X1   g079(.A1(KEYINPUT76), .A2(G134gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(KEYINPUT76), .A2(G134gat), .ZN(new_n282));
  OAI21_X1  g081(.A(G127gat), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G134gat), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n283), .B(KEYINPUT77), .C1(G127gat), .C2(new_n284), .ZN(new_n285));
  OR2_X1    g084(.A1(new_n283), .A2(KEYINPUT77), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n280), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT1), .B1(new_n284), .B2(G127gat), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n275), .B(new_n288), .C1(G127gat), .C2(new_n284), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n270), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n290), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n292), .B(new_n228), .C1(new_n268), .C2(new_n269), .ZN(new_n293));
  NAND2_X1  g092(.A1(G227gat), .A2(G233gat), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n291), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT34), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT34), .ZN(new_n297));
  XOR2_X1   g096(.A(new_n294), .B(KEYINPUT64), .Z(new_n298));
  NAND4_X1  g097(.A1(new_n291), .A2(new_n297), .A3(new_n293), .A4(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n298), .B1(new_n291), .B2(new_n293), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT32), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G15gat), .B(G43gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(G71gat), .B(G99gat), .ZN(new_n306));
  XOR2_X1   g105(.A(new_n305), .B(new_n306), .Z(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(new_n301), .B2(KEYINPUT33), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n296), .B(new_n299), .C1(new_n302), .C2(new_n301), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n304), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n309), .B1(new_n304), .B2(new_n310), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n202), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n304), .A2(new_n310), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(new_n308), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n304), .A2(new_n309), .A3(new_n310), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n315), .A2(KEYINPUT36), .A3(new_n316), .ZN(new_n317));
  XOR2_X1   g116(.A(G8gat), .B(G36gat), .Z(new_n318));
  XNOR2_X1  g117(.A(new_n318), .B(G64gat), .ZN(new_n319));
  XOR2_X1   g118(.A(new_n319), .B(G92gat), .Z(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT79), .B(G204gat), .ZN(new_n322));
  OR2_X1    g121(.A1(new_n322), .A2(G197gat), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT22), .ZN(new_n324));
  INV_X1    g123(.A(G211gat), .ZN(new_n325));
  INV_X1    g124(.A(G218gat), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n322), .A2(G197gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n323), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT80), .ZN(new_n330));
  XNOR2_X1  g129(.A(G211gat), .B(G218gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n329), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n330), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n334), .A2(new_n323), .A3(new_n327), .A4(new_n328), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n337));
  NAND2_X1  g136(.A1(G226gat), .A2(G233gat), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n338), .B(KEYINPUT81), .Z(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n270), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n227), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n342), .B1(new_n252), .B2(new_n267), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(new_n339), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n336), .B1(new_n341), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n336), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n270), .A2(new_n339), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n340), .B1(new_n343), .B2(KEYINPUT29), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n321), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n227), .B(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n252), .A2(new_n267), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT72), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n252), .A2(KEYINPUT72), .A3(new_n267), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n352), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n337), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n344), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n346), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n348), .B1(new_n357), .B2(new_n340), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n336), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n360), .A2(new_n362), .A3(new_n320), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n350), .A2(new_n363), .A3(KEYINPUT30), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT30), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n365), .B(new_n321), .C1(new_n345), .C2(new_n349), .ZN(new_n366));
  XNOR2_X1  g165(.A(G155gat), .B(G162gat), .ZN(new_n367));
  XOR2_X1   g166(.A(G141gat), .B(G148gat), .Z(new_n368));
  AND2_X1   g167(.A1(KEYINPUT82), .A2(KEYINPUT2), .ZN(new_n369));
  NOR2_X1   g168(.A1(KEYINPUT82), .A2(KEYINPUT2), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n367), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G141gat), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT83), .B1(new_n373), .B2(G148gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n373), .A2(G148gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n373), .A2(KEYINPUT83), .A3(G148gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(G155gat), .A2(G162gat), .ZN(new_n378));
  OR2_X1    g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n376), .A2(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(KEYINPUT2), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n381), .B(KEYINPUT84), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n372), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n383), .A2(new_n287), .A3(new_n289), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT4), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT4), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n383), .A2(new_n287), .A3(new_n386), .A4(new_n289), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(G225gat), .A2(G233gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n389), .B(KEYINPUT85), .Z(new_n390));
  NAND2_X1  g189(.A1(new_n384), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n377), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n382), .A2(new_n367), .A3(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n372), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n395), .A2(KEYINPUT3), .B1(new_n287), .B2(new_n289), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT3), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n383), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n388), .A2(new_n391), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n290), .A2(new_n395), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT86), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n402), .A3(new_n384), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n290), .A2(KEYINPUT86), .A3(new_n395), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n403), .A2(new_n390), .A3(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n400), .A2(new_n405), .A3(KEYINPUT5), .ZN(new_n406));
  AOI22_X1  g205(.A1(new_n385), .A2(new_n387), .B1(new_n396), .B2(new_n398), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT5), .ZN(new_n408));
  INV_X1    g207(.A(new_n390), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n406), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT0), .B(G57gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(G85gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(G1gat), .B(G29gat), .ZN(new_n414));
  XOR2_X1   g213(.A(new_n413), .B(new_n414), .Z(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT6), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n406), .A2(new_n415), .A3(new_n410), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n411), .A2(KEYINPUT6), .A3(new_n416), .ZN(new_n421));
  AOI22_X1  g220(.A1(new_n364), .A2(new_n366), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(G78gat), .B(G106gat), .ZN(new_n424));
  XOR2_X1   g223(.A(new_n424), .B(G22gat), .Z(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT29), .B1(new_n383), .B2(new_n397), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n427), .A2(new_n336), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT88), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT29), .B1(new_n333), .B2(new_n335), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n395), .B1(new_n431), .B2(KEYINPUT3), .ZN(new_n432));
  OAI21_X1  g231(.A(KEYINPUT88), .B1(new_n427), .B2(new_n336), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT87), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n329), .A2(new_n331), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n323), .A2(new_n332), .A3(new_n327), .A4(new_n328), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n337), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n383), .B1(new_n438), .B2(new_n397), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n435), .B1(new_n439), .B2(new_n428), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n434), .A2(G228gat), .A3(G233gat), .A4(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT31), .B(G50gat), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT87), .B1(new_n439), .B2(new_n428), .ZN(new_n444));
  NAND2_X1  g243(.A1(G228gat), .A2(G233gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n441), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n443), .B1(new_n441), .B2(new_n446), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n426), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n441), .A2(new_n446), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n442), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n441), .A2(new_n443), .A3(new_n446), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n425), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  AOI22_X1  g254(.A1(new_n313), .A2(new_n317), .B1(new_n423), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n403), .A2(new_n404), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n409), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n458), .A2(KEYINPUT91), .A3(KEYINPUT39), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n388), .A2(new_n399), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(new_n390), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT91), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n390), .B1(new_n403), .B2(new_n404), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT39), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n459), .A2(new_n461), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT92), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT40), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR3_X1   g268(.A1(new_n407), .A2(KEYINPUT39), .A3(new_n409), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n415), .B(KEYINPUT89), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT90), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT90), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n474), .B(new_n471), .C1(new_n461), .C2(KEYINPUT39), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n466), .A2(new_n469), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n471), .B1(new_n406), .B2(new_n410), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n466), .A2(new_n473), .A3(new_n475), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(new_n467), .A3(new_n468), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n479), .A2(new_n366), .A3(new_n364), .A4(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(KEYINPUT93), .B(KEYINPUT37), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(new_n345), .B2(new_n349), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n360), .A2(new_n362), .A3(KEYINPUT37), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n485), .A3(new_n320), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT38), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n419), .A2(new_n418), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n421), .B1(new_n488), .B2(new_n477), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT38), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n347), .A2(new_n346), .A3(new_n348), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n492), .B(KEYINPUT37), .C1(new_n346), .C2(new_n359), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n484), .A2(new_n491), .A3(new_n493), .A4(new_n320), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n487), .A2(new_n490), .A3(new_n350), .A4(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n482), .A2(new_n495), .A3(new_n454), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n315), .A2(new_n422), .A3(new_n454), .A4(new_n316), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n364), .A2(new_n366), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT35), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n499), .A2(new_n500), .A3(new_n489), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n311), .A2(new_n312), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n502), .A3(new_n454), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n456), .A2(new_n496), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT104), .ZN(new_n505));
  XOR2_X1   g304(.A(G57gat), .B(G64gat), .Z(new_n506));
  INV_X1    g305(.A(KEYINPUT9), .ZN(new_n507));
  INV_X1    g306(.A(G71gat), .ZN(new_n508));
  INV_X1    g307(.A(G78gat), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(G71gat), .B(G78gat), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n506), .A2(new_n512), .A3(new_n510), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n517), .A2(KEYINPUT21), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(new_n325), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n518), .B(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(G1gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT97), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n524), .A2(KEYINPUT97), .A3(G1gat), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n527), .B(new_n528), .C1(KEYINPUT16), .C2(new_n525), .ZN(new_n529));
  INV_X1    g328(.A(G8gat), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n524), .A2(G1gat), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n530), .B1(new_n531), .B2(KEYINPUT98), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n529), .B(new_n532), .Z(new_n533));
  INV_X1    g332(.A(KEYINPUT101), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n516), .B(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT21), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n216), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n533), .A2(new_n536), .A3(new_n216), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n538), .A2(new_n539), .B1(G231gat), .B2(G233gat), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n533), .A2(new_n536), .A3(new_n216), .ZN(new_n541));
  NAND2_X1  g340(.A1(G231gat), .A2(G233gat), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n541), .A2(new_n537), .A3(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G127gat), .B(G155gat), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n544), .B(KEYINPUT20), .Z(new_n545));
  NOR3_X1   g344(.A1(new_n540), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n545), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n538), .A2(new_n539), .A3(G231gat), .A4(G233gat), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n542), .B1(new_n541), .B2(new_n537), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n522), .B1(new_n546), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n545), .B1(new_n540), .B2(new_n543), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n548), .A2(new_n549), .A3(new_n547), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n552), .A2(new_n521), .A3(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(G85gat), .A2(G92gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT7), .ZN(new_n557));
  NAND2_X1  g356(.A1(G99gat), .A2(G106gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT103), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT103), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(G99gat), .A3(G106gat), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n559), .A2(new_n561), .A3(KEYINPUT8), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n557), .B(new_n562), .C1(G85gat), .C2(G92gat), .ZN(new_n563));
  XOR2_X1   g362(.A(G99gat), .B(G106gat), .Z(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G43gat), .B(G50gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT15), .ZN(new_n567));
  NAND2_X1  g366(.A1(G29gat), .A2(G36gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT14), .ZN(new_n569));
  INV_X1    g368(.A(G29gat), .ZN(new_n570));
  INV_X1    g369(.A(G36gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n567), .B1(new_n568), .B2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n567), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n566), .A2(KEYINPUT15), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n573), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n579), .B1(KEYINPUT95), .B2(new_n572), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n580), .B1(KEYINPUT95), .B2(new_n572), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(new_n581), .A3(new_n568), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT96), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n578), .A2(new_n581), .A3(KEYINPUT96), .A4(new_n568), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n575), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT17), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI211_X1 g387(.A(KEYINPUT17), .B(new_n575), .C1(new_n584), .C2(new_n585), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n565), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n591), .B(KEYINPUT102), .Z(new_n592));
  INV_X1    g391(.A(KEYINPUT41), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OR2_X1    g393(.A1(new_n586), .A2(new_n565), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n590), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n597), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n590), .A2(new_n599), .A3(new_n594), .A4(new_n595), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n592), .A2(new_n593), .ZN(new_n602));
  XNOR2_X1  g401(.A(G190gat), .B(G218gat), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n602), .B(new_n603), .Z(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n598), .A2(new_n604), .A3(new_n600), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n505), .B1(new_n555), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n608), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n551), .A2(new_n554), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n610), .A2(new_n611), .A3(KEYINPUT104), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n504), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n533), .B1(new_n588), .B2(new_n589), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n533), .A2(new_n586), .ZN(new_n616));
  NAND2_X1  g415(.A1(G229gat), .A2(G233gat), .ZN(new_n617));
  OR2_X1    g416(.A1(KEYINPUT99), .A2(KEYINPUT18), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n615), .A2(new_n616), .A3(new_n617), .A4(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(KEYINPUT99), .A2(KEYINPUT18), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n533), .B(new_n586), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n617), .B(KEYINPUT13), .Z(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n619), .A2(new_n620), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n621), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(KEYINPUT11), .B(G169gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(G197gat), .ZN(new_n628));
  XOR2_X1   g427(.A(G113gat), .B(G141gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(KEYINPUT94), .Z(new_n631));
  XOR2_X1   g430(.A(new_n631), .B(KEYINPUT12), .Z(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n626), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n621), .A2(new_n632), .A3(new_n624), .A4(new_n625), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT108), .ZN(new_n637));
  NAND2_X1  g436(.A1(G230gat), .A2(G233gat), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n638), .B(KEYINPUT106), .Z(new_n639));
  INV_X1    g438(.A(new_n564), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n563), .B(new_n640), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n640), .A2(KEYINPUT105), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n641), .A2(new_n517), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n517), .A2(new_n642), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(new_n565), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT10), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n643), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n535), .A2(KEYINPUT10), .A3(new_n641), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n639), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n643), .A2(new_n645), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n639), .ZN(new_n652));
  XNOR2_X1  g451(.A(G120gat), .B(G148gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(G204gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT107), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(new_n221), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n650), .A2(new_n652), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n657), .B1(new_n650), .B2(new_n652), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n637), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n660), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n662), .A2(KEYINPUT108), .A3(new_n658), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n636), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n614), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n420), .A2(new_n421), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT109), .B(G1gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1324gat));
  INV_X1    g471(.A(new_n668), .ZN(new_n673));
  INV_X1    g472(.A(new_n499), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT16), .B(G8gat), .Z(new_n675));
  NAND3_X1  g474(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT110), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(KEYINPUT42), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT42), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n676), .A2(new_n677), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(G8gat), .B1(new_n668), .B2(new_n499), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n682), .A2(KEYINPUT111), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(KEYINPUT111), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n679), .B(new_n681), .C1(new_n683), .C2(new_n684), .ZN(G1325gat));
  AOI21_X1  g484(.A(G15gat), .B1(new_n673), .B2(new_n502), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n313), .A2(new_n317), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n688), .A2(G15gat), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n686), .B1(new_n673), .B2(new_n689), .ZN(G1326gat));
  NOR2_X1   g489(.A1(new_n668), .A2(new_n454), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT43), .B(G22gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  NOR4_X1   g492(.A1(new_n504), .A2(new_n611), .A3(new_n610), .A4(new_n666), .ZN(new_n694));
  INV_X1    g493(.A(new_n669), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(new_n570), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(KEYINPUT112), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT112), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n694), .A2(new_n698), .A3(new_n570), .A4(new_n695), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT45), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n703), .B1(new_n504), .B2(new_n610), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n423), .A2(new_n455), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n687), .A2(new_n496), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n498), .A2(new_n503), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n708), .A2(KEYINPUT44), .A3(new_n608), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n704), .A2(new_n709), .A3(new_n555), .A4(new_n667), .ZN(new_n710));
  OAI21_X1  g509(.A(G29gat), .B1(new_n710), .B2(new_n669), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n697), .A2(KEYINPUT45), .A3(new_n699), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n702), .A2(new_n711), .A3(new_n712), .ZN(G1328gat));
  NAND3_X1  g512(.A1(new_n694), .A2(new_n571), .A3(new_n674), .ZN(new_n714));
  XOR2_X1   g513(.A(new_n714), .B(KEYINPUT46), .Z(new_n715));
  OAI21_X1  g514(.A(G36gat), .B1(new_n710), .B2(new_n499), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(G1329gat));
  OAI21_X1  g516(.A(G43gat), .B1(new_n710), .B2(new_n687), .ZN(new_n718));
  INV_X1    g517(.A(G43gat), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n694), .A2(new_n719), .A3(new_n502), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(KEYINPUT47), .B1(new_n721), .B2(KEYINPUT113), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT113), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT47), .ZN(new_n724));
  AOI211_X1 g523(.A(new_n723), .B(new_n724), .C1(new_n718), .C2(new_n720), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n722), .A2(new_n725), .ZN(G1330gat));
  OAI21_X1  g525(.A(G50gat), .B1(new_n710), .B2(new_n454), .ZN(new_n727));
  INV_X1    g526(.A(G50gat), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n694), .A2(new_n728), .A3(new_n455), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1331gat));
  NOR2_X1   g531(.A1(new_n636), .A2(new_n665), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n614), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n669), .ZN(new_n735));
  XOR2_X1   g534(.A(KEYINPUT114), .B(G57gat), .Z(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1332gat));
  NOR2_X1   g536(.A1(new_n734), .A2(new_n499), .ZN(new_n738));
  NOR2_X1   g537(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n739));
  AND2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n741), .B1(new_n738), .B2(new_n739), .ZN(G1333gat));
  INV_X1    g541(.A(new_n502), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n508), .B1(new_n734), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n688), .A2(G71gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n734), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g546(.A1(new_n734), .A2(new_n454), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(new_n509), .ZN(G1335gat));
  NAND4_X1  g548(.A1(new_n704), .A2(new_n709), .A3(new_n555), .A4(new_n733), .ZN(new_n750));
  INV_X1    g549(.A(G85gat), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n750), .A2(new_n751), .A3(new_n669), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n708), .A2(KEYINPUT115), .A3(new_n608), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n555), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n634), .A2(new_n635), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n610), .B1(new_n706), .B2(new_n707), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n756), .B2(KEYINPUT115), .ZN(new_n757));
  OAI21_X1  g556(.A(KEYINPUT51), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n611), .B1(new_n756), .B2(KEYINPUT115), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT115), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n504), .B2(new_n610), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n759), .A2(new_n760), .A3(new_n755), .A4(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n758), .A2(new_n763), .A3(new_n695), .A4(new_n664), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n752), .B1(new_n764), .B2(new_n751), .ZN(G1336gat));
  NOR2_X1   g564(.A1(new_n499), .A2(G92gat), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n758), .A2(new_n763), .A3(new_n664), .A4(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G92gat), .B1(new_n750), .B2(new_n499), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(KEYINPUT52), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n767), .A2(new_n771), .A3(new_n768), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(G1337gat));
  OR3_X1    g572(.A1(new_n750), .A2(KEYINPUT116), .A3(new_n687), .ZN(new_n774));
  XOR2_X1   g573(.A(KEYINPUT117), .B(G99gat), .Z(new_n775));
  OAI21_X1  g574(.A(KEYINPUT116), .B1(new_n750), .B2(new_n687), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n743), .A2(new_n775), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n758), .A2(new_n763), .A3(new_n664), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1338gat));
  NOR2_X1   g579(.A1(new_n454), .A2(G106gat), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n758), .A2(new_n763), .A3(new_n664), .A4(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(G106gat), .B1(new_n750), .B2(new_n454), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT53), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n782), .A2(new_n786), .A3(new_n783), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(G1339gat));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n647), .A2(new_n639), .A3(new_n648), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(KEYINPUT54), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(new_n649), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n647), .A2(new_n648), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794));
  INV_X1    g593(.A(new_n639), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n656), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n789), .B1(new_n792), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n657), .B1(new_n649), .B2(new_n794), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n799), .B(KEYINPUT55), .C1(new_n649), .C2(new_n791), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(new_n658), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT118), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n798), .A2(KEYINPUT118), .A3(new_n800), .A4(new_n658), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n636), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n617), .B1(new_n615), .B2(new_n616), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n622), .A2(new_n623), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n630), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n635), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n664), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n608), .B1(new_n805), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n803), .A2(new_n804), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n813), .A2(new_n608), .A3(new_n809), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n555), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n609), .A2(new_n612), .A3(new_n755), .A4(new_n665), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n743), .A2(new_n455), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n819), .A2(new_n669), .A3(new_n674), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n636), .ZN(new_n821));
  XOR2_X1   g620(.A(KEYINPUT119), .B(G113gat), .Z(new_n822));
  XNOR2_X1  g621(.A(new_n821), .B(new_n822), .ZN(G1340gat));
  NAND2_X1  g622(.A1(new_n820), .A2(new_n664), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(G120gat), .ZN(G1341gat));
  AND2_X1   g624(.A1(new_n817), .A2(new_n818), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n674), .A2(new_n669), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(new_n555), .ZN(new_n829));
  NOR2_X1   g628(.A1(KEYINPUT120), .A2(G127gat), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n829), .B(new_n830), .ZN(G1342gat));
  OR2_X1    g630(.A1(new_n281), .A2(new_n282), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n820), .A2(new_n832), .A3(new_n608), .ZN(new_n833));
  XNOR2_X1  g632(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(G134gat), .B1(new_n828), .B2(new_n610), .ZN(new_n836));
  AND2_X1   g635(.A1(KEYINPUT121), .A2(KEYINPUT56), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n835), .B(new_n836), .C1(new_n833), .C2(new_n837), .ZN(G1343gat));
  NAND2_X1  g637(.A1(new_n687), .A2(new_n827), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n801), .B1(new_n634), .B2(new_n635), .ZN(new_n840));
  AND3_X1   g639(.A1(new_n664), .A2(new_n635), .A3(new_n808), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n610), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n813), .A2(new_n608), .A3(new_n809), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n611), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AND4_X1   g643(.A1(new_n609), .A2(new_n612), .A3(new_n755), .A4(new_n665), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n455), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n839), .B1(new_n846), .B2(KEYINPUT57), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n817), .A2(new_n848), .A3(new_n455), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n847), .A2(new_n849), .A3(new_n636), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(G141gat), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n688), .A2(new_n669), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n810), .B1(new_n755), .B2(new_n812), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n610), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n611), .B1(new_n856), .B2(new_n843), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n455), .B(new_n854), .C1(new_n857), .C2(new_n845), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n755), .A2(G141gat), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n454), .B1(new_n815), .B2(new_n816), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(KEYINPUT122), .A3(new_n854), .ZN(new_n863));
  AND4_X1   g662(.A1(new_n499), .A2(new_n860), .A3(new_n861), .A4(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n858), .A2(new_n674), .ZN(new_n865));
  AOI22_X1  g664(.A1(new_n850), .A2(G141gat), .B1(new_n865), .B2(new_n861), .ZN(new_n866));
  OAI22_X1  g665(.A1(new_n853), .A2(new_n864), .B1(new_n866), .B2(new_n852), .ZN(G1344gat));
  NOR2_X1   g666(.A1(new_n665), .A2(G148gat), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n860), .A2(new_n499), .A3(new_n863), .A4(new_n868), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n869), .A2(KEYINPUT123), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n869), .A2(KEYINPUT123), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n843), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n845), .B1(new_n873), .B2(new_n555), .ZN(new_n874));
  OAI21_X1  g673(.A(KEYINPUT57), .B1(new_n874), .B2(new_n454), .ZN(new_n875));
  INV_X1    g674(.A(new_n839), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n610), .A2(new_n801), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(new_n809), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n611), .B1(new_n842), .B2(new_n878), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n848), .B(new_n455), .C1(new_n879), .C2(new_n845), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n875), .A2(new_n664), .A3(new_n876), .A4(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n872), .B1(new_n881), .B2(G148gat), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n847), .A2(new_n849), .A3(new_n664), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n883), .A2(new_n872), .A3(G148gat), .ZN(new_n884));
  OAI22_X1  g683(.A1(new_n870), .A2(new_n871), .B1(new_n882), .B2(new_n884), .ZN(G1345gat));
  AND4_X1   g684(.A1(G155gat), .A2(new_n847), .A3(new_n849), .A4(new_n611), .ZN(new_n886));
  INV_X1    g685(.A(G155gat), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n860), .A2(new_n499), .A3(new_n863), .A4(new_n611), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(G1346gat));
  NAND3_X1  g688(.A1(new_n847), .A2(new_n849), .A3(new_n608), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(G162gat), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n610), .A2(G162gat), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n860), .A2(new_n499), .A3(new_n863), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n891), .A2(new_n893), .A3(KEYINPUT124), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1347gat));
  NOR2_X1   g697(.A1(new_n695), .A2(new_n499), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n819), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n231), .A2(new_n232), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n901), .A2(new_n902), .A3(new_n636), .ZN(new_n903));
  OR2_X1    g702(.A1(new_n903), .A2(KEYINPUT125), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n826), .A2(new_n899), .ZN(new_n905));
  OAI21_X1  g704(.A(G169gat), .B1(new_n905), .B2(new_n755), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n903), .A2(KEYINPUT125), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n904), .A2(new_n906), .A3(new_n907), .ZN(G1348gat));
  NAND2_X1  g707(.A1(new_n901), .A2(new_n664), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(G176gat), .ZN(G1349gat));
  OAI21_X1  g709(.A(G183gat), .B1(new_n905), .B2(new_n555), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT60), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n901), .A2(new_n611), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n911), .B(new_n912), .C1(new_n203), .C2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n216), .B1(new_n901), .B2(new_n611), .ZN(new_n915));
  NOR4_X1   g714(.A1(new_n819), .A2(new_n203), .A3(new_n555), .A4(new_n900), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT60), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n914), .A2(new_n917), .ZN(G1350gat));
  NAND4_X1  g717(.A1(new_n817), .A2(new_n818), .A3(new_n608), .A4(new_n899), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(G190gat), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(KEYINPUT126), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n919), .A2(new_n922), .A3(G190gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n921), .A2(KEYINPUT61), .A3(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT61), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n920), .A2(KEYINPUT126), .A3(new_n925), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n924), .B(new_n926), .C1(new_n204), .C2(new_n919), .ZN(G1351gat));
  NOR2_X1   g726(.A1(new_n688), .A2(new_n900), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n880), .B(new_n928), .C1(new_n862), .C2(new_n848), .ZN(new_n929));
  OAI21_X1  g728(.A(G197gat), .B1(new_n929), .B2(new_n755), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n862), .A2(new_n928), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n931), .A2(KEYINPUT127), .ZN(new_n932));
  INV_X1    g731(.A(G197gat), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(KEYINPUT127), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n930), .B1(new_n935), .B2(new_n755), .ZN(G1352gat));
  OR3_X1    g735(.A1(new_n931), .A2(G204gat), .A3(new_n665), .ZN(new_n937));
  OR2_X1    g736(.A1(new_n937), .A2(KEYINPUT62), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n875), .A2(new_n664), .A3(new_n880), .ZN(new_n939));
  INV_X1    g738(.A(new_n928), .ZN(new_n940));
  OAI21_X1  g739(.A(G204gat), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n937), .A2(KEYINPUT62), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n938), .A2(new_n941), .A3(new_n942), .ZN(G1353gat));
  NAND4_X1  g742(.A1(new_n932), .A2(new_n325), .A3(new_n611), .A4(new_n934), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n875), .A2(new_n611), .A3(new_n880), .A4(new_n928), .ZN(new_n945));
  AOI21_X1  g744(.A(KEYINPUT63), .B1(new_n945), .B2(G211gat), .ZN(new_n946));
  OAI211_X1 g745(.A(KEYINPUT63), .B(G211gat), .C1(new_n929), .C2(new_n555), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n944), .B1(new_n946), .B2(new_n948), .ZN(G1354gat));
  NOR3_X1   g748(.A1(new_n929), .A2(new_n326), .A3(new_n610), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n932), .A2(new_n608), .A3(new_n934), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n950), .B1(new_n951), .B2(new_n326), .ZN(G1355gat));
endmodule


