//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 1 1 0 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n778,
    new_n779, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  AND2_X1   g006(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n193));
  INV_X1    g007(.A(G134), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(G137), .ZN(new_n195));
  OR2_X1    g009(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n196));
  AOI21_X1  g010(.A(new_n193), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(G137), .ZN(new_n198));
  INV_X1    g012(.A(G137), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G134), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n198), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  OAI21_X1  g016(.A(G131), .B1(new_n197), .B2(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n201), .B1(new_n200), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n195), .A2(new_n193), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n205), .A2(new_n206), .A3(new_n207), .A4(new_n198), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n203), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(new_n210), .B2(G107), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(G104), .ZN(new_n214));
  INV_X1    g028(.A(G101), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(G107), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n211), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n210), .A2(G107), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n213), .A2(G104), .ZN(new_n219));
  OAI21_X1  g033(.A(G101), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G143), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT1), .B1(new_n221), .B2(G146), .ZN(new_n222));
  INV_X1    g036(.A(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G143), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n221), .A2(G146), .ZN(new_n225));
  AOI22_X1  g039(.A1(new_n222), .A2(G128), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G128), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n228), .A2(new_n224), .A3(new_n225), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n217), .B(new_n220), .C1(new_n226), .C2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT10), .ZN(new_n231));
  AND3_X1   g045(.A1(new_n230), .A2(KEYINPUT76), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT76), .B1(new_n230), .B2(new_n231), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n224), .A2(new_n225), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT65), .B(G128), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT1), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n237), .B1(G143), .B2(new_n223), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n235), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(G143), .B(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(new_n228), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n231), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT77), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n217), .A2(new_n220), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n243), .B1(new_n217), .B2(new_n220), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n242), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n211), .A2(new_n214), .A3(new_n216), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT75), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n247), .A2(new_n248), .A3(G101), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n248), .B1(new_n247), .B2(G101), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n217), .A2(KEYINPUT4), .ZN(new_n251));
  NOR3_X1   g065(.A1(new_n249), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT0), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n224), .B(new_n225), .C1(new_n253), .C2(new_n227), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n253), .A2(new_n227), .ZN(new_n255));
  NOR2_X1   g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n254), .B1(new_n257), .B2(new_n240), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n247), .A2(new_n259), .A3(G101), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n246), .B1(new_n252), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n209), .B1(new_n234), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n217), .A2(new_n220), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT77), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n217), .A2(new_n220), .A3(new_n243), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n247), .A2(G101), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(KEYINPUT75), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n217), .A2(KEYINPUT4), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n247), .A2(new_n248), .A3(G101), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n258), .A2(new_n260), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n267), .A2(new_n242), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n226), .A2(new_n229), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n231), .B1(new_n275), .B2(new_n264), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT76), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n230), .A2(KEYINPUT76), .A3(new_n231), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n209), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n274), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(G110), .B(G140), .ZN(new_n283));
  INV_X1    g097(.A(G953), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n284), .A2(G227), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n283), .B(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n263), .A2(new_n282), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n239), .A2(new_n241), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n217), .A2(new_n220), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n230), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n209), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT12), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n292), .A2(KEYINPUT12), .A3(new_n209), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n282), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT78), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n282), .A3(KEYINPUT78), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n289), .B1(new_n302), .B2(new_n286), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n192), .B1(new_n303), .B2(G469), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT69), .B(G902), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n297), .A2(new_n282), .A3(new_n287), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n287), .B1(new_n263), .B2(new_n282), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT79), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AOI211_X1 g123(.A(KEYINPUT79), .B(new_n287), .C1(new_n263), .C2(new_n282), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n190), .B(new_n305), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n189), .B1(new_n304), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(G237), .A2(G953), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(G143), .A3(G214), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(G143), .B1(new_n313), .B2(G214), .ZN(new_n316));
  OAI21_X1  g130(.A(G131), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT17), .ZN(new_n318));
  INV_X1    g132(.A(G237), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(new_n284), .A3(G214), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n221), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(new_n207), .A3(new_n314), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n317), .A2(new_n318), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G125), .ZN(new_n325));
  INV_X1    g139(.A(G125), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G140), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT72), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n325), .A2(new_n327), .A3(new_n328), .A4(KEYINPUT16), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n325), .A2(new_n327), .A3(KEYINPUT16), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT72), .B1(new_n325), .B2(KEYINPUT16), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G146), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n223), .B(new_n329), .C1(new_n330), .C2(new_n331), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n321), .A2(new_n314), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(KEYINPUT17), .A3(G131), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n323), .A2(new_n333), .A3(new_n334), .A4(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(G113), .B(G122), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(new_n210), .ZN(new_n339));
  NAND2_X1  g153(.A1(KEYINPUT18), .A2(G131), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n325), .A2(new_n327), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G146), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n325), .A2(new_n327), .A3(new_n223), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n335), .A2(new_n341), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT86), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n315), .A2(new_n316), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n346), .B1(new_n347), .B2(new_n340), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n335), .A2(KEYINPUT86), .A3(new_n341), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n337), .A2(new_n339), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n317), .A2(new_n322), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT19), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n342), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n325), .A2(new_n327), .A3(KEYINPUT19), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n333), .B(new_n352), .C1(new_n356), .C2(G146), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n339), .B1(new_n357), .B2(new_n350), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n351), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(G475), .A2(G902), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT20), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT87), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n364), .B1(new_n351), .B2(new_n358), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n337), .A2(new_n350), .A3(new_n339), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n325), .A2(new_n327), .A3(KEYINPUT16), .ZN(new_n367));
  OR3_X1    g181(.A1(new_n326), .A2(KEYINPUT16), .A3(G140), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n368), .A3(KEYINPUT72), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n223), .B1(new_n369), .B2(new_n329), .ZN(new_n370));
  AOI21_X1  g184(.A(G146), .B1(new_n354), .B2(new_n355), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n347), .A2(new_n346), .A3(new_n340), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT86), .B1(new_n335), .B2(new_n341), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AOI22_X1  g189(.A1(new_n372), .A2(new_n352), .B1(new_n375), .B2(new_n345), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n366), .B(KEYINPUT87), .C1(new_n376), .C2(new_n339), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n365), .A2(new_n360), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n363), .B1(new_n378), .B2(KEYINPUT20), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n339), .B1(new_n337), .B2(new_n350), .ZN(new_n381));
  OR2_X1    g195(.A1(new_n351), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n191), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G475), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  AOI211_X1 g199(.A(new_n284), .B(new_n305), .C1(G234), .C2(G237), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT21), .B(G898), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G952), .ZN(new_n389));
  AOI211_X1 g203(.A(G953), .B(new_n389), .C1(G234), .C2(G237), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  XOR2_X1   g206(.A(new_n392), .B(KEYINPUT89), .Z(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G217), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n187), .A2(new_n395), .A3(G953), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G122), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G116), .ZN(new_n399));
  INV_X1    g213(.A(G116), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(G122), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n399), .B(new_n401), .C1(KEYINPUT14), .C2(new_n213), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n213), .B1(new_n399), .B2(KEYINPUT14), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n400), .A2(G122), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n398), .A2(G116), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n227), .A2(KEYINPUT65), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT65), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G128), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n407), .A2(new_n409), .A3(G143), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n221), .A2(G128), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n410), .A2(new_n194), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n194), .B1(new_n410), .B2(new_n411), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n402), .B(new_n406), .C1(new_n412), .C2(new_n413), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n407), .A2(new_n409), .A3(G143), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT13), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(new_n227), .B2(G143), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n221), .A2(KEYINPUT13), .A3(G128), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G134), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n410), .A2(new_n194), .A3(new_n411), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n399), .A2(new_n401), .A3(G107), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n213), .B1(new_n404), .B2(new_n405), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n420), .A2(new_n421), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT88), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n414), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n425), .B1(new_n414), .B2(new_n424), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n397), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n414), .A2(new_n424), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT88), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n414), .A2(new_n424), .A3(new_n425), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n430), .A2(new_n396), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n428), .A2(new_n432), .A3(new_n305), .ZN(new_n433));
  INV_X1    g247(.A(G478), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n434), .A2(KEYINPUT15), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n433), .B(new_n435), .ZN(new_n436));
  NOR3_X1   g250(.A1(new_n385), .A2(new_n394), .A3(new_n436), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n312), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT81), .ZN(new_n439));
  INV_X1    g253(.A(G119), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT66), .B1(new_n440), .B2(G116), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT66), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(new_n400), .A3(G119), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n440), .A2(G116), .ZN(new_n445));
  INV_X1    g259(.A(G113), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT2), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT2), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G113), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n444), .A2(new_n445), .A3(new_n450), .ZN(new_n451));
  OAI21_X1  g265(.A(G113), .B1(new_n445), .B2(KEYINPUT5), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n400), .A2(G119), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n441), .B2(new_n443), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n452), .B1(new_n454), .B2(KEYINPUT5), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT80), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n451), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT5), .ZN(new_n458));
  AOI211_X1 g272(.A(new_n458), .B(new_n453), .C1(new_n443), .C2(new_n441), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT80), .B1(new_n459), .B2(new_n452), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n457), .A2(new_n267), .A3(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n454), .B(new_n450), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n272), .A2(new_n462), .A3(new_n260), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n439), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n461), .A2(new_n463), .A3(new_n439), .ZN(new_n466));
  XNOR2_X1  g280(.A(G110), .B(G122), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n465), .A2(KEYINPUT6), .A3(new_n466), .A4(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT6), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n461), .A2(new_n463), .A3(new_n467), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT82), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n461), .A2(new_n463), .A3(KEYINPUT82), .A4(new_n467), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n470), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n461), .A2(new_n463), .A3(new_n439), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n476), .A2(new_n464), .A3(new_n467), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n469), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n258), .A2(G125), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n407), .A2(new_n409), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n222), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n229), .B1(new_n235), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n479), .B1(new_n482), .B2(G125), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n284), .A2(G224), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n483), .B(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n478), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(KEYINPUT84), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n479), .B(new_n487), .C1(G125), .C2(new_n482), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n484), .A2(KEYINPUT7), .ZN(new_n489));
  XOR2_X1   g303(.A(new_n488), .B(new_n489), .Z(new_n490));
  AND2_X1   g304(.A1(new_n459), .A2(KEYINPUT83), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n459), .A2(KEYINPUT83), .ZN(new_n492));
  NOR3_X1   g306(.A1(new_n491), .A2(new_n492), .A3(new_n452), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n291), .B1(new_n493), .B2(new_n451), .ZN(new_n494));
  XOR2_X1   g308(.A(new_n467), .B(KEYINPUT8), .Z(new_n495));
  AND2_X1   g309(.A1(new_n457), .A2(new_n460), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n495), .B1(new_n496), .B2(new_n264), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n490), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n473), .A2(new_n474), .ZN(new_n499));
  AOI21_X1  g313(.A(G902), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n486), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(G210), .B1(G237), .B2(G902), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n486), .A2(new_n500), .A3(new_n502), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(G214), .B1(G237), .B2(G902), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT85), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AND3_X1   g322(.A1(new_n486), .A2(new_n500), .A3(new_n502), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n502), .B1(new_n486), .B2(new_n500), .ZN(new_n510));
  OAI211_X1 g324(.A(KEYINPUT85), .B(new_n507), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n438), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT90), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT85), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n509), .A2(new_n510), .ZN(new_n517));
  INV_X1    g331(.A(new_n507), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n511), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(KEYINPUT90), .A3(new_n438), .ZN(new_n521));
  AND2_X1   g335(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n208), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n199), .A2(G134), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n524), .B1(new_n193), .B2(new_n195), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n207), .B1(new_n525), .B2(new_n205), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n258), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n454), .A2(new_n450), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n451), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(G131), .B1(new_n195), .B2(new_n524), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n290), .A2(new_n208), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n527), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT28), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n208), .A2(new_n530), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n536), .A2(new_n482), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n235), .B1(new_n255), .B2(new_n256), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n203), .A2(new_n208), .B1(new_n538), .B2(new_n254), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n462), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n533), .B1(new_n540), .B2(new_n532), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT68), .B1(new_n535), .B2(new_n541), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n537), .A2(new_n539), .A3(new_n462), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n529), .B1(new_n527), .B2(new_n531), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT28), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT68), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XOR2_X1   g361(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n548));
  NAND2_X1  g362(.A1(new_n313), .A2(G210), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n548), .B(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT26), .B(G101), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n550), .B(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n542), .A2(new_n547), .A3(new_n553), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n537), .A2(new_n539), .A3(KEYINPUT30), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT30), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n556), .B1(new_n527), .B2(new_n531), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n462), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n532), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT29), .B1(new_n559), .B2(new_n552), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n545), .A2(new_n534), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n553), .A2(KEYINPUT29), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n305), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI211_X1 g378(.A(KEYINPUT70), .B(G472), .C1(new_n561), .C2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT70), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n564), .B1(new_n554), .B2(new_n560), .ZN(new_n567));
  INV_X1    g381(.A(G472), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n542), .A2(new_n547), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n558), .A2(new_n532), .A3(new_n553), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT31), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT30), .B1(new_n537), .B2(new_n539), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n527), .A2(new_n556), .A3(new_n531), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n543), .B1(new_n576), .B2(new_n462), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(KEYINPUT31), .A3(new_n553), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n570), .A2(new_n552), .B1(new_n573), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(G472), .A2(G902), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT32), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n573), .A2(new_n578), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n546), .B1(new_n545), .B2(new_n534), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n541), .A2(KEYINPUT68), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n552), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT32), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(new_n588), .A3(new_n580), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n565), .A2(new_n569), .B1(new_n582), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT25), .ZN(new_n591));
  INV_X1    g405(.A(new_n305), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT22), .B(G137), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n284), .A2(G221), .A3(G234), .ZN(new_n594));
  XOR2_X1   g408(.A(new_n593), .B(new_n594), .Z(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT23), .B1(new_n227), .B2(G119), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n440), .B2(G128), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT23), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n407), .A2(new_n409), .A3(G119), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(G110), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT24), .B(G110), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT71), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n236), .A2(new_n605), .A3(G119), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT71), .B1(new_n227), .B2(G119), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n236), .B2(G119), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n604), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n334), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n602), .B(new_n610), .C1(new_n611), .C2(new_n370), .ZN(new_n612));
  INV_X1    g426(.A(new_n600), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n606), .B(new_n603), .C1(new_n613), .C2(new_n608), .ZN(new_n614));
  INV_X1    g428(.A(G110), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n598), .B(new_n615), .C1(new_n599), .C2(new_n600), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n344), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n332), .B2(G146), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n612), .A2(new_n620), .A3(KEYINPUT73), .ZN(new_n621));
  AOI21_X1  g435(.A(KEYINPUT73), .B1(new_n612), .B2(new_n620), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n596), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n612), .A2(new_n620), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n595), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n592), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n591), .B1(new_n626), .B2(KEYINPUT74), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT74), .ZN(new_n628));
  INV_X1    g442(.A(new_n625), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT73), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n612), .A2(new_n620), .A3(KEYINPUT73), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n629), .B1(new_n633), .B2(new_n596), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n628), .B(KEYINPUT25), .C1(new_n634), .C2(new_n592), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n395), .B1(new_n305), .B2(G234), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n627), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n634), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n636), .A2(G902), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n590), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n522), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT91), .B(G101), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G3));
  NAND3_X1  g459(.A1(new_n504), .A2(KEYINPUT92), .A3(new_n505), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT92), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n518), .B1(new_n510), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n383), .A2(G475), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n592), .A2(new_n434), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT93), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n428), .A2(new_n432), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT33), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n428), .A2(new_n432), .A3(new_n654), .A4(KEYINPUT33), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n433), .A2(new_n434), .ZN(new_n660));
  OAI22_X1  g474(.A1(new_n651), .A2(new_n379), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(KEYINPUT94), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT94), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n394), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n650), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n587), .A2(new_n305), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(G472), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n587), .A2(new_n580), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n669), .A2(new_n670), .A3(new_n640), .A4(new_n637), .ZN(new_n671));
  INV_X1    g485(.A(new_n192), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n297), .A2(new_n282), .A3(KEYINPUT78), .ZN(new_n673));
  AOI21_X1  g487(.A(KEYINPUT78), .B1(new_n297), .B2(new_n282), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n286), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n288), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n311), .B(new_n672), .C1(new_n190), .C2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n188), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n671), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n667), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT34), .B(G104), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G6));
  OR2_X1    g497(.A1(new_n378), .A2(KEYINPUT20), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n378), .A2(KEYINPUT20), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n651), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n393), .B(KEYINPUT95), .Z(new_n687));
  NAND3_X1  g501(.A1(new_n686), .A2(new_n436), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT96), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n650), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(new_n680), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT35), .B(G107), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G9));
  AND2_X1   g508(.A1(new_n669), .A2(new_n670), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n596), .A2(KEYINPUT36), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n633), .B(new_n696), .Z(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n639), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n637), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT97), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n522), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT37), .B(G110), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT98), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n703), .B(new_n705), .ZN(G12));
  XNOR2_X1  g520(.A(new_n378), .B(KEYINPUT20), .ZN(new_n707));
  INV_X1    g521(.A(G900), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n386), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n391), .ZN(new_n710));
  XOR2_X1   g524(.A(new_n710), .B(KEYINPUT99), .Z(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n707), .A2(new_n384), .A3(new_n436), .A4(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT100), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n686), .A2(KEYINPUT100), .A3(new_n436), .A4(new_n712), .ZN(new_n716));
  AND4_X1   g530(.A1(new_n646), .A2(new_n648), .A3(new_n715), .A4(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n699), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n590), .A2(new_n678), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G128), .ZN(G30));
  XOR2_X1   g535(.A(KEYINPUT102), .B(KEYINPUT39), .Z(new_n722));
  XNOR2_X1  g536(.A(new_n711), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n312), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(KEYINPUT40), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n506), .B(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n385), .A2(new_n436), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n699), .A2(new_n728), .A3(new_n518), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n559), .A2(new_n553), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n543), .A2(new_n544), .ZN(new_n731));
  AOI21_X1  g545(.A(G902), .B1(new_n731), .B2(new_n552), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n568), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n582), .B2(new_n589), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n729), .A2(new_n735), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n725), .A2(new_n727), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n221), .ZN(G45));
  NOR2_X1   g552(.A1(new_n661), .A2(new_n711), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n646), .A2(new_n648), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT103), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT103), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n646), .A2(new_n648), .A3(new_n742), .A4(new_n739), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n741), .A2(new_n719), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G146), .ZN(G48));
  OAI21_X1  g559(.A(new_n305), .B1(new_n309), .B2(new_n310), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(G469), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n747), .A2(new_n188), .A3(new_n311), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n590), .A2(new_n641), .A3(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n667), .A2(new_n750), .ZN(new_n751));
  XOR2_X1   g565(.A(KEYINPUT41), .B(G113), .Z(new_n752));
  XNOR2_X1  g566(.A(new_n751), .B(new_n752), .ZN(G15));
  NOR2_X1   g567(.A1(new_n691), .A2(new_n750), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n400), .ZN(G18));
  AND3_X1   g569(.A1(new_n747), .A2(new_n188), .A3(new_n311), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n646), .A2(new_n756), .A3(new_n648), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n590), .A2(new_n718), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n757), .A2(new_n437), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G119), .ZN(G21));
  INV_X1    g574(.A(KEYINPUT105), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n649), .A2(new_n728), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n641), .A2(KEYINPUT104), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT104), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n637), .A2(new_n764), .A3(new_n640), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n562), .A2(new_n552), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n581), .B1(new_n583), .B2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n668), .B2(G472), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n766), .A2(new_n687), .A3(new_n756), .A4(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n761), .B1(new_n762), .B2(new_n770), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n766), .A2(new_n769), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n649), .A2(new_n728), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n756), .A2(new_n687), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n772), .A2(new_n773), .A3(KEYINPUT105), .A4(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G122), .ZN(G24));
  AND3_X1   g591(.A1(new_n739), .A2(new_n769), .A3(new_n699), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n757), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G125), .ZN(G27));
  NAND3_X1  g594(.A1(new_n504), .A2(new_n507), .A3(new_n505), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(new_n678), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n642), .A2(new_n782), .A3(new_n739), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT42), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n582), .A2(new_n589), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT106), .ZN(new_n787));
  AOI22_X1  g601(.A1(new_n786), .A2(new_n787), .B1(new_n569), .B2(new_n565), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n582), .A2(KEYINPUT106), .A3(new_n589), .ZN(new_n789));
  AOI22_X1  g603(.A1(new_n788), .A2(new_n789), .B1(new_n763), .B2(new_n765), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n661), .A2(new_n784), .A3(new_n711), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n312), .A2(new_n517), .A3(new_n791), .A4(new_n507), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT107), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n588), .B1(new_n587), .B2(new_n580), .ZN(new_n795));
  AOI211_X1 g609(.A(KEYINPUT32), .B(new_n581), .C1(new_n583), .C2(new_n586), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n787), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n565), .A2(new_n569), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n797), .A2(new_n798), .A3(new_n789), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n766), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT107), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n800), .A2(new_n801), .A3(new_n792), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n785), .B1(new_n794), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G131), .ZN(G33));
  NAND4_X1  g618(.A1(new_n642), .A2(new_n782), .A3(new_n715), .A4(new_n716), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G134), .ZN(G36));
  NAND2_X1  g620(.A1(new_n303), .A2(KEYINPUT45), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT45), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n676), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n807), .A2(new_n809), .A3(G469), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT108), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n807), .A2(new_n809), .A3(KEYINPUT108), .A4(G469), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n192), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OR3_X1    g628(.A1(new_n814), .A2(KEYINPUT109), .A3(KEYINPUT46), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT109), .B1(new_n814), .B2(KEYINPUT46), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n814), .A2(KEYINPUT46), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n815), .A2(new_n311), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n818), .A2(new_n188), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n695), .A2(new_n718), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n651), .A2(new_n379), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT110), .ZN(new_n822));
  OAI221_X1 g636(.A(new_n821), .B1(new_n822), .B2(KEYINPUT43), .C1(new_n660), .C2(new_n659), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n659), .A2(new_n660), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n385), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(KEYINPUT110), .B(KEYINPUT43), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n820), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT44), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n828), .A2(KEYINPUT111), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n781), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n831), .B1(new_n828), .B2(new_n829), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT111), .B1(new_n828), .B2(new_n829), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n830), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n819), .A2(new_n834), .A3(new_n723), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(G137), .ZN(G39));
  XOR2_X1   g650(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n837));
  AND3_X1   g651(.A1(new_n818), .A2(new_n188), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT112), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(KEYINPUT47), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n818), .B2(new_n188), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n831), .A2(new_n590), .A3(new_n641), .A4(new_n739), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n838), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(new_n324), .ZN(G42));
  AND2_X1   g658(.A1(new_n827), .A2(new_n390), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n781), .A2(new_n748), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n845), .A2(new_n790), .A3(new_n846), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n847), .B(KEYINPUT48), .Z(new_n848));
  NOR2_X1   g662(.A1(new_n641), .A2(new_n391), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n846), .A2(new_n734), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n850), .B1(new_n665), .B2(new_n663), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n845), .A2(new_n772), .ZN(new_n852));
  INV_X1    g666(.A(new_n757), .ZN(new_n853));
  OAI211_X1 g667(.A(G952), .B(new_n284), .C1(new_n852), .C2(new_n853), .ZN(new_n854));
  OR3_X1    g668(.A1(new_n848), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n727), .A2(new_n518), .A3(new_n756), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT50), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n845), .A2(new_n699), .A3(new_n769), .A4(new_n846), .ZN(new_n859));
  INV_X1    g673(.A(new_n850), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n821), .A3(new_n824), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n858), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT51), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n747), .A2(new_n311), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n189), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n866), .B1(new_n838), .B2(new_n841), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n852), .A2(new_n781), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n855), .B1(new_n864), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT115), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n818), .A2(new_n188), .A3(new_n837), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n871), .B(new_n872), .C1(new_n819), .C2(new_n840), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT115), .B1(new_n838), .B2(new_n841), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n873), .A2(new_n874), .A3(new_n866), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n862), .B1(new_n875), .B2(new_n868), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n870), .B1(new_n876), .B2(KEYINPUT51), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT116), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT116), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n879), .B(new_n870), .C1(new_n876), .C2(KEYINPUT51), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n515), .B(new_n521), .C1(new_n702), .C2(new_n642), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n749), .B(new_n650), .C1(new_n690), .C2(new_n666), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n821), .A2(new_n436), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n671), .A2(new_n678), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n520), .A2(new_n687), .A3(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n882), .A2(new_n885), .A3(new_n759), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n662), .B(new_n687), .C1(new_n508), .C2(new_n512), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT113), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n520), .A2(KEYINPUT113), .A3(new_n662), .A4(new_n687), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(new_n679), .A3(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n881), .A2(new_n886), .A3(new_n891), .A4(new_n776), .ZN(new_n892));
  AOI22_X1  g706(.A1(new_n719), .A2(new_n717), .B1(new_n757), .B2(new_n778), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT52), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n734), .A2(new_n699), .A3(new_n711), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n773), .A2(new_n312), .A3(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n893), .A2(new_n894), .A3(new_n744), .A4(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n686), .ZN(new_n898));
  NOR4_X1   g712(.A1(new_n781), .A2(new_n436), .A3(new_n898), .A4(new_n711), .ZN(new_n899));
  AOI22_X1  g713(.A1(new_n899), .A2(new_n719), .B1(new_n778), .B2(new_n782), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n803), .A2(new_n897), .A3(new_n805), .A4(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n892), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n893), .A2(new_n744), .A3(new_n896), .ZN(new_n903));
  XOR2_X1   g717(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n904));
  AND2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT53), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n903), .A2(KEYINPUT52), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT53), .ZN(new_n910));
  NOR4_X1   g724(.A1(new_n892), .A2(new_n901), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(KEYINPUT54), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n892), .ZN(new_n913));
  INV_X1    g727(.A(new_n901), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT53), .A4(new_n906), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT54), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n892), .A2(new_n901), .A3(new_n909), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n915), .B(new_n916), .C1(new_n917), .C2(KEYINPUT53), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n878), .A2(new_n880), .A3(new_n912), .A4(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(G952), .A2(G953), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT117), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n865), .B(KEYINPUT49), .ZN(new_n923));
  AND4_X1   g737(.A1(new_n507), .A2(new_n734), .A3(new_n188), .A4(new_n825), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n727), .A2(new_n923), .A3(new_n766), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n922), .A2(new_n925), .ZN(G75));
  NAND2_X1  g740(.A1(new_n902), .A2(new_n908), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n910), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n305), .B1(new_n928), .B2(new_n915), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n503), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT56), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n478), .B(new_n485), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT55), .Z(new_n933));
  AND3_X1   g747(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(new_n930), .B2(new_n931), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n389), .A2(G953), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT118), .ZN(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n934), .A2(new_n935), .A3(new_n938), .ZN(G51));
  NOR2_X1   g753(.A1(new_n309), .A2(new_n310), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT53), .B1(new_n902), .B2(new_n908), .ZN(new_n941));
  NOR4_X1   g755(.A1(new_n892), .A2(new_n901), .A3(new_n905), .A4(new_n910), .ZN(new_n942));
  OAI21_X1  g756(.A(KEYINPUT54), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n918), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n192), .B(KEYINPUT57), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n940), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OR2_X1    g760(.A1(new_n946), .A2(KEYINPUT119), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n812), .A2(new_n813), .ZN(new_n948));
  AOI22_X1  g762(.A1(new_n946), .A2(KEYINPUT119), .B1(new_n948), .B2(new_n929), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n938), .B1(new_n947), .B2(new_n949), .ZN(G54));
  AND2_X1   g764(.A1(KEYINPUT58), .A2(G475), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n592), .B(new_n951), .C1(new_n941), .C2(new_n942), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n365), .A2(new_n377), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n938), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(new_n953), .B2(new_n952), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n955), .B(KEYINPUT120), .Z(G60));
  INV_X1    g770(.A(KEYINPUT121), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n657), .A2(new_n658), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(G478), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT59), .Z(new_n961));
  NOR2_X1   g775(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n957), .B1(new_n944), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n962), .ZN(new_n964));
  AOI211_X1 g778(.A(KEYINPUT121), .B(new_n964), .C1(new_n943), .C2(new_n918), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n961), .B1(new_n912), .B2(new_n918), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n937), .B1(new_n967), .B2(new_n958), .ZN(new_n968));
  OAI21_X1  g782(.A(KEYINPUT122), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n961), .ZN(new_n970));
  INV_X1    g784(.A(new_n918), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n913), .A2(new_n914), .A3(new_n906), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(new_n910), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n917), .A2(KEYINPUT53), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n916), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n970), .B1(new_n971), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n938), .B1(new_n976), .B2(new_n959), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT122), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n977), .B(new_n978), .C1(new_n963), .C2(new_n965), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n969), .A2(new_n979), .ZN(G63));
  XNOR2_X1  g794(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n981));
  NAND2_X1  g795(.A1(G217), .A2(G902), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n983), .B1(new_n928), .B2(new_n915), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n697), .ZN(new_n985));
  OAI211_X1 g799(.A(new_n985), .B(new_n937), .C1(new_n638), .C2(new_n984), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT123), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n986), .A2(new_n987), .A3(KEYINPUT61), .ZN(new_n988));
  AOI21_X1  g802(.A(KEYINPUT61), .B1(new_n986), .B2(new_n987), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n988), .A2(new_n989), .ZN(G66));
  INV_X1    g804(.A(new_n387), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n284), .B1(new_n991), .B2(G224), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(new_n892), .B2(new_n284), .ZN(new_n993));
  INV_X1    g807(.A(new_n478), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n994), .B1(G898), .B2(new_n284), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n993), .B(new_n995), .Z(G69));
  OR3_X1    g810(.A1(new_n838), .A2(new_n841), .A3(new_n842), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n893), .A2(new_n744), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n737), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT62), .ZN(new_n1000));
  INV_X1    g814(.A(new_n724), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n883), .A2(new_n661), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n1001), .A2(new_n642), .A3(new_n831), .A4(new_n1002), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n997), .A2(new_n1000), .A3(new_n835), .A4(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n284), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n576), .B(new_n356), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n819), .A2(new_n723), .A3(new_n773), .A4(new_n790), .ZN(new_n1008));
  AND4_X1   g822(.A1(new_n744), .A2(new_n803), .A3(new_n805), .A4(new_n893), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n1008), .A2(new_n835), .A3(new_n1009), .ZN(new_n1010));
  OR3_X1    g824(.A1(new_n1010), .A2(G953), .A3(new_n843), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n1006), .B1(G900), .B2(G953), .ZN(new_n1012));
  AOI22_X1  g826(.A1(new_n1007), .A2(KEYINPUT125), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(KEYINPUT126), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n284), .B1(G227), .B2(G900), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1006), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1016), .B1(new_n1004), .B2(new_n284), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT125), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .A4(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1015), .A2(new_n1014), .ZN(new_n1021));
  OR2_X1    g835(.A1(new_n1015), .A2(new_n1014), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1023), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1024));
  AND2_X1   g838(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1025));
  OAI211_X1 g839(.A(new_n1021), .B(new_n1022), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  AND2_X1   g840(.A1(new_n1020), .A2(new_n1026), .ZN(G72));
  NAND2_X1  g841(.A1(G472), .A2(G902), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1028), .B(KEYINPUT63), .Z(new_n1029));
  OR2_X1    g843(.A1(new_n1010), .A2(new_n843), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1029), .B1(new_n1030), .B2(new_n892), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1031), .A2(new_n552), .A3(new_n577), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1029), .B1(new_n1004), .B2(new_n892), .ZN(new_n1033));
  INV_X1    g847(.A(new_n730), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n938), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g849(.A(new_n571), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n577), .A2(new_n553), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1029), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g852(.A(new_n1038), .B(KEYINPUT127), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1039), .B1(new_n907), .B2(new_n911), .ZN(new_n1040));
  AND3_X1   g854(.A1(new_n1032), .A2(new_n1035), .A3(new_n1040), .ZN(G57));
endmodule


