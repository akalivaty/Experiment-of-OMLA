//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n616, new_n617, new_n619,
    new_n620, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT66), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G221), .A3(G218), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  AND3_X1   g033(.A1(KEYINPUT68), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n459));
  AOI21_X1  g034(.A(KEYINPUT3), .B1(KEYINPUT68), .B2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n461), .A2(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G137), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(G101), .A3(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n467), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(new_n464), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(G160));
  NAND2_X1  g045(.A1(new_n462), .A2(G136), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n464), .A2(G112), .ZN(new_n472));
  OAI21_X1  g047(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(G2105), .B1(new_n459), .B2(new_n460), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT69), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n474), .B1(new_n476), .B2(G124), .ZN(G162));
  OAI211_X1 g052(.A(G126), .B(G2105), .C1(new_n459), .C2(new_n460), .ZN(new_n478));
  OR2_X1    g053(.A1(G102), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G114), .C2(new_n464), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n464), .A2(G138), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT70), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT4), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(new_n467), .C1(new_n483), .C2(new_n484), .ZN(new_n486));
  OAI211_X1 g061(.A(G138), .B(new_n464), .C1(new_n459), .C2(new_n460), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n481), .B1(new_n486), .B2(new_n488), .ZN(G164));
  INV_X1    g064(.A(G543), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(KEYINPUT5), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT5), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G543), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n490), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT6), .B(G651), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  XOR2_X1   g074(.A(KEYINPUT72), .B(G88), .Z(new_n500));
  NAND2_X1  g075(.A1(new_n497), .A2(G543), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n499), .A2(new_n500), .B1(G50), .B2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n496), .A2(G62), .ZN(new_n505));
  NAND2_X1  g080(.A1(G75), .A2(G543), .ZN(new_n506));
  XOR2_X1   g081(.A(new_n506), .B(KEYINPUT73), .Z(new_n507));
  AOI21_X1  g082(.A(new_n504), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G166));
  NAND2_X1  g086(.A1(new_n499), .A2(G89), .ZN(new_n512));
  AND3_X1   g087(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT75), .B(G51), .ZN(new_n514));
  OAI221_X1 g089(.A(new_n512), .B1(KEYINPUT7), .B2(new_n513), .C1(new_n501), .C2(new_n514), .ZN(new_n515));
  AOI211_X1 g090(.A(KEYINPUT74), .B(new_n491), .C1(new_n494), .C2(new_n495), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT74), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n494), .A2(new_n495), .ZN(new_n518));
  INV_X1    g093(.A(new_n491), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G63), .ZN(new_n522));
  NAND3_X1  g097(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n504), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n515), .A2(new_n524), .ZN(G168));
  INV_X1    g100(.A(G64), .ZN(new_n526));
  NOR3_X1   g101(.A1(new_n516), .A2(new_n520), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(G77), .A2(G543), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(KEYINPUT76), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n531));
  AND3_X1   g106(.A1(new_n490), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n532));
  AOI21_X1  g107(.A(KEYINPUT71), .B1(new_n490), .B2(KEYINPUT5), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n519), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT74), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n496), .A2(new_n517), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g112(.A(new_n531), .B(new_n528), .C1(new_n537), .C2(new_n526), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n530), .A2(G651), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT77), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT77), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n530), .A2(new_n538), .A3(new_n541), .A4(G651), .ZN(new_n542));
  XNOR2_X1  g117(.A(KEYINPUT78), .B(G52), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n502), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n544), .B1(new_n498), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n540), .A2(new_n542), .A3(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  XOR2_X1   g124(.A(KEYINPUT79), .B(G43), .Z(new_n550));
  NAND2_X1  g125(.A1(new_n502), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n496), .A2(G81), .A3(new_n497), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(G68), .A2(G543), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n556), .B1(new_n521), .B2(G56), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n554), .B1(new_n557), .B2(new_n504), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  OR3_X1    g140(.A1(new_n501), .A2(KEYINPUT80), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT80), .B1(new_n501), .B2(new_n565), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n566), .A2(KEYINPUT9), .A3(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT9), .ZN(new_n569));
  OAI211_X1 g144(.A(KEYINPUT80), .B(new_n569), .C1(new_n501), .C2(new_n565), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n496), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n572));
  INV_X1    g147(.A(G91), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n572), .A2(new_n504), .B1(new_n573), .B2(new_n498), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G299));
  INV_X1    g151(.A(G168), .ZN(G286));
  INV_X1    g152(.A(KEYINPUT81), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n510), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n503), .A2(new_n509), .A3(KEYINPUT81), .ZN(new_n580));
  AND2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(G303));
  AOI22_X1  g156(.A1(new_n499), .A2(G87), .B1(G49), .B2(new_n502), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G288));
  AOI22_X1  g159(.A1(new_n496), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n504), .ZN(new_n586));
  INV_X1    g161(.A(G86), .ZN(new_n587));
  INV_X1    g162(.A(G48), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n498), .A2(new_n587), .B1(new_n588), .B2(new_n501), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n504), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n498), .A2(new_n594), .B1(new_n595), .B2(new_n501), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G290));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OR3_X1    g174(.A1(new_n498), .A2(KEYINPUT82), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(KEYINPUT82), .B1(new_n498), .B2(new_n599), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n602), .B(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n502), .A2(G54), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n496), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(new_n504), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT83), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G171), .B2(new_n609), .ZN(G284));
  OAI21_X1  g186(.A(new_n610), .B1(G171), .B2(new_n609), .ZN(G321));
  NAND2_X1  g187(.A1(G299), .A2(new_n609), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n609), .B2(G168), .ZN(G297));
  OAI21_X1  g189(.A(new_n613), .B1(new_n609), .B2(G168), .ZN(G280));
  INV_X1    g190(.A(G860), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n608), .B1(G559), .B2(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT84), .Z(G148));
  OR2_X1    g193(.A1(new_n608), .A2(G559), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g196(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g197(.A1(new_n476), .A2(G123), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT85), .Z(new_n624));
  NAND2_X1  g199(.A1(new_n462), .A2(G135), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n464), .A2(G111), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n624), .B(new_n625), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n628), .A2(G2096), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(G2096), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n464), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2100), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n629), .A2(new_n630), .A3(new_n634), .ZN(G156));
  XNOR2_X1  g210(.A(G2427), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2430), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  OR2_X1    g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n638), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(KEYINPUT14), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n641), .B(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2443), .B(G2446), .Z(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(G14), .B1(new_n646), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n651), .B1(new_n650), .B2(new_n646), .ZN(G401));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT87), .ZN(new_n654));
  NOR2_X1   g229(.A1(G2072), .A2(G2078), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n442), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n654), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT18), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n654), .A2(new_n656), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n656), .B(KEYINPUT17), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n661), .B(new_n658), .C1(new_n654), .C2(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n662), .A2(new_n654), .A3(new_n657), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n660), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2096), .B(G2100), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT88), .ZN(new_n669));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n671), .A2(KEYINPUT89), .ZN(new_n672));
  XOR2_X1   g247(.A(G1971), .B(G1976), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(KEYINPUT89), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT20), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n669), .A2(new_n670), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n678), .B1(new_n671), .B2(new_n674), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n674), .A2(KEYINPUT90), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT91), .ZN(new_n683));
  XOR2_X1   g258(.A(G1981), .B(G1986), .Z(new_n684));
  XNOR2_X1  g259(.A(G1991), .B(G1996), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n683), .B(new_n688), .ZN(G229));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  AND3_X1   g265(.A1(new_n690), .A2(KEYINPUT92), .A3(G25), .ZN(new_n691));
  AOI21_X1  g266(.A(KEYINPUT92), .B1(new_n690), .B2(G25), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n462), .A2(G131), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n464), .A2(G107), .ZN(new_n694));
  OAI21_X1  g269(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n476), .B2(G119), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT93), .Z(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT94), .Z(new_n699));
  AOI211_X1 g274(.A(new_n691), .B(new_n692), .C1(new_n699), .C2(G29), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT35), .B(G1991), .Z(new_n701));
  OR2_X1    g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(G23), .B(G288), .S(G16), .Z(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT33), .B(G1976), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(KEYINPUT95), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(KEYINPUT95), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G22), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G166), .B2(new_n708), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G1971), .ZN(new_n711));
  NOR2_X1   g286(.A1(G6), .A2(G16), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n590), .B2(G16), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT32), .B(G1981), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n711), .A2(new_n715), .ZN(new_n716));
  AND3_X1   g291(.A1(new_n706), .A2(new_n707), .A3(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT34), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n700), .A2(new_n701), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n708), .A2(G24), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n597), .B2(new_n708), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT36), .ZN(new_n723));
  OAI22_X1  g298(.A1(new_n722), .A2(G1986), .B1(KEYINPUT97), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G1986), .B2(new_n722), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n702), .A2(new_n719), .A3(new_n720), .A4(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n717), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n726), .B1(KEYINPUT34), .B2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT96), .ZN(new_n729));
  OAI21_X1  g304(.A(KEYINPUT97), .B1(new_n729), .B2(new_n723), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n728), .A2(new_n730), .ZN(new_n732));
  NOR2_X1   g307(.A1(G168), .A2(new_n708), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n708), .B2(G21), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G1966), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n735), .A2(KEYINPUT102), .B1(KEYINPUT103), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(KEYINPUT102), .B2(new_n735), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n736), .A2(KEYINPUT103), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n738), .B(new_n739), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n690), .A2(G35), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G162), .B2(new_n690), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT29), .Z(new_n743));
  INV_X1    g318(.A(G2090), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n708), .A2(G20), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT23), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n575), .B2(new_n708), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G1956), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT105), .ZN(new_n751));
  NOR2_X1   g326(.A1(G4), .A2(G16), .ZN(new_n752));
  INV_X1    g327(.A(new_n608), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(G16), .ZN(new_n754));
  INV_X1    g329(.A(G1348), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n708), .A2(G19), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n559), .B2(new_n708), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT98), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G1341), .ZN(new_n760));
  INV_X1    g335(.A(G34), .ZN(new_n761));
  OR2_X1    g336(.A1(new_n761), .A2(KEYINPUT24), .ZN(new_n762));
  AOI21_X1  g337(.A(G29), .B1(new_n761), .B2(KEYINPUT24), .ZN(new_n763));
  AOI22_X1  g338(.A1(G160), .A2(G29), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(G2084), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT101), .Z(new_n766));
  AND2_X1   g341(.A1(new_n690), .A2(G33), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n462), .A2(G139), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT25), .Z(new_n770));
  AOI22_X1  g345(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n771));
  OAI211_X1 g346(.A(new_n768), .B(new_n770), .C1(new_n464), .C2(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n767), .B1(new_n772), .B2(G29), .ZN(new_n773));
  INV_X1    g348(.A(G2072), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT31), .B(G11), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT30), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n777), .A2(G28), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n690), .B1(new_n777), .B2(G28), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n775), .B(new_n776), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n764), .A2(G2084), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n773), .A2(new_n774), .ZN(new_n782));
  OR4_X1    g357(.A1(new_n766), .A2(new_n780), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n628), .A2(new_n690), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT104), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n743), .A2(new_n744), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n690), .A2(G26), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT28), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n462), .A2(G140), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT99), .Z(new_n790));
  OR2_X1    g365(.A1(G104), .A2(G2105), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n791), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT100), .Z(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(new_n476), .B2(G128), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n788), .B1(new_n795), .B2(G29), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G2067), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n690), .A2(G32), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n462), .A2(G141), .ZN(new_n799));
  NAND3_X1  g374(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT26), .Z(new_n801));
  NAND3_X1  g376(.A1(new_n464), .A2(G105), .A3(G2104), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n799), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G129), .B2(new_n476), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n798), .B1(new_n804), .B2(new_n690), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT27), .B(G1996), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n690), .A2(G27), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(G164), .B2(new_n690), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(G2078), .Z(new_n810));
  NAND4_X1  g385(.A1(new_n786), .A2(new_n797), .A3(new_n807), .A4(new_n810), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n783), .A2(new_n785), .A3(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n751), .A2(new_n756), .A3(new_n760), .A4(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(G171), .A2(new_n708), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G5), .B2(new_n708), .ZN(new_n815));
  INV_X1    g390(.A(G1961), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AND2_X1   g392(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  NOR4_X1   g393(.A1(new_n740), .A2(new_n813), .A3(new_n817), .A4(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n731), .A2(new_n732), .A3(new_n819), .ZN(G150));
  INV_X1    g395(.A(G150), .ZN(G311));
  NAND2_X1  g396(.A1(G80), .A2(G543), .ZN(new_n822));
  INV_X1    g397(.A(G67), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n537), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n496), .A2(G93), .A3(new_n497), .ZN(new_n825));
  INV_X1    g400(.A(G55), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(new_n501), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT106), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n825), .B(KEYINPUT106), .C1(new_n826), .C2(new_n501), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n824), .A2(G651), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(new_n616), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT110), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT109), .B(KEYINPUT37), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n753), .A2(G559), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT38), .Z(new_n837));
  OAI211_X1 g412(.A(KEYINPUT107), .B(new_n554), .C1(new_n557), .C2(new_n504), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(new_n831), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT108), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT107), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n840), .B1(new_n558), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n535), .A2(G56), .A3(new_n536), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n504), .B1(new_n843), .B2(new_n555), .ZN(new_n844));
  OAI211_X1 g419(.A(new_n841), .B(new_n840), .C1(new_n844), .C2(new_n553), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n839), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n841), .B1(new_n844), .B2(new_n553), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT108), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n849), .A2(new_n831), .A3(new_n838), .A4(new_n845), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n837), .B(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n853), .A2(KEYINPUT39), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n616), .B1(new_n853), .B2(KEYINPUT39), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n835), .B1(new_n854), .B2(new_n855), .ZN(G145));
  INV_X1    g431(.A(KEYINPUT111), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n481), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n478), .A2(new_n480), .A3(KEYINPUT111), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n486), .A2(new_n488), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n795), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n698), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n462), .A2(G142), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n464), .A2(G118), .ZN(new_n866));
  OAI21_X1  g441(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(new_n476), .B2(G130), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(new_n632), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n804), .B(new_n772), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n864), .B(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(G162), .B(G160), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n628), .B(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(G37), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n873), .A2(new_n875), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(KEYINPUT40), .Z(G395));
  OR2_X1    g456(.A1(new_n831), .A2(G868), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n597), .B(G305), .ZN(new_n883));
  XNOR2_X1  g458(.A(G166), .B(G288), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(new_n884), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(KEYINPUT114), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n885), .A2(KEYINPUT113), .A3(new_n887), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT113), .B1(new_n885), .B2(new_n887), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n889), .B1(new_n893), .B2(new_n886), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n619), .B(new_n851), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n575), .B1(new_n603), .B2(new_n607), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT41), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n603), .A2(new_n575), .A3(new_n607), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n899), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n901), .A2(new_n896), .ZN(new_n902));
  XNOR2_X1  g477(.A(KEYINPUT112), .B(KEYINPUT41), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n895), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n902), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n905), .B1(new_n906), .B2(new_n895), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n894), .B(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n882), .B1(new_n908), .B2(new_n609), .ZN(G295));
  OAI21_X1  g484(.A(new_n882), .B1(new_n908), .B2(new_n609), .ZN(G331));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n912));
  AND4_X1   g487(.A1(G168), .A2(new_n540), .A3(new_n542), .A4(new_n547), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n546), .B1(new_n539), .B2(KEYINPUT77), .ZN(new_n914));
  AOI21_X1  g489(.A(G168), .B1(new_n914), .B2(new_n542), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n850), .B(new_n847), .C1(new_n913), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(G301), .A2(G286), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n914), .A2(G168), .A3(new_n542), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n851), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n916), .A2(new_n919), .A3(KEYINPUT115), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n918), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT115), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n921), .A2(new_n922), .A3(new_n850), .A4(new_n847), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n920), .A2(new_n904), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT116), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT116), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n920), .A2(new_n904), .A3(new_n923), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n916), .A2(new_n919), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n902), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n925), .A2(new_n892), .A3(new_n927), .A4(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n925), .A2(new_n927), .A3(new_n930), .ZN(new_n933));
  AOI21_X1  g508(.A(G37), .B1(new_n933), .B2(new_n893), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT117), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n932), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n924), .A2(KEYINPUT116), .B1(new_n902), .B2(new_n929), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n892), .B1(new_n937), .B2(new_n927), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT117), .B1(new_n938), .B2(G37), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n912), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n906), .A2(new_n898), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n928), .B(new_n941), .C1(new_n906), .C2(new_n903), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n906), .B1(new_n920), .B2(new_n923), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n942), .B1(new_n943), .B2(KEYINPUT118), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT118), .ZN(new_n945));
  AOI211_X1 g520(.A(new_n945), .B(new_n906), .C1(new_n920), .C2(new_n923), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n893), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n947), .A2(new_n912), .A3(new_n877), .A4(new_n931), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT119), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n931), .A2(new_n877), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n951), .A2(KEYINPUT119), .A3(new_n912), .A4(new_n947), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n911), .B1(new_n940), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT43), .B1(new_n936), .B2(new_n939), .ZN(new_n955));
  AND3_X1   g530(.A1(new_n951), .A2(KEYINPUT43), .A3(new_n947), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT44), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n954), .A2(new_n957), .ZN(G397));
  AOI21_X1  g533(.A(G1384), .B1(new_n860), .B2(new_n861), .ZN(new_n959));
  OR2_X1    g534(.A1(new_n959), .A2(KEYINPUT45), .ZN(new_n960));
  INV_X1    g535(.A(new_n469), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n961), .A2(new_n463), .A3(G40), .A4(new_n465), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G2067), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n795), .B(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n964), .B1(new_n966), .B2(new_n804), .ZN(new_n967));
  OR3_X1    g542(.A1(new_n964), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT46), .B1(new_n964), .B2(G1996), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT47), .ZN(new_n971));
  INV_X1    g546(.A(new_n701), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n698), .B(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n963), .ZN(new_n974));
  INV_X1    g549(.A(new_n966), .ZN(new_n975));
  XOR2_X1   g550(.A(new_n804), .B(G1996), .Z(new_n976));
  OAI21_X1  g551(.A(new_n963), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(G290), .A2(G1986), .ZN(new_n979));
  XOR2_X1   g554(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(new_n963), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n980), .ZN(new_n982));
  INV_X1    g557(.A(new_n979), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n982), .B1(new_n983), .B2(new_n964), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n978), .A2(new_n981), .A3(new_n984), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n699), .A2(new_n972), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(new_n977), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n987), .B1(G2067), .B2(new_n795), .ZN(new_n988));
  AOI211_X1 g563(.A(new_n971), .B(new_n985), .C1(new_n963), .C2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G40), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n466), .A2(new_n990), .A3(new_n469), .ZN(new_n991));
  NOR2_X1   g566(.A1(G164), .A2(G1384), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n991), .B1(new_n992), .B2(KEYINPUT45), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n994), .A2(G1384), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n862), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(KEYINPUT120), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT120), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n862), .A2(new_n998), .A3(new_n995), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n993), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(G1971), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1002), .A2(new_n991), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n959), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(G2090), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT121), .B1(new_n1001), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n579), .A2(G8), .A3(new_n580), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT55), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT121), .ZN(new_n1012));
  OAI221_X1 g587(.A(new_n1012), .B1(new_n1006), .B2(G2090), .C1(new_n1000), .C2(G1971), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1008), .A2(new_n1011), .A3(new_n1013), .A4(G8), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT122), .ZN(new_n1015));
  INV_X1    g590(.A(G8), .ZN(new_n1016));
  INV_X1    g591(.A(new_n992), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n962), .B1(new_n1017), .B2(new_n994), .ZN(new_n1018));
  INV_X1    g593(.A(new_n999), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n998), .B1(new_n862), .B2(new_n995), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1971), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1021), .A2(new_n1022), .B1(new_n1023), .B2(new_n744), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1016), .B1(new_n1024), .B2(new_n1012), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT122), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1025), .A2(new_n1026), .A3(new_n1011), .A4(new_n1008), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1015), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n995), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n960), .B(new_n991), .C1(G164), .C2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n736), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(G2084), .B2(new_n1006), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT123), .B(G8), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(G305), .A2(G1981), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT49), .ZN(new_n1037));
  INV_X1    g612(.A(G1981), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n590), .A2(new_n1038), .ZN(new_n1039));
  OR3_X1    g614(.A1(new_n1036), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n959), .A2(new_n991), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n1034), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1037), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1040), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(G1976), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT52), .B1(G288), .B2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1043), .B(new_n1047), .C1(new_n1046), .C2(G288), .ZN(new_n1048));
  NOR2_X1   g623(.A1(G288), .A2(new_n1046), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT52), .B1(new_n1042), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1045), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT63), .ZN(new_n1052));
  NOR4_X1   g627(.A1(new_n1035), .A2(new_n1051), .A3(new_n1052), .A4(G286), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1025), .A2(new_n1008), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1028), .B(new_n1053), .C1(new_n1011), .C2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1051), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n991), .B1(new_n1017), .B2(KEYINPUT50), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n959), .A2(new_n1004), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1057), .A2(new_n1058), .A3(G2090), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1034), .B1(new_n1001), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n1010), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1056), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1035), .A2(G286), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1028), .A2(KEYINPUT124), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n1052), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1062), .B1(new_n1015), .B2(new_n1027), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT124), .B1(new_n1067), .B2(new_n1064), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1055), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT125), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1028), .A2(new_n1051), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1045), .A2(new_n1046), .A3(new_n583), .A4(new_n582), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(G1981), .B2(G305), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1071), .B1(new_n1043), .B2(new_n1073), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1069), .A2(new_n1070), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1070), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1067), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1032), .A2(G8), .ZN(new_n1078));
  NOR2_X1   g653(.A1(G168), .A2(new_n1033), .ZN(new_n1079));
  OAI221_X1 g654(.A(KEYINPUT51), .B1(new_n1078), .B2(new_n1079), .C1(new_n1035), .C2(G168), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1079), .A2(KEYINPUT51), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1035), .A2(new_n1081), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  XOR2_X1   g658(.A(G301), .B(KEYINPUT54), .Z(new_n1084));
  OR2_X1    g659(.A1(new_n1021), .A2(G2078), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n1086));
  AOI22_X1  g661(.A1(new_n1085), .A2(new_n1086), .B1(new_n816), .B2(new_n1006), .ZN(new_n1087));
  AOI211_X1 g662(.A(new_n1086), .B(G2078), .C1(new_n997), .C2(new_n999), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1088), .A2(new_n991), .A3(new_n960), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1084), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  OR3_X1    g665(.A1(new_n1030), .A2(new_n1086), .A3(G2078), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1087), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1090), .B1(new_n1092), .B2(new_n1084), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n575), .B(KEYINPUT57), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT56), .B(G2072), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1000), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(G1956), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1094), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1096), .A2(new_n1094), .A3(new_n1098), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1100), .A2(new_n1101), .A3(KEYINPUT126), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT126), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT61), .B1(new_n1099), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1041), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1006), .A2(new_n755), .B1(new_n1106), .B2(new_n965), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1107), .A2(KEYINPUT60), .A3(new_n608), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n608), .B1(new_n1107), .B2(KEYINPUT60), .ZN(new_n1109));
  OAI22_X1  g684(.A1(new_n1108), .A2(new_n1109), .B1(KEYINPUT60), .B2(new_n1107), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1100), .A2(new_n1101), .A3(KEYINPUT61), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT58), .B(G1341), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n1021), .A2(G1996), .B1(new_n1106), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(new_n559), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT59), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(new_n1116), .A3(new_n559), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1105), .A2(new_n1110), .A3(new_n1111), .A4(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1107), .A2(new_n608), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1099), .B1(new_n1120), .B2(new_n1101), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1093), .B1(new_n1119), .B2(new_n1121), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n1092), .A2(KEYINPUT62), .A3(G301), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1083), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1092), .A2(G301), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(KEYINPUT62), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1077), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1075), .A2(new_n1076), .A3(new_n1128), .ZN(new_n1129));
  AND2_X1   g704(.A1(G290), .A2(G1986), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n963), .B1(new_n1130), .B2(new_n979), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n978), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n989), .B1(new_n1129), .B2(new_n1132), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g708(.A1(new_n940), .A2(new_n953), .ZN(new_n1135));
  INV_X1    g709(.A(new_n880), .ZN(new_n1136));
  INV_X1    g710(.A(G319), .ZN(new_n1137));
  NOR4_X1   g711(.A1(G229), .A2(new_n1137), .A3(G401), .A4(G227), .ZN(new_n1138));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g713(.A1(new_n1135), .A2(new_n1139), .ZN(G308));
  OAI211_X1 g714(.A(new_n1136), .B(new_n1138), .C1(new_n940), .C2(new_n953), .ZN(G225));
endmodule


