//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939;
  INV_X1    g000(.A(KEYINPUT32), .ZN(new_n187));
  INV_X1    g001(.A(G472), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT31), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G143), .ZN(new_n194));
  OAI21_X1  g008(.A(G128), .B1(new_n192), .B2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(G146), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n197), .A3(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n195), .A2(KEYINPUT0), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n196), .A2(new_n197), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT0), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G128), .ZN(new_n203));
  AND2_X1   g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT11), .ZN(new_n205));
  INV_X1    g019(.A(G134), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(G137), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(G137), .ZN(new_n208));
  INV_X1    g022(.A(G137), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT11), .A3(G134), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G131), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n207), .A2(new_n210), .A3(new_n213), .A4(new_n208), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT65), .B1(new_n206), .B2(G137), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(new_n209), .A3(G134), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n216), .A2(new_n218), .A3(new_n208), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G131), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n220), .A2(new_n214), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT66), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(G143), .B(G146), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n198), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n199), .ZN(new_n229));
  OAI22_X1  g043(.A1(new_n228), .A2(new_n229), .B1(new_n197), .B2(new_n226), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n204), .A2(new_n215), .B1(new_n221), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(G116), .B(G119), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n232), .A2(KEYINPUT67), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT2), .B(G113), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n233), .B(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(KEYINPUT69), .B(G237), .ZN(new_n238));
  INV_X1    g052(.A(G953), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(G210), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT26), .B(G101), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n237), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT30), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n248), .B1(new_n231), .B2(KEYINPUT64), .ZN(new_n249));
  INV_X1    g063(.A(new_n215), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n200), .A2(new_n203), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n226), .A2(new_n197), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n253));
  OAI21_X1  g067(.A(G128), .B1(new_n201), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n252), .B1(new_n254), .B2(new_n199), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n220), .A2(new_n214), .ZN(new_n256));
  OAI22_X1  g070(.A1(new_n250), .A2(new_n251), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT64), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT30), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n249), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n236), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n247), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AOI211_X1 g076(.A(KEYINPUT68), .B(new_n236), .C1(new_n249), .C2(new_n259), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n246), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n221), .A2(new_n230), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n215), .A2(new_n203), .A3(new_n200), .ZN(new_n268));
  AOI211_X1 g082(.A(KEYINPUT64), .B(new_n248), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT30), .B1(new_n257), .B2(new_n258), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n261), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT68), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n247), .B(new_n261), .C1(new_n269), .C2(new_n270), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n245), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT71), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n190), .B1(new_n266), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT28), .B1(new_n231), .B2(new_n236), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n257), .A2(new_n261), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n237), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n277), .B1(new_n279), .B2(KEYINPUT28), .ZN(new_n280));
  OAI22_X1  g094(.A1(new_n264), .A2(KEYINPUT31), .B1(new_n280), .B2(new_n244), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n188), .B(new_n189), .C1(new_n276), .C2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n272), .A2(new_n273), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT71), .B1(new_n285), .B2(new_n246), .ZN(new_n286));
  AOI211_X1 g100(.A(new_n265), .B(new_n245), .C1(new_n272), .C2(new_n273), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT31), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n280), .A2(new_n244), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n289), .B1(new_n274), .B2(new_n190), .ZN(new_n290));
  AOI21_X1  g104(.A(G902), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT72), .B1(new_n291), .B2(new_n188), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n187), .B1(new_n284), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n282), .A2(new_n187), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n285), .A2(new_n237), .ZN(new_n296));
  INV_X1    g110(.A(new_n244), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT29), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n280), .A2(new_n244), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n301), .B(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n189), .B1(new_n300), .B2(new_n299), .ZN(new_n304));
  OAI21_X1  g118(.A(G472), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n293), .A2(new_n295), .A3(new_n305), .ZN(new_n306));
  OR2_X1    g120(.A1(KEYINPUT76), .A2(G140), .ZN(new_n307));
  NAND2_X1  g121(.A1(KEYINPUT76), .A2(G140), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(G125), .A3(new_n308), .ZN(new_n309));
  AND2_X1   g123(.A1(KEYINPUT77), .A2(G125), .ZN(new_n310));
  NOR2_X1   g124(.A1(KEYINPUT77), .A2(G125), .ZN(new_n311));
  OAI21_X1  g125(.A(G140), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n312), .A3(KEYINPUT16), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT78), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT78), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n309), .A2(new_n312), .A3(new_n315), .A4(KEYINPUT16), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n310), .A2(new_n311), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT16), .ZN(new_n319));
  INV_X1    g133(.A(G140), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n317), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n193), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT79), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n317), .A2(G146), .A3(new_n321), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n198), .A2(G119), .ZN(new_n327));
  INV_X1    g141(.A(G119), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G128), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT23), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n328), .A2(KEYINPUT23), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n330), .B1(G128), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  OR2_X1    g147(.A1(new_n333), .A2(KEYINPUT75), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(KEYINPUT75), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n334), .A2(G110), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT74), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n329), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n328), .A2(KEYINPUT74), .A3(G128), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n338), .A2(new_n339), .B1(G119), .B2(new_n198), .ZN(new_n340));
  XOR2_X1   g154(.A(KEYINPUT24), .B(G110), .Z(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n317), .A2(KEYINPUT79), .A3(G146), .A4(new_n321), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n326), .A2(new_n336), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  OAI22_X1  g158(.A1(new_n333), .A2(G110), .B1(new_n340), .B2(new_n341), .ZN(new_n345));
  OR2_X1    g159(.A1(G125), .A2(G140), .ZN(new_n346));
  NAND2_X1  g160(.A1(G125), .A2(G140), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n346), .A2(KEYINPUT80), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(KEYINPUT80), .B1(new_n346), .B2(new_n347), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n193), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n325), .A2(new_n345), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n344), .A2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(KEYINPUT81), .B(KEYINPUT22), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n353), .B(G137), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n239), .A2(G221), .A3(G234), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n354), .B(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n356), .B(KEYINPUT82), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT83), .B1(new_n352), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n344), .A2(new_n351), .A3(new_n356), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n352), .A2(KEYINPUT83), .A3(new_n357), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT25), .B1(new_n362), .B2(G902), .ZN(new_n363));
  INV_X1    g177(.A(G217), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(G234), .B2(new_n189), .ZN(new_n365));
  INV_X1    g179(.A(new_n361), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n366), .A2(new_n358), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT25), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n367), .A2(new_n368), .A3(new_n189), .A4(new_n360), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n363), .A2(new_n365), .A3(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n367), .A2(KEYINPUT84), .A3(new_n360), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT84), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n362), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n365), .A2(G902), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n371), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(G110), .B(G140), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n239), .A2(G227), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G104), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT3), .B1(new_n381), .B2(G107), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT3), .ZN(new_n383));
  INV_X1    g197(.A(G107), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(new_n384), .A3(G104), .ZN(new_n385));
  INV_X1    g199(.A(G101), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n381), .A2(G107), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n382), .A2(new_n385), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT85), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n388), .B(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n384), .A2(G104), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n386), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT86), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n392), .B(new_n393), .ZN(new_n394));
  OAI22_X1  g208(.A1(new_n228), .A2(new_n229), .B1(new_n222), .B2(new_n197), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n390), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT87), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT10), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n397), .B1(new_n396), .B2(new_n398), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n382), .A2(new_n385), .A3(new_n387), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G101), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n390), .A2(KEYINPUT4), .A3(new_n403), .ZN(new_n404));
  OR2_X1    g218(.A1(new_n403), .A2(KEYINPUT4), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(new_n204), .A3(new_n405), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n390), .A2(KEYINPUT10), .A3(new_n230), .A4(new_n394), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n250), .B1(new_n401), .B2(new_n409), .ZN(new_n410));
  NOR4_X1   g224(.A1(new_n408), .A2(new_n399), .A3(new_n400), .A4(new_n215), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n380), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT88), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n396), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n230), .B1(new_n390), .B2(new_n394), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(new_n250), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(KEYINPUT12), .ZN(new_n419));
  INV_X1    g233(.A(new_n411), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(new_n420), .A3(new_n379), .ZN(new_n421));
  OAI211_X1 g235(.A(KEYINPUT88), .B(new_n380), .C1(new_n410), .C2(new_n411), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n414), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G469), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(new_n189), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n419), .A2(new_n420), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n380), .ZN(new_n427));
  OR3_X1    g241(.A1(new_n410), .A2(new_n411), .A3(new_n380), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(new_n428), .A3(G469), .ZN(new_n429));
  NAND2_X1  g243(.A1(G469), .A2(G902), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n425), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  XOR2_X1   g245(.A(KEYINPUT9), .B(G234), .Z(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(G221), .B1(new_n433), .B2(G902), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n230), .A2(new_n318), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT91), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT91), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n438), .B1(new_n251), .B2(new_n318), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n437), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G224), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT7), .B1(new_n441), .B2(G953), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G116), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n444), .A2(KEYINPUT5), .A3(G119), .ZN(new_n445));
  INV_X1    g259(.A(G113), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n232), .A2(KEYINPUT5), .ZN(new_n448));
  AOI22_X1  g262(.A1(new_n447), .A2(new_n448), .B1(new_n235), .B2(new_n232), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n390), .A2(new_n449), .A3(new_n394), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n404), .A2(new_n261), .A3(new_n405), .ZN(new_n452));
  XNOR2_X1  g266(.A(G110), .B(G122), .ZN(new_n453));
  XOR2_X1   g267(.A(new_n453), .B(KEYINPUT90), .Z(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  XOR2_X1   g269(.A(KEYINPUT92), .B(KEYINPUT8), .Z(new_n456));
  XNOR2_X1  g270(.A(new_n454), .B(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n449), .B1(new_n390), .B2(new_n394), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n457), .B1(new_n450), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n442), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n437), .B(new_n460), .C1(new_n436), .C2(new_n439), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n443), .A2(new_n455), .A3(new_n459), .A4(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n189), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT93), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n451), .A2(new_n452), .ZN(new_n465));
  INV_X1    g279(.A(new_n454), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(KEYINPUT6), .A3(new_n455), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n441), .A2(G953), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n440), .B(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT6), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n465), .A2(new_n471), .A3(new_n466), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n468), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT93), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n462), .A2(new_n474), .A3(new_n189), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n464), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(G210), .B1(G237), .B2(G902), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n464), .A2(new_n473), .A3(new_n477), .A4(new_n475), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(G214), .B1(G237), .B2(G902), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n482), .B(KEYINPUT89), .ZN(new_n483));
  NAND2_X1  g297(.A1(G234), .A2(G237), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(G952), .A3(new_n239), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(KEYINPUT100), .ZN(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  XOR2_X1   g301(.A(KEYINPUT21), .B(G898), .Z(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n484), .A2(G902), .A3(G953), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n487), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n481), .A2(new_n483), .A3(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(G128), .B(G143), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(new_n206), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n444), .A2(KEYINPUT14), .A3(G122), .ZN(new_n497));
  XNOR2_X1  g311(.A(G116), .B(G122), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  OAI211_X1 g313(.A(G107), .B(new_n497), .C1(new_n499), .C2(KEYINPUT14), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n496), .B(new_n500), .C1(G107), .C2(new_n499), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n495), .A2(KEYINPUT13), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n191), .A2(G128), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n502), .B(G134), .C1(KEYINPUT13), .C2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n498), .B(new_n384), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n495), .A2(new_n206), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n432), .A2(G217), .A3(new_n239), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n510), .A2(new_n189), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT15), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n512), .A2(KEYINPUT99), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n512), .A2(KEYINPUT99), .ZN(new_n514));
  OAI21_X1  g328(.A(G478), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n511), .B(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT98), .ZN(new_n517));
  XNOR2_X1  g331(.A(G113), .B(G122), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(new_n381), .ZN(new_n519));
  AND2_X1   g333(.A1(KEYINPUT69), .A2(G237), .ZN(new_n520));
  NOR2_X1   g334(.A1(KEYINPUT69), .A2(G237), .ZN(new_n521));
  OAI211_X1 g335(.A(G214), .B(new_n239), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n191), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n238), .A2(G143), .A3(G214), .A4(new_n239), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(KEYINPUT18), .A3(G131), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT94), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n523), .A2(new_n524), .ZN(new_n528));
  NAND2_X1  g342(.A1(KEYINPUT18), .A2(G131), .ZN(new_n529));
  XOR2_X1   g343(.A(new_n529), .B(KEYINPUT95), .Z(new_n530));
  NAND2_X1  g344(.A1(new_n309), .A2(new_n312), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(G146), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n528), .A2(new_n530), .B1(new_n350), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT94), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n525), .A2(new_n534), .A3(KEYINPUT18), .A4(G131), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n527), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n326), .A2(new_n343), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n525), .A2(G131), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n523), .A2(new_n524), .A3(new_n213), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  MUX2_X1   g355(.A(new_n541), .B(new_n539), .S(KEYINPUT17), .Z(new_n542));
  AOI21_X1  g356(.A(new_n537), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT19), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(new_n348), .B2(new_n349), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT96), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n531), .A2(KEYINPUT19), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT96), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n548), .B(new_n544), .C1(new_n348), .C2(new_n349), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n546), .A2(new_n193), .A3(new_n547), .A4(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n325), .A2(new_n550), .A3(new_n541), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n536), .ZN(new_n552));
  INV_X1    g366(.A(new_n519), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT97), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n552), .A2(KEYINPUT97), .A3(new_n553), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n519), .A2(new_n543), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(G475), .A2(G902), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n517), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n556), .A2(new_n557), .ZN(new_n562));
  AOI211_X1 g376(.A(new_n553), .B(new_n537), .C1(new_n538), .C2(new_n542), .ZN(new_n563));
  OAI211_X1 g377(.A(KEYINPUT98), .B(new_n559), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n561), .A2(new_n564), .A3(KEYINPUT20), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n543), .A2(new_n519), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n189), .B1(new_n566), .B2(new_n563), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G475), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT20), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n517), .B(new_n569), .C1(new_n558), .C2(new_n560), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n565), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  NOR4_X1   g385(.A1(new_n435), .A2(new_n494), .A3(new_n516), .A4(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n306), .A2(new_n376), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n573), .B(G101), .ZN(G3));
  OAI21_X1  g388(.A(KEYINPUT101), .B1(new_n291), .B2(new_n188), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT101), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n266), .A2(new_n275), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n281), .B1(new_n577), .B2(KEYINPUT31), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n576), .B(G472), .C1(new_n578), .C2(G902), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n282), .A2(new_n283), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n291), .A2(KEYINPUT72), .A3(new_n188), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AND3_X1   g397(.A1(new_n580), .A2(new_n376), .A3(new_n583), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n431), .A2(new_n434), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G478), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(new_n189), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n511), .A2(new_n587), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT102), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n591), .B1(new_n508), .B2(new_n592), .ZN(new_n593));
  XOR2_X1   g407(.A(new_n510), .B(new_n593), .Z(new_n594));
  AOI211_X1 g408(.A(new_n588), .B(new_n590), .C1(new_n594), .C2(G478), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n571), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n481), .ZN(new_n598));
  INV_X1    g412(.A(new_n482), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n598), .A2(new_n599), .A3(new_n492), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n586), .A2(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT34), .B(G104), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(KEYINPUT103), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n602), .B(new_n604), .ZN(G6));
  INV_X1    g419(.A(new_n516), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n571), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n584), .A2(new_n585), .A3(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT35), .B(G107), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G9));
  NOR2_X1   g425(.A1(new_n357), .A2(KEYINPUT36), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n352), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n374), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n370), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n572), .A2(new_n583), .A3(new_n580), .A4(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT104), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT37), .B(G110), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G12));
  INV_X1    g433(.A(G900), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n487), .B1(new_n620), .B2(new_n491), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n571), .A2(new_n606), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n599), .B1(new_n479), .B2(new_n480), .ZN(new_n623));
  AND3_X1   g437(.A1(new_n585), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n306), .A2(new_n624), .A3(new_n615), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G128), .ZN(G30));
  AOI22_X1  g440(.A1(new_n266), .A2(new_n275), .B1(new_n297), .B2(new_n279), .ZN(new_n627));
  OAI21_X1  g441(.A(G472), .B1(new_n627), .B2(G902), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n293), .A2(new_n295), .A3(new_n628), .ZN(new_n629));
  AND4_X1   g443(.A1(new_n482), .A2(new_n629), .A3(new_n516), .A4(new_n571), .ZN(new_n630));
  INV_X1    g444(.A(new_n615), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n481), .A2(KEYINPUT105), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT105), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n479), .B2(new_n480), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n635), .A2(KEYINPUT38), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n635), .A2(KEYINPUT38), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n630), .A2(new_n631), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT106), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n621), .B(KEYINPUT39), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n585), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT40), .ZN(new_n645));
  OR3_X1    g459(.A1(new_n640), .A2(new_n641), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n641), .B1(new_n640), .B2(new_n645), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(new_n191), .ZN(G45));
  NOR3_X1   g463(.A1(new_n435), .A2(new_n599), .A3(new_n598), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n596), .A2(new_n621), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n306), .A2(new_n615), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G146), .ZN(G48));
  NAND2_X1  g467(.A1(new_n370), .A2(new_n375), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n294), .B1(new_n583), .B2(new_n187), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n654), .B1(new_n655), .B2(new_n305), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n423), .A2(new_n189), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(G469), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n658), .A2(new_n425), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n434), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n601), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT41), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G113), .ZN(G15));
  INV_X1    g478(.A(new_n660), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n665), .A2(new_n608), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n656), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G116), .ZN(G18));
  AOI21_X1  g482(.A(new_n631), .B1(new_n655), .B2(new_n305), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n565), .A2(new_n568), .A3(new_n570), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(new_n493), .A3(new_n606), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n658), .A2(new_n623), .A3(new_n434), .A4(new_n425), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(KEYINPUT107), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n672), .A2(KEYINPUT107), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n671), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n669), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G119), .ZN(G21));
  XNOR2_X1  g492(.A(new_n291), .B(new_n188), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(new_n654), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n571), .A2(new_n516), .A3(new_n623), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(KEYINPUT108), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT108), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n571), .A2(new_n623), .A3(new_n683), .A4(new_n516), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n660), .A2(new_n492), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G122), .ZN(G24));
  NOR2_X1   g503(.A1(new_n631), .A2(new_n679), .ZN(new_n690));
  INV_X1    g504(.A(new_n675), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n690), .B(new_n651), .C1(new_n691), .C2(new_n673), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G125), .ZN(G27));
  NAND3_X1  g507(.A1(new_n479), .A2(new_n482), .A3(new_n480), .ZN(new_n694));
  OR2_X1    g508(.A1(new_n694), .A2(KEYINPUT109), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(KEYINPUT109), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n697), .A2(new_n435), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n306), .A2(new_n376), .A3(new_n651), .A4(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT42), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT111), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n282), .A2(new_n702), .A3(new_n187), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n702), .B1(new_n282), .B2(new_n187), .ZN(new_n705));
  OAI211_X1 g519(.A(KEYINPUT110), .B(new_n295), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n282), .A2(new_n187), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT111), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n708), .B(new_n703), .C1(new_n709), .C2(new_n294), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n706), .A2(new_n710), .A3(new_n305), .ZN(new_n711));
  INV_X1    g525(.A(new_n651), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n712), .A2(new_n435), .A3(new_n697), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n711), .A2(new_n713), .A3(KEYINPUT42), .A4(new_n376), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n701), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT112), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G131), .ZN(G33));
  AND3_X1   g531(.A1(new_n656), .A2(new_n622), .A3(new_n698), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(new_n206), .ZN(G36));
  NAND2_X1  g533(.A1(new_n670), .A2(new_n595), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n670), .A2(KEYINPUT43), .A3(new_n595), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n580), .A2(new_n583), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n724), .A2(new_n725), .A3(new_n615), .ZN(new_n726));
  OR2_X1    g540(.A1(new_n726), .A2(KEYINPUT44), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n427), .A2(new_n428), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(KEYINPUT45), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(G469), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(KEYINPUT46), .A3(new_n430), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT46), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n732), .B(G469), .C1(new_n729), .C2(G902), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n731), .A2(new_n425), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n434), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n642), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n726), .A2(KEYINPUT44), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n697), .B(KEYINPUT113), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n727), .A2(new_n736), .A3(new_n737), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G137), .ZN(G39));
  XOR2_X1   g554(.A(new_n735), .B(KEYINPUT47), .Z(new_n741));
  NOR2_X1   g555(.A1(new_n697), .A2(new_n376), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n306), .A2(new_n712), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G140), .ZN(G42));
  INV_X1    g559(.A(new_n494), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n516), .B(KEYINPUT114), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n596), .B1(new_n571), .B2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n584), .A2(new_n746), .A3(new_n585), .A4(new_n748), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n749), .A2(new_n573), .A3(new_n616), .ZN(new_n750));
  INV_X1    g564(.A(new_n621), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n565), .A2(new_n568), .A3(new_n570), .A4(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n747), .ZN(new_n753));
  OR3_X1    g567(.A1(new_n752), .A2(new_n753), .A3(KEYINPUT115), .ZN(new_n754));
  OAI21_X1  g568(.A(KEYINPUT115), .B1(new_n752), .B2(new_n753), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n756), .B1(new_n655), .B2(new_n305), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n712), .A2(new_n679), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n615), .B(new_n698), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  AOI22_X1  g573(.A1(new_n656), .A2(new_n666), .B1(new_n686), .B2(new_n687), .ZN(new_n760));
  AOI22_X1  g574(.A1(new_n669), .A2(new_n676), .B1(new_n656), .B2(new_n661), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n750), .A2(new_n759), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n718), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n715), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n652), .A2(new_n625), .A3(new_n692), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n431), .A2(new_n370), .A3(new_n434), .A4(new_n614), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n767), .B1(new_n682), .B2(new_n684), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n629), .A2(new_n751), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT116), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n629), .A2(new_n768), .A3(new_n771), .A4(new_n751), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n766), .A2(KEYINPUT52), .A3(new_n770), .A4(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n770), .A2(new_n772), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n652), .A2(new_n625), .A3(new_n692), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n765), .A2(new_n778), .A3(KEYINPUT53), .ZN(new_n779));
  AOI21_X1  g593(.A(KEYINPUT53), .B1(new_n765), .B2(new_n778), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n621), .B1(new_n655), .B2(new_n628), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n771), .B1(new_n784), .B2(new_n768), .ZN(new_n785));
  AND4_X1   g599(.A1(new_n771), .A2(new_n629), .A3(new_n751), .A4(new_n768), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT52), .B1(new_n787), .B2(new_n766), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n775), .A2(new_n774), .A3(new_n776), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n718), .B1(new_n701), .B2(new_n714), .ZN(new_n791));
  AND4_X1   g605(.A1(new_n662), .A2(new_n677), .A3(new_n667), .A4(new_n688), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n791), .A2(new_n792), .A3(new_n759), .A4(new_n750), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n783), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n765), .A2(new_n778), .A3(KEYINPUT53), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT54), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n782), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n486), .B1(new_n722), .B2(new_n723), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n798), .A2(new_n680), .ZN(new_n799));
  INV_X1    g613(.A(new_n659), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n434), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n738), .B(new_n799), .C1(new_n741), .C2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n629), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n660), .A2(new_n697), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n803), .A2(new_n376), .A3(new_n487), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n595), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n798), .A2(new_n804), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n806), .A2(new_n670), .B1(new_n690), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n638), .A2(new_n798), .A3(new_n665), .A4(new_n680), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT50), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n482), .B1(KEYINPUT117), .B2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n815), .A3(KEYINPUT50), .ZN(new_n816));
  OAI22_X1  g630(.A1(new_n810), .A2(new_n813), .B1(KEYINPUT117), .B2(new_n811), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n802), .A2(KEYINPUT51), .A3(new_n809), .A4(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n711), .A2(new_n376), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(new_n808), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT48), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n819), .A2(G952), .A3(new_n239), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n797), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n799), .B1(new_n673), .B2(new_n691), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n818), .A2(new_n809), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT118), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n818), .A2(new_n809), .A3(KEYINPUT118), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n829), .A3(new_n802), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT51), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n830), .A2(KEYINPUT119), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT119), .B1(new_n830), .B2(new_n831), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OR2_X1    g648(.A1(new_n805), .A2(new_n596), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n824), .A2(new_n825), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  OR2_X1    g650(.A1(G952), .A2(G953), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XOR2_X1   g652(.A(new_n659), .B(KEYINPUT49), .Z(new_n839));
  NOR3_X1   g653(.A1(new_n639), .A2(new_n839), .A3(new_n720), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n376), .A2(new_n434), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n840), .A2(new_n483), .A3(new_n803), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n838), .A2(new_n842), .ZN(G75));
  NOR2_X1   g657(.A1(new_n239), .A2(G952), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n468), .A2(new_n472), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(new_n470), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT55), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n189), .B1(new_n794), .B2(new_n795), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(G210), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT56), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n847), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n852));
  XNOR2_X1  g666(.A(new_n848), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n478), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n847), .A2(new_n850), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n844), .B(new_n851), .C1(new_n854), .C2(new_n855), .ZN(G51));
  NAND3_X1  g670(.A1(new_n853), .A2(G469), .A3(new_n729), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n430), .B(KEYINPUT57), .Z(new_n858));
  NAND2_X1  g672(.A1(new_n797), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n423), .B(KEYINPUT121), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n844), .B1(new_n857), .B2(new_n861), .ZN(G54));
  OR2_X1    g676(.A1(new_n848), .A2(KEYINPUT120), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n848), .A2(KEYINPUT120), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n863), .A2(KEYINPUT58), .A3(G475), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n558), .ZN(new_n866));
  INV_X1    g680(.A(new_n558), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n853), .A2(KEYINPUT58), .A3(G475), .A4(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n844), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(G60));
  INV_X1    g684(.A(new_n594), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n588), .B(KEYINPUT59), .Z(new_n872));
  NAND4_X1  g686(.A1(new_n797), .A2(KEYINPUT122), .A3(new_n871), .A4(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n781), .B1(new_n779), .B2(new_n780), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n794), .A2(KEYINPUT54), .A3(new_n795), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n874), .A2(new_n875), .A3(new_n872), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n844), .B1(new_n876), .B2(new_n594), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n874), .A2(new_n875), .A3(new_n871), .A4(new_n872), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n873), .A2(new_n877), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT123), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n873), .A2(new_n877), .A3(KEYINPUT123), .A4(new_n880), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(G63));
  NAND2_X1  g699(.A1(new_n794), .A2(new_n795), .ZN(new_n886));
  NAND2_X1  g700(.A1(G217), .A2(G902), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(KEYINPUT60), .Z(new_n888));
  NAND3_X1  g702(.A1(new_n886), .A2(new_n613), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n886), .A2(new_n888), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n371), .A2(new_n373), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n889), .A2(new_n869), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT61), .B1(new_n889), .B2(new_n894), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n893), .B(new_n895), .ZN(G66));
  OAI21_X1  g710(.A(G953), .B1(new_n489), .B2(new_n441), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n792), .A2(new_n750), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n897), .B1(new_n899), .B2(G953), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n845), .B1(G898), .B2(new_n239), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n900), .B(new_n901), .ZN(G69));
  AND3_X1   g716(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n260), .B(new_n903), .Z(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT126), .ZN(new_n906));
  AOI21_X1  g720(.A(G227), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(G953), .B1(new_n907), .B2(new_n620), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n904), .A2(new_n620), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n906), .B1(new_n909), .B2(G953), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n646), .A2(new_n647), .A3(new_n766), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT62), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n912), .B(new_n913), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n744), .A2(new_n739), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n656), .A2(new_n643), .A3(new_n698), .A4(new_n748), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n914), .A2(new_n904), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  AND2_X1   g731(.A1(new_n739), .A2(new_n766), .ZN(new_n918));
  OR2_X1    g732(.A1(new_n918), .A2(KEYINPUT125), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(KEYINPUT125), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n919), .A2(new_n744), .A3(new_n791), .A4(new_n920), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n736), .A2(new_n820), .A3(new_n685), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n905), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n917), .A2(new_n923), .A3(new_n239), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n924), .A2(new_n908), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n911), .B1(new_n925), .B2(new_n910), .ZN(G72));
  INV_X1    g740(.A(new_n296), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n927), .A2(new_n297), .ZN(new_n928));
  AND4_X1   g742(.A1(new_n899), .A2(new_n914), .A3(new_n915), .A4(new_n916), .ZN(new_n929));
  NAND2_X1  g743(.A1(G472), .A2(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT63), .Z(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n928), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n927), .A2(new_n297), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT127), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n921), .A2(new_n898), .A3(new_n922), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n935), .B1(new_n936), .B2(new_n932), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n577), .A2(new_n298), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n886), .A2(new_n931), .A3(new_n938), .ZN(new_n939));
  AND4_X1   g753(.A1(new_n869), .A2(new_n933), .A3(new_n937), .A4(new_n939), .ZN(G57));
endmodule


