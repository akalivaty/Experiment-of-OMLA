//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 0 1 0 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:20 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT0), .Z(new_n208));
  XNOR2_X1  g0008(.A(KEYINPUT66), .B(G244), .ZN(new_n209));
  AOI22_X1  g0009(.A1(new_n209), .A2(G77), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G50), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT67), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n215), .A2(new_n216), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G87), .A2(G250), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G58), .A2(G232), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  AND2_X1   g0021(.A1(G97), .A2(G257), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n205), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT68), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n201), .A2(KEYINPUT64), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n229), .A2(G50), .A3(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT65), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n208), .B(new_n225), .C1(new_n228), .C2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G68), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT69), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(KEYINPUT70), .B(G107), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n245), .B(new_n249), .ZN(G351));
  INV_X1    g0050(.A(G1), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(G41), .B2(G45), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT71), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G41), .ZN(new_n256));
  OAI211_X1 g0056(.A(G1), .B(G13), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n251), .B(KEYINPUT71), .C1(G41), .C2(G45), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n254), .A2(G238), .A3(new_n257), .A4(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n252), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT77), .ZN(new_n264));
  XNOR2_X1  g0064(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT13), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(G226), .A3(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n267), .A2(G232), .A3(G1698), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G97), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT75), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT75), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G33), .A3(G97), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n269), .A2(new_n270), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT76), .ZN(new_n278));
  INV_X1    g0078(.A(new_n257), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT76), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n269), .A2(new_n270), .A3(new_n276), .A4(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n278), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  AND3_X1   g0082(.A1(new_n265), .A2(new_n266), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n266), .B1(new_n265), .B2(new_n282), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G169), .ZN(new_n286));
  OAI21_X1  g0086(.A(KEYINPUT14), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(G179), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT14), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n289), .B(G169), .C1(new_n283), .C2(new_n284), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n287), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n251), .A2(G20), .ZN(new_n292));
  INV_X1    g0092(.A(G13), .ZN(new_n293));
  OAI21_X1  g0093(.A(KEYINPUT73), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT73), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n295), .A2(new_n251), .A3(G13), .A4(G20), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n213), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n299), .B(KEYINPUT12), .ZN(new_n300));
  NAND3_X1  g0100(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n226), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n255), .A2(G20), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G77), .ZN(new_n305));
  OAI22_X1  g0105(.A1(new_n304), .A2(new_n305), .B1(new_n227), .B2(G68), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n227), .A2(new_n255), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(new_n211), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n302), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n309), .B(KEYINPUT11), .ZN(new_n310));
  INV_X1    g0110(.A(new_n302), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n297), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n312), .B1(new_n251), .B2(G20), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G68), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n300), .A2(new_n310), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n291), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT78), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n285), .A2(G190), .ZN(new_n318));
  INV_X1    g0118(.A(new_n315), .ZN(new_n319));
  INV_X1    g0119(.A(G200), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n318), .B(new_n319), .C1(new_n320), .C2(new_n285), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n316), .A2(new_n317), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n298), .A2(new_n211), .ZN(new_n323));
  INV_X1    g0123(.A(new_n312), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n211), .B1(new_n251), .B2(G20), .ZN(new_n325));
  OR2_X1    g0125(.A1(new_n325), .A2(KEYINPUT74), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(KEYINPUT74), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n324), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  XNOR2_X1  g0128(.A(KEYINPUT8), .B(G58), .ZN(new_n329));
  INV_X1    g0129(.A(G150), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n329), .A2(new_n304), .B1(new_n330), .B2(new_n307), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n227), .B1(new_n201), .B2(new_n211), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n302), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n333), .A2(KEYINPUT72), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n333), .A2(KEYINPUT72), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n323), .B(new_n328), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT9), .ZN(new_n338));
  NOR2_X1   g0138(.A1(G222), .A2(G1698), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n268), .A2(G223), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n267), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n341), .B(new_n279), .C1(G77), .C2(new_n267), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n254), .A2(new_n257), .A3(new_n258), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n342), .B(new_n262), .C1(new_n212), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G200), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT9), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n336), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G190), .ZN(new_n348));
  OR2_X1    g0148(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND4_X1  g0149(.A1(new_n338), .A2(new_n345), .A3(new_n347), .A4(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT10), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n344), .A2(G179), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n344), .A2(new_n286), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n336), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n313), .A2(G77), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n298), .A2(new_n305), .ZN(new_n356));
  XOR2_X1   g0156(.A(KEYINPUT15), .B(G87), .Z(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(new_n304), .ZN(new_n359));
  OAI22_X1  g0159(.A1(new_n329), .A2(new_n307), .B1(new_n227), .B2(new_n305), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n302), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AND3_X1   g0161(.A1(new_n355), .A2(new_n356), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n267), .A2(G238), .A3(G1698), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n267), .A2(G232), .A3(new_n268), .ZN(new_n364));
  INV_X1    g0164(.A(G107), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n363), .B(new_n364), .C1(new_n365), .C2(new_n267), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n279), .ZN(new_n367));
  INV_X1    g0167(.A(new_n343), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n209), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n262), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(G200), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n362), .B(new_n371), .C1(new_n348), .C2(new_n370), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n355), .A2(new_n356), .A3(new_n361), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n370), .A2(new_n286), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n373), .B(new_n374), .C1(G179), .C2(new_n370), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n351), .A2(new_n354), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n317), .B1(new_n316), .B2(new_n321), .ZN(new_n378));
  AND2_X1   g0178(.A1(KEYINPUT3), .A2(G33), .ZN(new_n379));
  NOR2_X1   g0179(.A1(KEYINPUT3), .A2(G33), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT7), .B1(new_n381), .B2(new_n227), .ZN(new_n382));
  OR2_X1    g0182(.A1(KEYINPUT3), .A2(G33), .ZN(new_n383));
  NAND2_X1  g0183(.A1(KEYINPUT3), .A2(G33), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n383), .A2(KEYINPUT7), .A3(new_n227), .A4(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(G68), .B1(new_n382), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G159), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n307), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  AND3_X1   g0190(.A1(KEYINPUT79), .A2(G58), .A3(G68), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT79), .B1(G58), .B2(G68), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n227), .B1(new_n393), .B2(new_n202), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n387), .A2(new_n390), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT16), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n383), .A2(new_n227), .A3(new_n384), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n385), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n394), .B1(new_n401), .B2(G68), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n403), .A3(new_n390), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n311), .B1(new_n397), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n329), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n298), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n313), .B2(new_n329), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  OAI211_X1 g0210(.A(G223), .B(new_n268), .C1(new_n379), .C2(new_n380), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT80), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT80), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n267), .A2(new_n413), .A3(G223), .A4(new_n268), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n267), .A2(G226), .A3(G1698), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G33), .A2(G87), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n412), .A2(new_n414), .A3(new_n415), .A4(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n261), .B1(new_n417), .B2(new_n279), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n368), .A2(G232), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n320), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n405), .A2(new_n410), .A3(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT81), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT17), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n418), .A2(G190), .A3(new_n419), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n421), .A2(new_n422), .A3(new_n423), .A4(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n403), .B1(new_n402), .B2(new_n390), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n213), .B1(new_n400), .B2(new_n385), .ZN(new_n427));
  NOR4_X1   g0227(.A1(new_n427), .A2(KEYINPUT16), .A3(new_n394), .A4(new_n389), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n302), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n417), .A2(new_n279), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(new_n262), .A3(new_n419), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G200), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n429), .A2(new_n424), .A3(new_n409), .A4(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT17), .B1(new_n433), .B2(KEYINPUT81), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n425), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n429), .A2(new_n409), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n431), .A2(G169), .ZN(new_n437));
  INV_X1    g0237(.A(G179), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n437), .B1(new_n438), .B2(new_n431), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT18), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n436), .A2(new_n439), .A3(KEYINPUT18), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n435), .A2(new_n444), .ZN(new_n445));
  NOR4_X1   g0245(.A1(new_n322), .A2(new_n377), .A3(new_n378), .A4(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(G250), .B(G1698), .C1(new_n379), .C2(new_n380), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT83), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT83), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n267), .A2(new_n450), .A3(G250), .A4(G1698), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G283), .ZN(new_n453));
  OAI211_X1 g0253(.A(G244), .B(new_n268), .C1(new_n379), .C2(new_n380), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n454), .A2(KEYINPUT82), .A3(KEYINPUT4), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT4), .B1(new_n454), .B2(KEYINPUT82), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n452), .B(new_n453), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT84), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n449), .A2(new_n451), .B1(G33), .B2(G283), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n460), .B(KEYINPUT84), .C1(new_n455), .C2(new_n456), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(new_n279), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(G45), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n463), .A2(G1), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n256), .A2(KEYINPUT5), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT5), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G41), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n464), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(new_n260), .ZN(new_n469));
  AND2_X1   g0269(.A1(new_n468), .A2(new_n257), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n469), .B1(new_n470), .B2(G257), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n462), .A2(G190), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT85), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n462), .A2(new_n471), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(G200), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n297), .A2(G97), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n255), .A2(G1), .ZN(new_n478));
  AOI211_X1 g0278(.A(new_n478), .B(new_n302), .C1(new_n294), .C2(new_n296), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G97), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n401), .A2(G107), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT6), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n481), .A2(new_n365), .ZN(new_n485));
  NOR2_X1   g0285(.A1(G97), .A2(G107), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n365), .A2(KEYINPUT6), .A3(G97), .ZN(new_n488));
  AND2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI221_X1 g0289(.A(new_n483), .B1(new_n227), .B2(new_n489), .C1(new_n305), .C2(new_n307), .ZN(new_n490));
  AOI211_X1 g0290(.A(new_n477), .B(new_n482), .C1(new_n490), .C2(new_n302), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n462), .A2(KEYINPUT85), .A3(G190), .A4(new_n471), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n474), .A2(new_n476), .A3(new_n491), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n475), .A2(new_n286), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n477), .B1(new_n490), .B2(new_n302), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(new_n481), .B2(new_n480), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n462), .A2(new_n438), .A3(new_n471), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n494), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n479), .A2(G107), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n303), .A2(G116), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n227), .A2(G107), .ZN(new_n502));
  XNOR2_X1  g0302(.A(new_n502), .B(KEYINPUT23), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n227), .B(G87), .C1(new_n379), .C2(new_n380), .ZN(new_n504));
  AND2_X1   g0304(.A1(new_n504), .A2(KEYINPUT22), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n504), .A2(KEYINPUT22), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n501), .B(new_n503), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT24), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g0309(.A(new_n504), .B(KEYINPUT22), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n510), .A2(KEYINPUT24), .A3(new_n501), .A4(new_n503), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n509), .A2(new_n302), .A3(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n297), .A2(G107), .ZN(new_n513));
  XNOR2_X1  g0313(.A(new_n513), .B(KEYINPUT25), .ZN(new_n514));
  OAI211_X1 g0314(.A(G250), .B(new_n268), .C1(new_n379), .C2(new_n380), .ZN(new_n515));
  OAI211_X1 g0315(.A(G257), .B(G1698), .C1(new_n379), .C2(new_n380), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G33), .A2(G294), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n279), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n470), .A2(G264), .ZN(new_n520));
  INV_X1    g0320(.A(new_n469), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G200), .ZN(new_n523));
  AND4_X1   g0323(.A1(new_n500), .A2(new_n512), .A3(new_n514), .A4(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n522), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G190), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n522), .A2(G169), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT89), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n525), .A2(G179), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n522), .A2(KEYINPUT89), .A3(G169), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n512), .A2(new_n500), .A3(new_n514), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n527), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n479), .A2(G116), .ZN(new_n538));
  INV_X1    g0338(.A(G116), .ZN(new_n539));
  AOI22_X1  g0339(.A1(new_n301), .A2(new_n226), .B1(G20), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n453), .B(new_n227), .C1(G33), .C2(new_n481), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT20), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n540), .A2(KEYINPUT20), .A3(new_n541), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n542), .B1(KEYINPUT88), .B2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT88), .ZN(new_n545));
  AOI211_X1 g0345(.A(new_n545), .B(KEYINPUT20), .C1(new_n540), .C2(new_n541), .ZN(new_n546));
  OAI221_X1 g0346(.A(new_n538), .B1(G116), .B2(new_n297), .C1(new_n544), .C2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(G303), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT87), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT87), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G303), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n383), .A2(new_n550), .A3(new_n552), .A4(new_n384), .ZN(new_n553));
  OAI211_X1 g0353(.A(G264), .B(G1698), .C1(new_n379), .C2(new_n380), .ZN(new_n554));
  OAI211_X1 g0354(.A(G257), .B(new_n268), .C1(new_n379), .C2(new_n380), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n279), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n468), .A2(G270), .A3(new_n257), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n557), .A2(G179), .A3(new_n521), .A4(new_n558), .ZN(new_n559));
  OR2_X1    g0359(.A1(new_n548), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n557), .A2(new_n521), .A3(new_n558), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G200), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n548), .B(new_n562), .C1(new_n348), .C2(new_n561), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n547), .A2(G169), .A3(new_n561), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT21), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n547), .A2(KEYINPUT21), .A3(G169), .A4(new_n561), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n560), .A2(new_n563), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n214), .A2(new_n268), .ZN(new_n569));
  INV_X1    g0369(.A(G244), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G1698), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n569), .B(new_n571), .C1(new_n379), .C2(new_n380), .ZN(new_n572));
  NAND2_X1  g0372(.A1(G33), .A2(G116), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n257), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n251), .A2(G45), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n575), .A2(new_n260), .ZN(new_n576));
  AND2_X1   g0376(.A1(G33), .A2(G41), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n575), .B(G250), .C1(new_n577), .C2(new_n226), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n574), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G190), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n297), .A2(new_n357), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n267), .A2(new_n227), .A3(G68), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT19), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n304), .B2(new_n481), .ZN(new_n585));
  AOI21_X1  g0385(.A(G20), .B1(new_n275), .B2(KEYINPUT19), .ZN(new_n586));
  NOR3_X1   g0386(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n583), .B(new_n585), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n582), .B1(new_n588), .B2(new_n302), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n572), .A2(new_n573), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n279), .ZN(new_n591));
  INV_X1    g0391(.A(new_n576), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n592), .A3(new_n578), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G200), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n479), .A2(G87), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n589), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n479), .A2(new_n357), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT86), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n591), .A2(new_n438), .A3(new_n592), .A4(new_n578), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n589), .A2(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n599), .B1(new_n580), .B2(G169), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT86), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n581), .A2(new_n596), .B1(new_n600), .B2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n568), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n499), .A2(new_n537), .A3(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n447), .A2(new_n606), .ZN(G372));
  INV_X1    g0407(.A(new_n354), .ZN(new_n608));
  AND2_X1   g0408(.A1(new_n316), .A2(new_n375), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n321), .A2(new_n435), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n444), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n608), .B1(new_n611), .B2(new_n351), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n535), .A2(new_n560), .A3(new_n567), .A4(new_n566), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n589), .A2(new_n594), .A3(new_n581), .A4(new_n595), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n589), .A2(new_n597), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n614), .B1(new_n615), .B2(new_n601), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n524), .B2(new_n526), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n493), .A2(new_n613), .A3(new_n498), .A4(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n615), .A2(new_n601), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n603), .A2(new_n494), .A3(new_n496), .A4(new_n497), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n619), .B1(new_n620), .B2(KEYINPUT26), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n491), .B1(new_n286), .B2(new_n475), .ZN(new_n622));
  INV_X1    g0422(.A(new_n616), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT26), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n622), .A2(new_n623), .A3(new_n624), .A4(new_n497), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n618), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n612), .B1(new_n447), .B2(new_n627), .ZN(G369));
  NAND3_X1  g0428(.A1(new_n560), .A2(new_n567), .A3(new_n566), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n293), .A2(G20), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  OR3_X1    g0431(.A1(new_n631), .A2(KEYINPUT27), .A3(G1), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT27), .B1(new_n631), .B2(G1), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n632), .A2(G213), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  XNOR2_X1  g0435(.A(KEYINPUT90), .B(G343), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n548), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n629), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n568), .B2(new_n638), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(G330), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(new_n637), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n534), .A2(new_n643), .ZN(new_n644));
  OAI22_X1  g0444(.A1(new_n536), .A2(new_n644), .B1(new_n535), .B2(new_n637), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n535), .A2(new_n643), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n629), .A2(new_n637), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n647), .B1(new_n649), .B2(new_n537), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n646), .A2(new_n650), .ZN(G399));
  INV_X1    g0451(.A(new_n206), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(G41), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n587), .A2(new_n539), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n653), .ZN(new_n656));
  OAI22_X1  g0456(.A1(new_n655), .A2(new_n251), .B1(new_n231), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n657), .B(KEYINPUT28), .ZN(new_n658));
  INV_X1    g0458(.A(G330), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n499), .A2(new_n537), .A3(new_n605), .A4(new_n637), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n519), .A2(new_n520), .ZN(new_n662));
  NOR3_X1   g0462(.A1(new_n559), .A2(new_n662), .A3(new_n593), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n462), .A2(new_n471), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT30), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT30), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n462), .A2(new_n663), .A3(new_n666), .A4(new_n471), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n525), .A2(new_n580), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n475), .A2(new_n669), .A3(new_n438), .A4(new_n561), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n671), .A2(KEYINPUT31), .A3(new_n643), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(KEYINPUT91), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT91), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n668), .A2(new_n675), .A3(new_n670), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n674), .A2(new_n643), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT31), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n673), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n661), .B1(new_n679), .B2(KEYINPUT92), .ZN(new_n680));
  AND3_X1   g0480(.A1(new_n668), .A2(new_n675), .A3(new_n670), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n675), .B1(new_n668), .B2(new_n670), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n681), .A2(new_n682), .A3(new_n637), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n672), .B1(new_n683), .B2(KEYINPUT31), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT92), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n659), .B1(new_n680), .B2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n626), .A2(new_n637), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT93), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(KEYINPUT93), .B1(new_n626), .B2(new_n637), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n691), .A2(KEYINPUT29), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT29), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT26), .B1(new_n498), .B2(new_n616), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n622), .A2(new_n624), .A3(new_n497), .A4(new_n603), .ZN(new_n696));
  INV_X1    g0496(.A(new_n619), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT94), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n695), .A2(new_n696), .A3(KEYINPUT94), .A4(new_n697), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(new_n618), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n694), .B1(new_n702), .B2(new_n637), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n693), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n688), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n658), .B1(new_n706), .B2(G1), .ZN(G364));
  AOI21_X1  g0507(.A(new_n251), .B1(new_n630), .B2(G45), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n653), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n642), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(G330), .B2(new_n640), .ZN(new_n712));
  INV_X1    g0512(.A(new_n710), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n226), .B1(G20), .B2(new_n286), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n348), .A2(G179), .A3(G200), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n227), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(G20), .A2(G179), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G190), .A2(G200), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n718), .A2(G294), .B1(new_n723), .B2(G311), .ZN(new_n724));
  INV_X1    g0524(.A(G326), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n348), .A2(new_n320), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n720), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n724), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT97), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(new_n267), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n719), .A2(new_n320), .A3(G190), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n731), .A2(KEYINPUT96), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(KEYINPUT96), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  XOR2_X1   g0535(.A(KEYINPUT33), .B(G317), .Z(new_n736));
  INV_X1    g0536(.A(G322), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n719), .A2(new_n348), .A3(G200), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  OAI22_X1  g0539(.A1(new_n735), .A2(new_n736), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n227), .A2(G179), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n726), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n740), .B1(G303), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n320), .A2(G190), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G283), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n741), .A2(new_n721), .ZN(new_n749));
  AND2_X1   g0549(.A1(new_n749), .A2(KEYINPUT98), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(KEYINPUT98), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G329), .ZN(new_n754));
  NAND4_X1  g0554(.A1(new_n730), .A2(new_n744), .A3(new_n748), .A4(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G58), .ZN(new_n756));
  OAI22_X1  g0556(.A1(new_n739), .A2(new_n756), .B1(new_n727), .B2(new_n211), .ZN(new_n757));
  INV_X1    g0557(.A(G87), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n742), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n746), .A2(new_n365), .ZN(new_n760));
  NOR4_X1   g0560(.A1(new_n757), .A2(new_n759), .A3(new_n760), .A4(new_n381), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n717), .A2(new_n481), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(G77), .B2(new_n723), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n749), .A2(new_n388), .ZN(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT95), .B(KEYINPUT32), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n734), .A2(G68), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n761), .A2(new_n763), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n715), .B1(new_n755), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(new_n714), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n232), .A2(new_n463), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n652), .A2(new_n267), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n774), .B(new_n775), .C1(new_n245), .C2(new_n463), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n267), .A2(G355), .A3(new_n206), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n776), .B(new_n777), .C1(G116), .C2(new_n206), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n713), .B(new_n769), .C1(new_n773), .C2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n772), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n779), .B1(new_n640), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n712), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(G396));
  OAI21_X1  g0583(.A(new_n376), .B1(new_n362), .B2(new_n637), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n375), .A2(new_n637), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n785), .A2(KEYINPUT100), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n785), .A2(KEYINPUT100), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n784), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n789), .B1(new_n691), .B2(new_n692), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n626), .A2(new_n788), .A3(new_n637), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(KEYINPUT101), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT101), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n626), .A2(new_n788), .A3(new_n793), .A4(new_n637), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n790), .A2(new_n795), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n796), .A2(new_n687), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n687), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n797), .A2(new_n713), .A3(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G283), .ZN(new_n800));
  INV_X1    g0600(.A(G311), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n735), .A2(new_n800), .B1(new_n752), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n746), .A2(new_n758), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n738), .A2(G294), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n267), .B1(new_n743), .B2(G107), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n727), .A2(new_n549), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n807), .B(new_n762), .C1(G116), .C2(new_n723), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n804), .A2(new_n805), .A3(new_n806), .A4(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n727), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n734), .A2(G150), .B1(G137), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n388), .B2(new_n722), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G143), .B2(new_n738), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT34), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G58), .B2(new_n718), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n743), .A2(G50), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n753), .A2(G132), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n815), .A2(new_n267), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n746), .A2(new_n213), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n809), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n714), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n713), .B1(new_n789), .B2(new_n770), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n714), .A2(new_n770), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT99), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n821), .B(new_n822), .C1(G77), .C2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n799), .A2(new_n825), .ZN(G384));
  OAI21_X1  g0626(.A(new_n446), .B1(new_n693), .B2(new_n703), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n612), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT104), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n681), .A2(new_n682), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT105), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n830), .A2(new_n831), .A3(KEYINPUT31), .A4(new_n643), .ZN(new_n832));
  NAND4_X1  g0632(.A1(new_n674), .A2(KEYINPUT31), .A3(new_n643), .A4(new_n676), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(KEYINPUT105), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n677), .A2(new_n678), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n832), .A2(new_n834), .A3(new_n835), .A4(new_n660), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n446), .A2(G330), .A3(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT40), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n316), .B(new_n321), .C1(new_n319), .C2(new_n637), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n291), .A2(new_n315), .A3(new_n643), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n789), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AND3_X1   g0641(.A1(new_n836), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g0642(.A1(KEYINPUT103), .A2(KEYINPUT16), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n396), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n302), .B1(new_n396), .B2(new_n843), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n409), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n445), .A2(new_n635), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n439), .B2(new_n635), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n433), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(KEYINPUT37), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n436), .B1(new_n439), .B2(new_n635), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n433), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n850), .B1(KEYINPUT37), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n847), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT38), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n847), .A2(KEYINPUT38), .A3(new_n853), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT37), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n852), .B(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n436), .A2(new_n635), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n435), .B2(new_n444), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n855), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n857), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n834), .A2(new_n835), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n660), .B1(new_n833), .B2(KEYINPUT105), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n864), .B(new_n841), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n842), .A2(new_n858), .B1(KEYINPUT40), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n837), .B1(new_n868), .B2(new_n659), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(KEYINPUT40), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n858), .A2(new_n836), .A3(new_n838), .A4(new_n841), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(new_n446), .A3(new_n836), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n829), .B(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n442), .A2(new_n443), .A3(new_n634), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n856), .A2(KEYINPUT39), .A3(new_n857), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n857), .A2(new_n863), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n877), .B1(KEYINPUT39), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n316), .A2(new_n643), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n876), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n375), .A2(new_n643), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n795), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n839), .A2(new_n840), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n885), .A2(new_n858), .A3(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n875), .B(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n251), .B2(new_n630), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n393), .A2(G77), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n231), .A2(new_n891), .B1(G50), .B2(new_n213), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(G1), .A3(new_n293), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT35), .ZN(new_n894));
  AOI211_X1 g0694(.A(new_n227), .B(new_n226), .C1(new_n489), .C2(new_n894), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n895), .B(G116), .C1(new_n894), .C2(new_n489), .ZN(new_n896));
  XOR2_X1   g0696(.A(KEYINPUT102), .B(KEYINPUT36), .Z(new_n897));
  XNOR2_X1  g0697(.A(new_n896), .B(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n890), .A2(new_n893), .A3(new_n898), .ZN(G367));
  OAI21_X1  g0699(.A(new_n499), .B1(new_n491), .B2(new_n637), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n900), .A2(new_n535), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n643), .B1(new_n901), .B2(new_n498), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n499), .A2(new_n537), .A3(new_n649), .A4(new_n613), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n903), .B(KEYINPUT42), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT43), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n637), .B1(new_n589), .B2(new_n595), .ZN(new_n906));
  MUX2_X1   g0706(.A(new_n616), .B(new_n697), .S(new_n906), .Z(new_n907));
  OAI22_X1  g0707(.A1(new_n902), .A2(new_n904), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n905), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n908), .B(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n900), .B1(new_n498), .B2(new_n637), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n911), .A2(new_n642), .A3(new_n645), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT106), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n653), .B(KEYINPUT41), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n649), .A2(new_n537), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n645), .B2(new_n649), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n642), .B1(new_n919), .B2(KEYINPUT107), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(KEYINPUT107), .B2(new_n919), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n646), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n705), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n911), .A2(new_n650), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT45), .Z(new_n925));
  NOR2_X1   g0725(.A1(new_n911), .A2(new_n650), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT44), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n923), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n917), .B1(new_n929), .B2(new_n706), .ZN(new_n930));
  OAI221_X1 g0730(.A(new_n915), .B1(new_n709), .B2(new_n930), .C1(new_n913), .C2(new_n910), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n907), .A2(new_n772), .ZN(new_n932));
  INV_X1    g0732(.A(new_n775), .ZN(new_n933));
  OAI221_X1 g0733(.A(new_n773), .B1(new_n206), .B2(new_n358), .C1(new_n240), .C2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n710), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT108), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n267), .B1(new_n735), .B2(new_n388), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(G143), .B2(new_n810), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n718), .A2(G68), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n939), .B1(new_n756), .B2(new_n742), .C1(new_n330), .C2(new_n739), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n940), .B1(G77), .B2(new_n747), .ZN(new_n941));
  AND2_X1   g0741(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(KEYINPUT110), .B(G137), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n942), .B1(new_n211), .B2(new_n722), .C1(new_n749), .C2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT46), .B1(new_n743), .B2(G116), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n743), .A2(KEYINPUT46), .A3(G116), .ZN(new_n947));
  AOI211_X1 g0747(.A(new_n946), .B(new_n947), .C1(G294), .C2(new_n734), .ZN(new_n948));
  INV_X1    g0748(.A(new_n749), .ZN(new_n949));
  AOI22_X1  g0749(.A1(G317), .A2(new_n949), .B1(new_n723), .B2(G283), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n746), .A2(new_n481), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n267), .B1(new_n718), .B2(G107), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n948), .A2(new_n950), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n550), .A2(new_n552), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n739), .A2(new_n955), .B1(new_n727), .B2(new_n801), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT109), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n945), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  XOR2_X1   g0758(.A(new_n958), .B(KEYINPUT47), .Z(new_n959));
  OAI211_X1 g0759(.A(new_n932), .B(new_n936), .C1(new_n959), .C2(new_n715), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n931), .A2(new_n960), .ZN(G387));
  NAND2_X1  g0761(.A1(new_n718), .A2(new_n357), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n949), .A2(G150), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n743), .A2(G77), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n810), .A2(G159), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n962), .A2(new_n963), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n966), .B1(G68), .B2(new_n723), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n381), .B(new_n951), .C1(new_n734), .C2(new_n406), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n967), .B(new_n968), .C1(new_n211), .C2(new_n739), .ZN(new_n969));
  INV_X1    g0769(.A(new_n955), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n970), .A2(new_n723), .B1(new_n738), .B2(G317), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n971), .B1(new_n737), .B2(new_n727), .C1(new_n735), .C2(new_n801), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT48), .ZN(new_n973));
  INV_X1    g0773(.A(G294), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n973), .B1(new_n800), .B2(new_n717), .C1(new_n974), .C2(new_n742), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT111), .Z(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT49), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n381), .B1(new_n749), .B2(new_n725), .C1(new_n539), .C2(new_n746), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT112), .Z(new_n979));
  OAI21_X1  g0779(.A(new_n969), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n713), .B1(new_n980), .B2(new_n714), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n775), .B1(new_n237), .B2(new_n463), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n654), .A2(new_n206), .A3(new_n267), .ZN(new_n983));
  AOI211_X1 g0783(.A(G45), .B(new_n654), .C1(G68), .C2(G77), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n329), .A2(G50), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT50), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n982), .A2(new_n983), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n206), .A2(G107), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n773), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n645), .A2(new_n780), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n981), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n922), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n653), .B1(new_n706), .B2(new_n992), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n991), .B1(new_n708), .B2(new_n922), .C1(new_n993), .C2(new_n923), .ZN(G393));
  XNOR2_X1  g0794(.A(new_n928), .B(new_n646), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n653), .B(new_n929), .C1(new_n995), .C2(new_n923), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n911), .A2(new_n780), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n810), .A2(G150), .B1(G159), .B2(new_n738), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT51), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(G77), .B2(new_n718), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n949), .A2(G143), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n381), .B1(new_n734), .B2(G50), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n722), .A2(new_n329), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n1003), .B(new_n803), .C1(G68), .C2(new_n743), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n810), .A2(G317), .B1(G311), .B2(new_n738), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n743), .A2(G283), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n717), .A2(new_n539), .B1(new_n722), .B2(new_n974), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1010), .B1(new_n734), .B2(new_n970), .ZN(new_n1011));
  AOI211_X1 g0811(.A(new_n267), .B(new_n760), .C1(G322), .C2(new_n949), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1008), .A2(new_n1009), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n715), .B1(new_n1005), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n773), .B1(new_n249), .B2(new_n933), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G97), .B2(new_n652), .ZN(new_n1016));
  NOR3_X1   g0816(.A1(new_n1014), .A2(new_n713), .A3(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n995), .A2(new_n709), .B1(new_n997), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n996), .A2(new_n1018), .ZN(G390));
  AOI21_X1  g0819(.A(new_n883), .B1(new_n792), .B2(new_n794), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n886), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n881), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n879), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n702), .A2(new_n637), .A3(new_n788), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n884), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n886), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n878), .A2(new_n880), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n660), .B1(new_n684), .B2(new_n685), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n679), .A2(KEYINPUT92), .ZN(new_n1030));
  OAI211_X1 g0830(.A(G330), .B(new_n841), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1023), .A2(new_n1028), .A3(new_n1031), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n1022), .A2(new_n879), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n836), .A2(G330), .A3(new_n841), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1032), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1035), .A2(new_n708), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n879), .A2(new_n770), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n718), .A2(G159), .B1(new_n747), .B2(G50), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n735), .B2(new_n944), .ZN(new_n1039));
  INV_X1    g0839(.A(G132), .ZN(new_n1040));
  INV_X1    g0840(.A(G125), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n267), .B1(new_n1040), .B2(new_n739), .C1(new_n752), .C2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(G128), .B2(new_n810), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n742), .A2(new_n330), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT53), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g0846(.A(KEYINPUT54), .B(G143), .Z(new_n1047));
  AOI211_X1 g0847(.A(new_n1039), .B(new_n1046), .C1(new_n723), .C2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n759), .B1(G116), .B2(new_n738), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n305), .B2(new_n717), .C1(new_n752), .C2(new_n974), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n381), .B1(new_n735), .B2(new_n365), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n727), .A2(new_n800), .B1(new_n722), .B2(new_n481), .ZN(new_n1052));
  NOR4_X1   g0852(.A1(new_n1050), .A2(new_n819), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n714), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n710), .B1(new_n824), .B2(new_n406), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT117), .ZN(new_n1056));
  AND3_X1   g0856(.A1(new_n1037), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT116), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n837), .A2(KEYINPUT114), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT114), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n446), .A2(new_n836), .A3(new_n1060), .A4(G330), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1059), .A2(new_n827), .A3(new_n612), .A4(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1025), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1031), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT115), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n836), .B2(G330), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n836), .A2(new_n1066), .A3(G330), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1068), .A2(new_n788), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1065), .B1(new_n1070), .B2(new_n1021), .ZN(new_n1071));
  OAI211_X1 g0871(.A(G330), .B(new_n788), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n1021), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1020), .B1(new_n1073), .B2(new_n1034), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1063), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1058), .B1(new_n1075), .B2(new_n1035), .ZN(new_n1076));
  AND3_X1   g0876(.A1(new_n1023), .A2(new_n1028), .A3(new_n1031), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1034), .B1(new_n1023), .B2(new_n1028), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1069), .A2(new_n788), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1021), .B1(new_n1080), .B2(new_n1067), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1025), .B1(new_n687), .B2(new_n841), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n886), .B1(new_n687), .B2(new_n788), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1034), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n885), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1062), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1079), .A2(new_n1087), .A3(KEYINPUT116), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1076), .A2(new_n1088), .B1(new_n1035), .B2(new_n1075), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1036), .B(new_n1057), .C1(new_n1089), .C2(new_n653), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(G378));
  NOR3_X1   g0891(.A1(new_n1075), .A2(new_n1035), .A3(new_n1058), .ZN(new_n1092));
  AOI21_X1  g0892(.A(KEYINPUT116), .B1(new_n1079), .B2(new_n1087), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1063), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n885), .A2(new_n858), .A3(new_n886), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1095), .B(new_n876), .C1(new_n881), .C2(new_n879), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n351), .A2(new_n354), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n337), .A2(new_n634), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n351), .B(new_n354), .C1(new_n337), .C2(new_n634), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1101), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n872), .B2(G330), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n659), .B(new_n1104), .C1(new_n870), .C2(new_n871), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1096), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1104), .B1(new_n868), .B2(new_n659), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n872), .A2(G330), .A3(new_n1105), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n888), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(KEYINPUT57), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n656), .B1(new_n1094), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT57), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1062), .B1(new_n1076), .B2(new_n1088), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1112), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1120));
  NOR3_X1   g0920(.A1(new_n1106), .A2(new_n1107), .A3(new_n1096), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n888), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n709), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n710), .B1(new_n824), .B2(G50), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT120), .ZN(new_n1125));
  INV_X1    g0925(.A(G124), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n255), .B1(new_n749), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n735), .A2(new_n1040), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n743), .A2(new_n1047), .B1(G128), .B2(new_n738), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT118), .Z(new_n1130));
  AOI211_X1 g0930(.A(new_n1128), .B(new_n1130), .C1(G137), .C2(new_n723), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n1131), .B1(new_n1041), .B2(new_n727), .C1(new_n330), .C2(new_n717), .ZN(new_n1132));
  XOR2_X1   g0932(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1133));
  AOI211_X1 g0933(.A(G41), .B(new_n1127), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1134), .B1(new_n388), .B2(new_n746), .C1(new_n1133), .C2(new_n1132), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n964), .A2(new_n256), .A3(new_n381), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n735), .A2(new_n481), .B1(new_n756), .B2(new_n746), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(G116), .B2(new_n810), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n738), .A2(G107), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n753), .A2(G283), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1138), .A2(new_n939), .A3(new_n1139), .A4(new_n1140), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1136), .B(new_n1141), .C1(new_n357), .C2(new_n723), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1142), .A2(KEYINPUT58), .ZN(new_n1143));
  OR2_X1    g0943(.A1(new_n1142), .A2(KEYINPUT58), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n211), .B1(new_n379), .B2(G41), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1135), .A2(new_n1143), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1125), .B1(new_n1146), .B2(new_n714), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1104), .A2(new_n770), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT121), .B1(new_n1123), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n708), .B1(new_n1108), .B2(new_n1111), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT121), .ZN(new_n1153));
  NOR3_X1   g0953(.A1(new_n1152), .A2(new_n1153), .A3(new_n1149), .ZN(new_n1154));
  OR2_X1    g0954(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1120), .A2(new_n1155), .ZN(G375));
  NOR2_X1   g0956(.A1(new_n824), .A2(G68), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n710), .B1(new_n886), .B2(new_n771), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n267), .B1(new_n723), .B2(G107), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n962), .B(new_n1159), .C1(new_n974), .C2(new_n727), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n753), .A2(G303), .B1(new_n734), .B2(G116), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1161), .B1(new_n305), .B2(new_n746), .C1(new_n481), .C2(new_n742), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1160), .B(new_n1162), .C1(G283), .C2(new_n738), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n734), .A2(new_n1047), .B1(G58), .B2(new_n747), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1164), .B1(new_n211), .B2(new_n717), .C1(new_n388), .C2(new_n742), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n381), .B1(new_n753), .B2(G128), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1166), .B1(new_n1040), .B2(new_n727), .C1(new_n330), .C2(new_n722), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1165), .B(new_n1167), .C1(new_n738), .C2(new_n943), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1163), .A2(new_n1168), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1157), .B(new_n1158), .C1(new_n714), .C2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1170), .B1(new_n1171), .B2(new_n709), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1083), .A2(new_n1086), .A3(new_n1062), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n916), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1172), .B1(new_n1174), .B2(new_n1087), .ZN(G381));
  NOR2_X1   g0975(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n1090), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n931), .A2(new_n960), .A3(new_n1018), .A4(new_n996), .ZN(new_n1179));
  NOR3_X1   g0979(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1180));
  XOR2_X1   g0980(.A(new_n1180), .B(KEYINPUT122), .Z(new_n1181));
  OR4_X1    g0981(.A1(G381), .A2(new_n1178), .A3(new_n1179), .A4(new_n1181), .ZN(G407));
  INV_X1    g0982(.A(G213), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n636), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1177), .A2(new_n1090), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(KEYINPUT123), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1185), .A2(KEYINPUT123), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(G407), .A2(G213), .A3(new_n1186), .A4(new_n1187), .ZN(G409));
  INV_X1    g0988(.A(new_n1184), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1036), .B1(new_n1089), .B2(new_n653), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1094), .A2(new_n916), .A3(new_n1112), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1152), .A2(new_n1149), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1057), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1189), .B(new_n1194), .C1(new_n1177), .C2(new_n1090), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1083), .A2(new_n1086), .A3(KEYINPUT60), .A4(new_n1062), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1075), .A2(new_n1196), .A3(new_n653), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT60), .ZN(new_n1198));
  AND2_X1   g0998(.A1(new_n1173), .A2(new_n1198), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT124), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n799), .A2(new_n1201), .A3(new_n825), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1200), .A2(new_n1172), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1202), .B(new_n1172), .C1(new_n1197), .C2(new_n1199), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1205), .A2(KEYINPUT124), .A3(G384), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1195), .A2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(KEYINPUT125), .B1(new_n1209), .B2(KEYINPUT63), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(G387), .A2(G390), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n1179), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(G393), .B(G396), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1212), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1211), .A2(new_n1213), .A3(new_n1179), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n1209), .B2(KEYINPUT63), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1184), .A2(G2897), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1204), .A2(new_n1206), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1219), .B1(new_n1204), .B2(new_n1206), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(KEYINPUT61), .B1(new_n1195), .B2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT125), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT63), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(new_n1195), .C2(new_n1208), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1210), .A2(new_n1218), .A3(new_n1223), .A4(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1184), .B1(G375), .B2(G378), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT62), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1228), .A2(new_n1229), .A3(new_n1194), .A4(new_n1207), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT62), .B1(new_n1195), .B2(new_n1208), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT126), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1195), .A2(new_n1222), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT61), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1233), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  AOI211_X1 g1036(.A(KEYINPUT126), .B(KEYINPUT61), .C1(new_n1195), .C2(new_n1222), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1232), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1217), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1227), .B1(new_n1238), .B2(new_n1239), .ZN(G405));
  XNOR2_X1  g1040(.A(new_n1217), .B(KEYINPUT127), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT127), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(G375), .A2(G378), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1178), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1208), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1178), .A3(new_n1207), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  MUX2_X1   g1047(.A(new_n1241), .B(new_n1242), .S(new_n1247), .Z(G402));
endmodule


