//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1206, new_n1207,
    new_n1208, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1278, new_n1279, new_n1280;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n203), .A2(G50), .ZN(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT64), .Z(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n210), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n212), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n215), .B(new_n220), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT65), .Z(new_n230));
  NOR2_X1   g0030(.A1(new_n228), .A2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  OAI21_X1  g0048(.A(G20), .B1(new_n203), .B2(G50), .ZN(new_n249));
  INV_X1    g0049(.A(G150), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n249), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT8), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G58), .ZN(new_n256));
  AND3_X1   g0056(.A1(new_n254), .A2(new_n256), .A3(KEYINPUT67), .ZN(new_n257));
  AOI21_X1  g0057(.A(KEYINPUT67), .B1(new_n254), .B2(new_n256), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n210), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n253), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(new_n218), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(G50), .B1(new_n210), .B2(G1), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n267), .B(KEYINPUT68), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(new_n265), .A3(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n270), .B1(G50), .B2(new_n269), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n266), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g0072(.A(new_n272), .B(KEYINPUT9), .Z(new_n273));
  INV_X1    g0073(.A(KEYINPUT71), .ZN(new_n274));
  INV_X1    g0074(.A(G41), .ZN(new_n275));
  INV_X1    g0075(.A(G45), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G1), .A3(G13), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n277), .A2(new_n279), .A3(G274), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n281), .B1(G226), .B2(new_n284), .ZN(new_n285));
  OR2_X1    g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(G223), .ZN(new_n290));
  INV_X1    g0090(.A(G77), .ZN(new_n291));
  OAI22_X1  g0091(.A1(new_n289), .A2(new_n290), .B1(new_n291), .B2(new_n288), .ZN(new_n292));
  AND2_X1   g0092(.A1(KEYINPUT3), .A2(G33), .ZN(new_n293));
  NOR2_X1   g0093(.A1(KEYINPUT3), .A2(G33), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n295), .A2(G1698), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n292), .B1(G222), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n285), .B1(new_n297), .B2(new_n279), .ZN(new_n298));
  INV_X1    g0098(.A(G190), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n274), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT69), .B(G200), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n300), .B1(new_n302), .B2(new_n298), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n273), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n304), .B(KEYINPUT10), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n272), .B1(new_n306), .B2(new_n298), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n307), .B1(G179), .B2(new_n298), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n251), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n311), .B1(new_n291), .B2(new_n260), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n264), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT72), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT72), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n312), .A2(new_n315), .A3(new_n264), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(KEYINPUT11), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT11), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n314), .A2(new_n319), .A3(new_n316), .ZN(new_n320));
  OR3_X1    g0120(.A1(new_n269), .A2(KEYINPUT12), .A3(G68), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT12), .B1(new_n269), .B2(G68), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n263), .B(new_n218), .C1(G1), .C2(new_n210), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n321), .A2(new_n322), .B1(new_n324), .B2(G68), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n318), .A2(new_n320), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT73), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n318), .A2(KEYINPUT73), .A3(new_n320), .A4(new_n325), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT13), .ZN(new_n330));
  INV_X1    g0130(.A(G238), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n280), .B1(new_n331), .B2(new_n283), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n233), .A2(G1698), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n288), .B(new_n334), .C1(G226), .C2(G1698), .ZN(new_n335));
  NAND2_X1  g0135(.A1(G33), .A2(G97), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n330), .B(new_n333), .C1(new_n337), .C2(new_n279), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n279), .B1(new_n335), .B2(new_n336), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT13), .B1(new_n339), .B2(new_n332), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT14), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n341), .A2(new_n342), .A3(G169), .ZN(new_n343));
  INV_X1    g0143(.A(G179), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n343), .B1(new_n344), .B2(new_n341), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n342), .B1(new_n341), .B2(G169), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n328), .B(new_n329), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n328), .A2(new_n329), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n338), .A2(G190), .A3(new_n340), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n341), .A2(G200), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  XOR2_X1   g0152(.A(new_n352), .B(KEYINPUT74), .Z(new_n353));
  INV_X1    g0153(.A(G244), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n280), .B1(new_n354), .B2(new_n283), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n296), .A2(G232), .ZN(new_n356));
  OAI221_X1 g0156(.A(new_n356), .B1(new_n206), .B2(new_n288), .C1(new_n331), .C2(new_n289), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n355), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n306), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n344), .ZN(new_n362));
  INV_X1    g0162(.A(new_n269), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n291), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n291), .B2(new_n323), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n255), .A2(G58), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n369), .A2(new_n251), .B1(G20), .B2(G77), .ZN(new_n370));
  XNOR2_X1  g0170(.A(KEYINPUT15), .B(G87), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n370), .B1(new_n260), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n365), .B1(new_n372), .B2(new_n264), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n361), .A2(new_n362), .A3(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT70), .ZN(new_n377));
  OAI211_X1 g0177(.A(new_n377), .B(new_n373), .C1(new_n359), .C2(new_n301), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n373), .B1(new_n359), .B2(new_n301), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n379), .A2(KEYINPUT70), .B1(G190), .B2(new_n359), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n376), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT16), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n286), .A2(new_n210), .A3(new_n287), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT7), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n286), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n287), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n202), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n201), .A2(new_n202), .ZN(new_n388));
  NOR2_X1   g0188(.A1(G58), .A2(G68), .ZN(new_n389));
  OAI21_X1  g0189(.A(G20), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n251), .A2(G159), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n382), .B1(new_n387), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT7), .B1(new_n295), .B2(new_n210), .ZN(new_n394));
  NOR4_X1   g0194(.A1(new_n293), .A2(new_n294), .A3(new_n384), .A4(G20), .ZN(new_n395));
  OAI21_X1  g0195(.A(G68), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n392), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(KEYINPUT16), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n393), .A2(new_n398), .A3(new_n264), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n269), .B1(new_n257), .B2(new_n258), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT75), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT67), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n366), .B2(new_n367), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n254), .A2(new_n256), .A3(KEYINPUT67), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n403), .A2(new_n404), .A3(new_n323), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n400), .A2(new_n401), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n401), .B1(new_n400), .B2(new_n405), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n399), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(G226), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G1698), .ZN(new_n411));
  OAI221_X1 g0211(.A(new_n411), .B1(G223), .B2(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G87), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n358), .ZN(new_n415));
  INV_X1    g0215(.A(G274), .ZN(new_n416));
  AND2_X1   g0216(.A1(G1), .A2(G13), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n416), .B1(new_n417), .B2(new_n278), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n284), .A2(G232), .B1(new_n277), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n415), .A2(new_n344), .A3(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n279), .B1(new_n412), .B2(new_n413), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n280), .B1(new_n233), .B2(new_n283), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n306), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n409), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT18), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n415), .A2(new_n299), .A3(new_n419), .ZN(new_n428));
  INV_X1    g0228(.A(G200), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n421), .B2(new_n422), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  AND3_X1   g0231(.A1(new_n399), .A2(new_n408), .A3(new_n431), .ZN(new_n432));
  XOR2_X1   g0232(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n424), .B1(new_n399), .B2(new_n408), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT18), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n399), .A2(new_n408), .A3(new_n431), .ZN(new_n438));
  NOR2_X1   g0238(.A1(KEYINPUT76), .A2(KEYINPUT17), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n427), .A2(new_n434), .A3(new_n437), .A4(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  AND4_X1   g0242(.A1(new_n310), .A2(new_n353), .A3(new_n381), .A4(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(G116), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n363), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n209), .A2(G33), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n265), .A2(G116), .A3(new_n269), .A4(new_n447), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n263), .A2(new_n218), .B1(G20), .B2(new_n445), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G283), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n450), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n449), .A2(KEYINPUT20), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT20), .B1(new_n449), .B2(new_n451), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n446), .B(new_n448), .C1(new_n452), .C2(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(G264), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n455));
  INV_X1    g0255(.A(G1698), .ZN(new_n456));
  OAI211_X1 g0256(.A(G257), .B(new_n456), .C1(new_n293), .C2(new_n294), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n286), .A2(G303), .A3(new_n287), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n455), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n358), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n276), .A2(G1), .ZN(new_n461));
  NAND2_X1  g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(KEYINPUT5), .A2(G41), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(G270), .A3(new_n279), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT78), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g0268(.A(KEYINPUT5), .B(G41), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n418), .A2(new_n461), .A3(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n465), .A2(KEYINPUT78), .A3(G270), .A4(new_n279), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n460), .A2(new_n468), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n454), .B1(new_n472), .B2(G200), .ZN(new_n473));
  AND2_X1   g0273(.A1(new_n468), .A2(new_n471), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n474), .A2(G190), .A3(new_n460), .A4(new_n470), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n472), .A2(G169), .A3(new_n454), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT21), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n472), .A2(KEYINPUT21), .A3(G169), .A4(new_n454), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n344), .B1(new_n459), .B2(new_n358), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n474), .A2(new_n470), .A3(new_n454), .A4(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n476), .A2(new_n479), .A3(new_n480), .A4(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT79), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n480), .A2(new_n482), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n486), .A2(KEYINPUT79), .A3(new_n479), .A4(new_n476), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n288), .A2(G244), .A3(G1698), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n288), .A2(G238), .A3(new_n456), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G116), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n358), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n418), .A2(new_n461), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n279), .B(G250), .C1(G1), .C2(new_n276), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n302), .ZN(new_n499));
  INV_X1    g0299(.A(new_n371), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n500), .A2(new_n269), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n265), .A2(new_n269), .A3(new_n447), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n288), .A2(new_n210), .A3(G68), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT19), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n210), .B1(new_n336), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(G87), .B2(new_n207), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n504), .B1(new_n260), .B2(new_n205), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n503), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI221_X4 g0308(.A(new_n501), .B1(new_n502), .B2(G87), .C1(new_n508), .C2(new_n264), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n496), .B1(new_n492), .B2(new_n358), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G190), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n499), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n344), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n501), .B1(new_n508), .B2(new_n264), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n502), .A2(new_n500), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n513), .B(new_n516), .C1(G169), .C2(new_n510), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n465), .A2(G257), .A3(new_n279), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n470), .ZN(new_n520));
  OAI211_X1 g0320(.A(G244), .B(new_n456), .C1(new_n293), .C2(new_n294), .ZN(new_n521));
  XNOR2_X1  g0321(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n288), .A2(KEYINPUT4), .A3(G244), .A4(new_n456), .ZN(new_n524));
  OAI211_X1 g0324(.A(G250), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n523), .A2(new_n524), .A3(new_n450), .A4(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n520), .B1(new_n526), .B2(new_n358), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n306), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT6), .ZN(new_n530));
  NOR3_X1   g0330(.A1(new_n530), .A2(new_n205), .A3(G107), .ZN(new_n531));
  XNOR2_X1  g0331(.A(G97), .B(G107), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n531), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  OAI22_X1  g0333(.A1(new_n533), .A2(new_n210), .B1(new_n291), .B2(new_n252), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n206), .B1(new_n385), .B2(new_n386), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n264), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n269), .A2(G97), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n537), .B1(new_n502), .B2(G97), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n536), .A2(new_n538), .B1(new_n527), .B2(new_n344), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT4), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n450), .B(new_n525), .C1(new_n521), .C2(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n521), .A2(new_n522), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n358), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n520), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(new_n299), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(G200), .B2(new_n527), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n536), .A2(new_n538), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n529), .A2(new_n539), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n518), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT83), .ZN(new_n550));
  OAI211_X1 g0350(.A(KEYINPUT82), .B(KEYINPUT25), .C1(new_n269), .C2(G107), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n363), .A2(new_n206), .ZN(new_n552));
  XNOR2_X1  g0352(.A(KEYINPUT82), .B(KEYINPUT25), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n265), .A2(new_n269), .A3(new_n447), .ZN(new_n554));
  OAI221_X1 g0354(.A(new_n551), .B1(new_n552), .B2(new_n553), .C1(new_n554), .C2(new_n206), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n465), .A2(G264), .A3(new_n279), .ZN(new_n557));
  AND2_X1   g0357(.A1(new_n557), .A2(new_n470), .ZN(new_n558));
  OAI211_X1 g0358(.A(G257), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n559));
  OAI211_X1 g0359(.A(G250), .B(new_n456), .C1(new_n293), .C2(new_n294), .ZN(new_n560));
  INV_X1    g0360(.A(G33), .ZN(new_n561));
  INV_X1    g0361(.A(G294), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n559), .B(new_n560), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n358), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n558), .A2(new_n564), .A3(G190), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n557), .A2(new_n470), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n566), .B1(new_n358), .B2(new_n563), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n556), .B(new_n565), .C1(new_n567), .C2(new_n429), .ZN(new_n568));
  OAI21_X1  g0368(.A(KEYINPUT81), .B1(new_n210), .B2(G107), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(KEYINPUT23), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT23), .ZN(new_n571));
  OAI211_X1 g0371(.A(KEYINPUT81), .B(new_n571), .C1(new_n210), .C2(G107), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n570), .A2(new_n572), .B1(G116), .B2(new_n261), .ZN(new_n573));
  AND2_X1   g0373(.A1(KEYINPUT80), .A2(KEYINPUT22), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n288), .A2(new_n210), .A3(G87), .A4(new_n574), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n210), .B(G87), .C1(new_n293), .C2(new_n294), .ZN(new_n576));
  NOR2_X1   g0376(.A1(KEYINPUT80), .A2(KEYINPUT22), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n573), .A2(new_n575), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT24), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT24), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n573), .A2(new_n582), .A3(new_n579), .A4(new_n575), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n265), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n550), .B1(new_n568), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n581), .A2(new_n583), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n264), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n555), .B1(new_n567), .B2(G190), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n558), .A2(new_n564), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G200), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n587), .A2(new_n588), .A3(KEYINPUT83), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n585), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n587), .A2(new_n556), .ZN(new_n593));
  AOI21_X1  g0393(.A(G169), .B1(new_n558), .B2(new_n564), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n594), .B1(new_n344), .B2(new_n567), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n549), .A2(new_n592), .A3(new_n597), .ZN(new_n598));
  NOR3_X1   g0398(.A1(new_n444), .A2(new_n488), .A3(new_n598), .ZN(G372));
  NAND2_X1  g0399(.A1(new_n486), .A2(new_n479), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n549), .B(new_n592), .C1(new_n600), .C2(new_n596), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n518), .A2(KEYINPUT26), .A3(new_n529), .A4(new_n539), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT26), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n512), .A2(new_n517), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n539), .A2(new_n529), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n602), .A2(KEYINPUT84), .A3(new_n606), .ZN(new_n607));
  OR2_X1    g0407(.A1(new_n606), .A2(KEYINPUT84), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n601), .A2(new_n517), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n443), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g0410(.A(new_n610), .B(KEYINPUT85), .Z(new_n611));
  INV_X1    g0411(.A(new_n305), .ZN(new_n612));
  XNOR2_X1  g0412(.A(new_n435), .B(KEYINPUT18), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n351), .A2(new_n376), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n347), .ZN(new_n616));
  INV_X1    g0416(.A(new_n433), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n438), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n618), .B1(new_n439), .B2(new_n438), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n614), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n308), .B1(new_n612), .B2(new_n620), .ZN(new_n621));
  XOR2_X1   g0421(.A(new_n621), .B(KEYINPUT86), .Z(new_n622));
  NAND2_X1  g0422(.A1(new_n611), .A2(new_n622), .ZN(G369));
  NAND3_X1  g0423(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n624));
  OR2_X1    g0424(.A1(new_n624), .A2(KEYINPUT27), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(KEYINPUT27), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(G213), .A3(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(G343), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n454), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g0430(.A(new_n630), .B(KEYINPUT87), .Z(new_n631));
  NOR2_X1   g0431(.A1(new_n488), .A2(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n600), .A2(new_n631), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(G330), .ZN(new_n635));
  OR3_X1    g0435(.A1(new_n634), .A2(KEYINPUT88), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(KEYINPUT88), .B1(new_n634), .B2(new_n635), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n597), .A2(new_n629), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n593), .A2(new_n629), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n596), .B1(new_n592), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n629), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n600), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n639), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n643), .A2(new_n650), .ZN(G399));
  INV_X1    g0451(.A(new_n213), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n652), .A2(G41), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G1), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n656), .B1(new_n216), .B2(new_n654), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n657), .B(KEYINPUT28), .ZN(new_n658));
  INV_X1    g0458(.A(new_n517), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(new_n602), .B2(new_n606), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n629), .B1(new_n601), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT29), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n609), .A2(new_n644), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n664), .B1(KEYINPUT29), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT30), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n567), .A2(new_n474), .A3(new_n510), .A4(new_n481), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n667), .B1(new_n668), .B2(new_n528), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n567), .A2(new_n510), .A3(G179), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n670), .A2(new_n472), .A3(new_n528), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n474), .A2(new_n510), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n481), .A2(new_n558), .A3(new_n564), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n672), .A2(KEYINPUT30), .A3(new_n527), .A4(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n669), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n629), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT31), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n675), .A2(KEYINPUT31), .A3(new_n629), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n629), .B1(new_n593), .B2(new_n595), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n592), .A2(new_n681), .A3(new_n548), .A4(new_n518), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT89), .B1(new_n488), .B2(new_n682), .ZN(new_n683));
  AND4_X1   g0483(.A1(new_n592), .A2(new_n681), .A3(new_n548), .A4(new_n518), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT89), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n485), .A2(new_n487), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n680), .B1(new_n683), .B2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(new_n635), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n666), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n658), .B1(new_n690), .B2(G1), .ZN(G364));
  AND2_X1   g0491(.A1(new_n210), .A2(G13), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n209), .B1(new_n692), .B2(G45), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n653), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n213), .A2(new_n288), .ZN(new_n696));
  INV_X1    g0496(.A(G355), .ZN(new_n697));
  OAI22_X1  g0497(.A1(new_n696), .A2(new_n697), .B1(G116), .B2(new_n213), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n652), .A2(new_n288), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n700), .B1(new_n217), .B2(new_n276), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n247), .A2(G45), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n698), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OR3_X1    g0503(.A1(KEYINPUT90), .A2(G13), .A3(G33), .ZN(new_n704));
  OAI21_X1  g0504(.A(KEYINPUT90), .B1(G13), .B2(G33), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G20), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n218), .B1(G20), .B2(new_n306), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n695), .B1(new_n703), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n302), .A2(KEYINPUT92), .A3(new_n344), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT92), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(new_n301), .B2(G179), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n713), .A2(G20), .A3(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n299), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n718), .A2(KEYINPUT93), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(KEYINPUT93), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(G303), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n295), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  XOR2_X1   g0523(.A(new_n723), .B(KEYINPUT95), .Z(new_n724));
  NOR2_X1   g0524(.A1(new_n210), .A2(new_n344), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n725), .B(KEYINPUT91), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n726), .A2(G190), .A3(G200), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n726), .A2(new_n299), .A3(G200), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n727), .A2(G311), .B1(new_n728), .B2(G322), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n725), .A2(G200), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n299), .ZN(new_n731));
  NOR2_X1   g0531(.A1(G190), .A2(G200), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(G20), .A3(new_n344), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n731), .A2(G326), .B1(G329), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n730), .A2(G190), .ZN(new_n736));
  XNOR2_X1  g0536(.A(KEYINPUT33), .B(G317), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n344), .A2(new_n429), .A3(G190), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G20), .ZN(new_n739));
  AOI22_X1  g0539(.A1(new_n736), .A2(new_n737), .B1(new_n739), .B2(G294), .ZN(new_n740));
  AND3_X1   g0540(.A1(new_n729), .A2(new_n735), .A3(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(G283), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n716), .A2(G190), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n724), .B(new_n741), .C1(new_n742), .C2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n721), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G87), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n743), .A2(G107), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n747), .A2(new_n288), .A3(new_n748), .ZN(new_n749));
  XOR2_X1   g0549(.A(new_n749), .B(KEYINPUT94), .Z(new_n750));
  INV_X1    g0550(.A(G159), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n733), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT32), .ZN(new_n753));
  AOI22_X1  g0553(.A1(new_n731), .A2(G50), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n728), .ZN(new_n755));
  INV_X1    g0555(.A(new_n727), .ZN(new_n756));
  OAI221_X1 g0556(.A(new_n754), .B1(new_n755), .B2(new_n201), .C1(new_n291), .C2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n739), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n205), .ZN(new_n759));
  INV_X1    g0559(.A(new_n736), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n760), .A2(new_n202), .B1(new_n753), .B2(new_n752), .ZN(new_n761));
  OR3_X1    g0561(.A1(new_n757), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n745), .B1(new_n750), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n712), .B1(new_n763), .B2(new_n709), .ZN(new_n764));
  INV_X1    g0564(.A(new_n634), .ZN(new_n765));
  INV_X1    g0565(.A(new_n708), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n695), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n768), .B1(new_n765), .B2(G330), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n767), .B1(new_n638), .B2(new_n769), .ZN(G396));
  NOR2_X1   g0570(.A1(new_n375), .A2(new_n629), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n380), .A2(new_n378), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n374), .A2(new_n629), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n771), .B1(new_n774), .B2(new_n375), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n665), .B(new_n775), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n776), .A2(new_n689), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n689), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n777), .A2(new_n768), .A3(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n706), .A2(new_n709), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n768), .B1(new_n291), .B2(new_n780), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n736), .A2(G150), .B1(new_n731), .B2(G137), .ZN(new_n782));
  INV_X1    g0582(.A(G143), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n782), .B1(new_n755), .B2(new_n783), .C1(new_n751), .C2(new_n756), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT34), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n743), .A2(G68), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n784), .A2(new_n785), .ZN(new_n789));
  INV_X1    g0589(.A(G132), .ZN(new_n790));
  OAI221_X1 g0590(.A(new_n288), .B1(new_n790), .B2(new_n733), .C1(new_n758), .C2(new_n201), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n746), .A2(G50), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n746), .A2(G107), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n743), .A2(G87), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n727), .A2(G116), .B1(new_n728), .B2(G294), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n288), .B(new_n759), .C1(G311), .C2(new_n734), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n736), .A2(G283), .B1(new_n731), .B2(G303), .ZN(new_n798));
  AND4_X1   g0598(.A1(new_n795), .A2(new_n796), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n792), .A2(new_n793), .B1(new_n794), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n709), .ZN(new_n801));
  OAI221_X1 g0601(.A(new_n781), .B1(new_n800), .B2(new_n801), .C1(new_n707), .C2(new_n775), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n779), .A2(new_n802), .ZN(G384));
  INV_X1    g0603(.A(new_n533), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n804), .A2(KEYINPUT35), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(KEYINPUT35), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n805), .A2(G116), .A3(new_n219), .A4(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT36), .Z(new_n808));
  OR3_X1    g0608(.A1(new_n216), .A2(new_n291), .A3(new_n388), .ZN(new_n809));
  INV_X1    g0609(.A(G50), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G68), .ZN(new_n811));
  AOI211_X1 g0611(.A(new_n209), .B(G13), .C1(new_n809), .C2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n328), .A2(new_n329), .A3(new_n629), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n347), .A2(new_n351), .A3(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n814), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n346), .B2(new_n345), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n609), .A2(new_n644), .A3(new_n775), .ZN(new_n820));
  INV_X1    g0620(.A(new_n771), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT38), .ZN(new_n823));
  AND3_X1   g0623(.A1(new_n403), .A2(new_n404), .A3(new_n323), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n363), .B1(new_n403), .B2(new_n404), .ZN(new_n825));
  OAI21_X1  g0625(.A(KEYINPUT75), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n400), .A2(new_n405), .A3(new_n401), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n396), .A2(new_n397), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n265), .B1(new_n829), .B2(new_n382), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n828), .B1(new_n830), .B2(new_n398), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(new_n627), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n823), .B1(new_n441), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n438), .B1(new_n831), .B2(new_n424), .ZN(new_n834));
  OAI21_X1  g0634(.A(KEYINPUT37), .B1(new_n834), .B2(new_n832), .ZN(new_n835));
  INV_X1    g0635(.A(new_n627), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n409), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT37), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n426), .A2(new_n837), .A3(new_n838), .A4(new_n438), .ZN(new_n839));
  AND3_X1   g0639(.A1(new_n835), .A2(KEYINPUT96), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT96), .B1(new_n835), .B2(new_n839), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n833), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n837), .B1(new_n619), .B2(new_n613), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT96), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n432), .A2(new_n435), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n838), .B1(new_n845), .B2(new_n837), .ZN(new_n846));
  AND4_X1   g0646(.A1(new_n838), .A2(new_n426), .A3(new_n837), .A4(new_n438), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n844), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n835), .A2(KEYINPUT96), .A3(new_n839), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n843), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n842), .B1(new_n850), .B2(KEYINPUT38), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n822), .A2(new_n851), .B1(new_n614), .B2(new_n627), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT97), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n842), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT39), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n848), .A2(new_n849), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n857), .A2(KEYINPUT97), .A3(new_n833), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n846), .A2(new_n847), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n823), .B1(new_n859), .B2(new_n843), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n855), .A2(new_n856), .A3(new_n858), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n851), .A2(KEYINPUT39), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT98), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n863), .B1(new_n861), .B2(new_n862), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n347), .A2(new_n629), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n853), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n443), .A2(new_n666), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n622), .A2(new_n869), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n868), .B(new_n870), .Z(new_n871));
  NOR2_X1   g0671(.A1(new_n444), .A2(new_n688), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT40), .ZN(new_n873));
  INV_X1    g0673(.A(new_n680), .ZN(new_n874));
  NOR3_X1   g0674(.A1(new_n488), .A2(KEYINPUT89), .A3(new_n682), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n685), .B1(new_n684), .B2(new_n686), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI22_X1  g0677(.A1(new_n380), .A2(new_n378), .B1(new_n374), .B2(new_n629), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n821), .B1(new_n878), .B2(new_n376), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n879), .B1(new_n815), .B2(new_n817), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n441), .A2(new_n832), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n840), .B2(new_n841), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n883), .A2(new_n823), .B1(new_n857), .B2(new_n833), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n873), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n818), .A2(new_n775), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n688), .A2(new_n886), .A3(new_n873), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n855), .A2(new_n858), .A3(new_n860), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n635), .B1(new_n872), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n891), .B1(new_n890), .B2(new_n872), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n871), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n209), .B2(new_n692), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n871), .A2(new_n892), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n813), .B1(new_n894), .B2(new_n895), .ZN(G367));
  INV_X1    g0696(.A(KEYINPUT101), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n548), .B1(new_n547), .B2(new_n644), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n539), .A2(new_n529), .A3(new_n629), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n897), .B1(new_n647), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n642), .A2(KEYINPUT101), .A3(new_n646), .A4(new_n900), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT42), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n605), .B1(new_n898), .B2(new_n597), .ZN(new_n907));
  OR2_X1    g0707(.A1(new_n907), .A2(KEYINPUT100), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n644), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n909), .B1(KEYINPUT100), .B2(new_n907), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n906), .A2(new_n911), .A3(KEYINPUT102), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT102), .B1(new_n906), .B2(new_n911), .ZN(new_n913));
  NOR3_X1   g0713(.A1(new_n903), .A2(KEYINPUT42), .A3(new_n905), .ZN(new_n914));
  OR3_X1    g0714(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT103), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n509), .A2(new_n644), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n659), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n604), .B2(new_n917), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT43), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n915), .A2(new_n916), .A3(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n919), .A2(KEYINPUT43), .ZN(new_n922));
  XNOR2_X1  g0722(.A(new_n922), .B(KEYINPUT99), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n916), .B1(new_n915), .B2(new_n920), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n643), .A2(new_n901), .ZN(new_n928));
  OR3_X1    g0728(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(new_n690), .ZN(new_n930));
  INV_X1    g0730(.A(new_n642), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n638), .B(new_n931), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(new_n646), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  XOR2_X1   g0734(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n935));
  NAND3_X1  g0735(.A1(new_n650), .A2(new_n900), .A3(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n935), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n937), .B1(new_n649), .B2(new_n901), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n649), .A2(KEYINPUT44), .A3(new_n901), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT44), .B1(new_n649), .B2(new_n901), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n936), .B(new_n938), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(new_n643), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n930), .B1(new_n934), .B2(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n653), .B(KEYINPUT41), .Z(new_n944));
  OAI21_X1  g0744(.A(new_n693), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n928), .B1(new_n926), .B2(new_n927), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n929), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n711), .B1(new_n652), .B2(new_n500), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n699), .A2(new_n239), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n768), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n744), .A2(new_n291), .ZN(new_n951));
  INV_X1    g0751(.A(G137), .ZN(new_n952));
  INV_X1    g0752(.A(new_n731), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n288), .B1(new_n733), .B2(new_n952), .C1(new_n953), .C2(new_n783), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n739), .A2(G68), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n760), .B2(new_n751), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n957), .B1(new_n810), .B2(new_n756), .C1(new_n250), .C2(new_n755), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n951), .B(new_n958), .C1(new_n746), .C2(G58), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n288), .B1(new_n734), .B2(G317), .ZN(new_n960));
  INV_X1    g0760(.A(G311), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n960), .B1(new_n953), .B2(new_n961), .C1(new_n562), .C2(new_n760), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n755), .A2(new_n722), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n727), .A2(G283), .B1(G107), .B2(new_n739), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n962), .B(new_n963), .C1(KEYINPUT105), .C2(new_n964), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n965), .B1(KEYINPUT105), .B2(new_n964), .C1(new_n205), .C2(new_n744), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT106), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT46), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n721), .A2(new_n445), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n969), .A2(new_n970), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n959), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n973), .A2(KEYINPUT47), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n709), .B1(new_n973), .B2(KEYINPUT47), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n950), .B1(new_n766), .B2(new_n919), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n947), .A2(new_n976), .ZN(G387));
  NOR2_X1   g0777(.A1(new_n933), .A2(new_n930), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n933), .A2(new_n930), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n979), .A2(new_n980), .A3(new_n653), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n696), .A2(new_n655), .B1(G107), .B2(new_n213), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n700), .B1(new_n236), .B2(G45), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n368), .A2(G50), .ZN(new_n984));
  XNOR2_X1  g0784(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n984), .B(new_n985), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n655), .B(new_n276), .C1(new_n202), .C2(new_n291), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT107), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(new_n988), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n982), .B1(new_n983), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n695), .B1(new_n992), .B2(new_n711), .ZN(new_n993));
  INV_X1    g0793(.A(G322), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n760), .A2(new_n961), .B1(new_n953), .B2(new_n994), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n995), .A2(KEYINPUT109), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(KEYINPUT109), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n727), .A2(G303), .B1(new_n728), .B2(G317), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n996), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT48), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n742), .B2(new_n758), .C1(new_n562), .C2(new_n721), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT110), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1002), .A2(KEYINPUT49), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(KEYINPUT49), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n744), .A2(new_n445), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n288), .B(new_n1005), .C1(G326), .C2(new_n734), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1003), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n288), .B1(new_n250), .B2(new_n733), .C1(new_n758), .C2(new_n371), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n728), .A2(G50), .B1(new_n259), .B2(new_n736), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n202), .B2(new_n756), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1008), .B(new_n1010), .C1(G159), .C2(new_n731), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n205), .B2(new_n744), .C1(new_n721), .C2(new_n291), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n801), .B1(new_n1007), .B2(new_n1012), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n993), .B(new_n1013), .C1(new_n931), .C2(new_n708), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n934), .B2(new_n694), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n981), .A2(new_n1015), .ZN(G393));
  AOI21_X1  g0816(.A(new_n654), .B1(new_n978), .B2(new_n942), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n978), .A2(new_n942), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n1018), .A2(KEYINPUT112), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1018), .A2(KEYINPUT112), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1017), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n901), .A2(new_n708), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n244), .A2(new_n700), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n710), .B1(new_n205), .B2(new_n213), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n695), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n758), .A2(new_n291), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n288), .B1(new_n733), .B2(new_n783), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n755), .A2(new_n751), .B1(new_n250), .B2(new_n953), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT51), .ZN(new_n1029));
  AOI211_X1 g0829(.A(new_n1026), .B(new_n1027), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n727), .A2(new_n369), .B1(G50), .B2(new_n736), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT111), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1030), .A2(new_n795), .A3(new_n1031), .A4(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n721), .A2(new_n202), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n721), .A2(new_n742), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n731), .A2(G317), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n755), .B2(new_n961), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT52), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n758), .A2(new_n445), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n295), .B1(new_n733), .B2(new_n994), .C1(new_n760), .C2(new_n722), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(G294), .C2(new_n727), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1040), .A2(new_n1043), .A3(new_n748), .A4(new_n1044), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n1034), .A2(new_n1035), .B1(new_n1036), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1025), .B1(new_n1046), .B2(new_n709), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n942), .A2(new_n694), .B1(new_n1022), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1021), .A2(new_n1048), .ZN(G390));
  NAND3_X1  g0849(.A1(new_n689), .A2(new_n775), .A3(new_n818), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(KEYINPUT113), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n1051), .A2(KEYINPUT113), .ZN(new_n1053));
  NOR2_X1   g0853(.A1(new_n822), .A2(new_n867), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n861), .A2(new_n862), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(KEYINPUT98), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1054), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n774), .A2(new_n375), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n771), .B1(new_n661), .B2(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n1060), .A2(new_n819), .B1(new_n347), .B2(new_n629), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n888), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1052), .B(new_n1053), .C1(new_n1058), .C2(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n864), .A2(new_n865), .B1(new_n822), .B2(new_n867), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1063), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n1065), .A2(KEYINPUT113), .A3(new_n1051), .A4(new_n1066), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n693), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n866), .A2(new_n707), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n259), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n768), .B1(new_n1071), .B2(new_n780), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n721), .A2(new_n250), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT53), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n288), .B1(new_n744), .B2(new_n810), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n1075), .A2(KEYINPUT114), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1075), .A2(KEYINPUT114), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n736), .A2(G137), .B1(G125), .B2(new_n734), .ZN(new_n1079));
  INV_X1    g0879(.A(G128), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1079), .B1(new_n1080), .B2(new_n953), .C1(new_n751), .C2(new_n758), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(KEYINPUT54), .B(G143), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n790), .A2(new_n755), .B1(new_n756), .B2(new_n1082), .ZN(new_n1083));
  NOR4_X1   g0883(.A1(new_n1077), .A2(new_n1078), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n727), .A2(G97), .B1(new_n728), .B2(G116), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n288), .B(new_n1026), .C1(G294), .C2(new_n734), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n736), .A2(G107), .B1(new_n731), .B2(G283), .ZN(new_n1087));
  AND4_X1   g0887(.A1(new_n787), .A2(new_n1085), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1074), .A2(new_n1084), .B1(new_n747), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1072), .B1(new_n1089), .B2(new_n801), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1070), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1069), .A2(KEYINPUT115), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT115), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n1068), .B2(new_n1091), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n443), .A2(new_n689), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n622), .A2(new_n869), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n820), .A2(new_n821), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n818), .B1(new_n689), .B2(new_n775), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1100), .B1(new_n1051), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1101), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(new_n1050), .A3(new_n1060), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1099), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1097), .A2(new_n1105), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n1106), .A2(new_n654), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1097), .A2(new_n1105), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1096), .A2(new_n1109), .ZN(G378));
  NAND3_X1  g0910(.A1(new_n885), .A2(new_n889), .A3(G330), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT118), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n885), .A2(new_n889), .A3(KEYINPUT118), .A4(G330), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n836), .B1(new_n266), .B2(new_n271), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT55), .Z(new_n1116));
  NAND2_X1  g0916(.A1(new_n309), .A2(new_n1116), .ZN(new_n1117));
  XOR2_X1   g0917(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1118));
  INV_X1    g0918(.A(new_n1116), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n305), .A2(new_n308), .A3(new_n1119), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1117), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1118), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1113), .A2(new_n1114), .A3(new_n1124), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n890), .A2(new_n1123), .A3(KEYINPUT118), .A4(G330), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n868), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1125), .A2(new_n868), .A3(new_n1126), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1129), .A2(KEYINPUT57), .A3(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1099), .B1(new_n1097), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n653), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT57), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1099), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1108), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1129), .A2(KEYINPUT119), .A3(new_n1130), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT119), .ZN(new_n1139));
  AND3_X1   g0939(.A1(new_n1125), .A2(new_n868), .A3(new_n1126), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n866), .A2(new_n867), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1125), .A2(new_n1126), .B1(new_n1141), .B2(new_n852), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1139), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1137), .A2(new_n1138), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1134), .B1(new_n1135), .B2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1143), .A2(new_n1138), .A3(new_n694), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1123), .A2(new_n706), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n780), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n695), .B1(G50), .B2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n288), .A2(G41), .ZN(new_n1150));
  AOI211_X1 g0950(.A(G50), .B(new_n1150), .C1(new_n561), .C2(new_n275), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n743), .A2(G58), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT116), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n206), .A2(new_n755), .B1(new_n756), .B2(new_n371), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n955), .B(new_n1150), .C1(new_n742), .C2(new_n733), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n760), .A2(new_n205), .B1(new_n953), .B2(new_n445), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  OAI211_X1 g0957(.A(new_n1153), .B(new_n1157), .C1(new_n721), .C2(new_n291), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT58), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1151), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n760), .A2(new_n790), .B1(new_n758), .B2(new_n250), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(G125), .B2(new_n731), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n727), .A2(G137), .B1(new_n728), .B2(G128), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(new_n721), .C2(new_n1082), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n743), .A2(G159), .ZN(new_n1166));
  AOI211_X1 g0966(.A(G33), .B(G41), .C1(new_n734), .C2(G124), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1160), .B1(new_n1159), .B2(new_n1158), .C1(new_n1168), .C2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1149), .B1(new_n1170), .B2(new_n709), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1147), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1146), .A2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1145), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(G375));
  NAND2_X1  g0975(.A1(new_n1136), .A2(new_n1132), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n944), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1099), .A2(new_n1102), .A3(new_n1104), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n693), .B(KEYINPUT120), .Z(new_n1180));
  NAND2_X1  g0980(.A1(new_n1132), .A2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n768), .B1(new_n202), .B2(new_n780), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n295), .B1(new_n733), .B2(new_n722), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n760), .A2(new_n445), .B1(new_n953), .B2(new_n562), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(new_n500), .C2(new_n739), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1185), .B1(new_n206), .B2(new_n756), .C1(new_n742), .C2(new_n755), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n951), .B(new_n1186), .C1(new_n746), .C2(G97), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1187), .A2(KEYINPUT121), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(KEYINPUT121), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n952), .A2(new_n755), .B1(new_n756), .B2(new_n250), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n288), .B1(new_n733), .B2(new_n1080), .C1(new_n760), .C2(new_n1082), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n953), .A2(new_n790), .B1(new_n758), .B2(new_n810), .ZN(new_n1192));
  NOR3_X1   g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1153), .B(new_n1193), .C1(new_n721), .C2(new_n751), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1188), .A2(new_n1189), .A3(new_n1194), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1182), .B1(new_n707), .B2(new_n818), .C1(new_n1195), .C2(new_n801), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1181), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1179), .A2(new_n1198), .ZN(G381));
  OR2_X1    g0999(.A1(G393), .A2(G396), .ZN(new_n1200));
  INV_X1    g1000(.A(G384), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1179), .A2(new_n1198), .A3(new_n1201), .ZN(new_n1202));
  NOR4_X1   g1002(.A1(G387), .A2(G390), .A3(new_n1200), .A4(new_n1202), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1095), .A2(new_n1093), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1203), .A2(new_n1204), .A3(new_n1174), .ZN(G407));
  NAND2_X1  g1005(.A1(new_n628), .A2(G213), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT122), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1174), .A2(new_n1204), .A3(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(G407), .A2(G213), .A3(new_n1208), .ZN(G409));
  AOI21_X1  g1009(.A(G390), .B1(new_n947), .B2(new_n976), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT125), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(G393), .A2(G396), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1200), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1212), .B1(new_n1200), .B2(new_n1213), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(G390), .A2(new_n947), .A3(new_n976), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1211), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1217), .ZN(new_n1219));
  OAI22_X1  g1019(.A1(new_n1219), .A2(new_n1210), .B1(new_n1215), .B2(new_n1214), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT61), .B1(new_n1218), .B2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1173), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1140), .A2(new_n1142), .A3(new_n1139), .ZN(new_n1223));
  AOI21_X1  g1023(.A(KEYINPUT119), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(KEYINPUT57), .B1(new_n1225), .B2(new_n1137), .ZN(new_n1226));
  OAI211_X1 g1026(.A(G378), .B(new_n1222), .C1(new_n1226), .C2(new_n1134), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1137), .A2(new_n1143), .A3(new_n1177), .A4(new_n1138), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1229), .A2(new_n1180), .B1(new_n1147), .B2(new_n1171), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1204), .A2(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1207), .B1(new_n1227), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1176), .A2(new_n653), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1178), .A2(KEYINPUT123), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT60), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1178), .A2(KEYINPUT123), .A3(KEYINPUT60), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1234), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1240), .A2(G384), .A3(new_n1198), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1201), .B1(new_n1239), .B2(new_n1197), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1233), .A2(KEYINPUT63), .A3(new_n1244), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1145), .A2(new_n1204), .A3(new_n1173), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1232), .ZN(new_n1247));
  OAI211_X1 g1047(.A(new_n1206), .B(new_n1244), .C1(new_n1246), .C2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT63), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1206), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1206), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(G2897), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1241), .A2(new_n1242), .A3(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT124), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1241), .A2(new_n1242), .A3(KEYINPUT124), .A4(new_n1253), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1243), .A2(G2897), .A3(new_n1207), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1251), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  NAND4_X1  g1060(.A1(new_n1221), .A2(new_n1245), .A3(new_n1250), .A4(new_n1260), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT61), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1263), .B1(new_n1264), .B2(new_n1233), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1241), .A2(new_n1242), .A3(KEYINPUT62), .ZN(new_n1266));
  AOI211_X1 g1066(.A(new_n1207), .B(new_n1266), .C1(new_n1227), .C2(new_n1232), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT62), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1267), .A2(KEYINPUT126), .B1(new_n1248), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT126), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1233), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1270), .B1(new_n1271), .B2(new_n1266), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1265), .B1(new_n1269), .B2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT127), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1262), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  AOI211_X1 g1075(.A(KEYINPUT127), .B(new_n1265), .C1(new_n1269), .C2(new_n1272), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1261), .B1(new_n1275), .B2(new_n1276), .ZN(G405));
  NAND2_X1  g1077(.A1(G375), .A2(new_n1204), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1278), .A2(new_n1227), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1279), .B(new_n1244), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1262), .B(new_n1280), .ZN(G402));
endmodule


