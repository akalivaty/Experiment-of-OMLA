//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT1), .B1(new_n188), .B2(G146), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G146), .ZN(new_n192));
  AOI22_X1  g006(.A1(new_n189), .A2(G128), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT64), .B1(new_n190), .B2(G143), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(new_n188), .A3(G146), .ZN(new_n196));
  AOI22_X1  g010(.A1(new_n194), .A2(new_n196), .B1(G143), .B2(new_n190), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n198), .B1(new_n191), .B2(KEYINPUT1), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n193), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(G125), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT0), .A2(G128), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT0), .A2(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n191), .A2(new_n192), .ZN(new_n206));
  AOI22_X1  g020(.A1(new_n197), .A2(new_n203), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n201), .B1(G125), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G224), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G953), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n208), .B(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(G110), .B(G122), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT4), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT78), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT78), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT3), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT79), .B(G107), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n219), .A2(new_n220), .A3(G104), .ZN(new_n221));
  INV_X1    g035(.A(G107), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n215), .B1(new_n222), .B2(G104), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(G104), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(KEYINPUT80), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n222), .A2(KEYINPUT79), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT79), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(G107), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(new_n229), .A3(G104), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT78), .B(KEYINPUT3), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n225), .B(KEYINPUT80), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n214), .B(G101), .C1(new_n226), .C2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G119), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G116), .ZN(new_n236));
  INV_X1    g050(.A(G116), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G119), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT2), .B(G113), .ZN(new_n240));
  OR2_X1    g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n240), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G101), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n225), .B1(new_n230), .B2(new_n231), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT80), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n244), .B1(new_n247), .B2(new_n232), .ZN(new_n248));
  OAI211_X1 g062(.A(new_n225), .B(new_n244), .C1(new_n230), .C2(new_n231), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT4), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n234), .B(new_n243), .C1(new_n248), .C2(new_n250), .ZN(new_n251));
  AND3_X1   g065(.A1(new_n236), .A2(new_n238), .A3(KEYINPUT5), .ZN(new_n252));
  OAI21_X1  g066(.A(G113), .B1(new_n236), .B2(KEYINPUT5), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n241), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(G104), .B1(new_n227), .B2(new_n229), .ZN(new_n255));
  INV_X1    g069(.A(new_n224), .ZN(new_n256));
  OAI21_X1  g070(.A(G101), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n249), .A2(new_n257), .ZN(new_n258));
  OR2_X1    g072(.A1(new_n254), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n251), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT86), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT86), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n251), .A2(new_n262), .A3(new_n259), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n213), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n213), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(KEYINPUT6), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  AND3_X1   g081(.A1(new_n251), .A2(new_n262), .A3(new_n259), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n262), .B1(new_n251), .B2(new_n259), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n265), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n212), .B1(new_n267), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT7), .B1(new_n209), .B2(G953), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n208), .B(new_n274), .ZN(new_n275));
  XOR2_X1   g089(.A(new_n213), .B(KEYINPUT8), .Z(new_n276));
  NAND2_X1  g090(.A1(new_n254), .A2(new_n258), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n276), .B1(new_n259), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n266), .ZN(new_n280));
  AOI21_X1  g094(.A(G902), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n187), .B1(new_n273), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n271), .B1(new_n270), .B2(new_n280), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n261), .A2(new_n263), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT6), .B1(new_n285), .B2(new_n265), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n211), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n287), .A2(KEYINPUT87), .A3(new_n281), .ZN(new_n288));
  OAI21_X1  g102(.A(G210), .B1(G237), .B2(G902), .ZN(new_n289));
  XOR2_X1   g103(.A(new_n289), .B(KEYINPUT88), .Z(new_n290));
  NAND3_X1  g104(.A1(new_n283), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n287), .A2(new_n281), .A3(new_n289), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT89), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT89), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n287), .A2(new_n294), .A3(new_n281), .A4(new_n289), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n291), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G478), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n297), .A2(KEYINPUT15), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT9), .B(G234), .ZN(new_n299));
  INV_X1    g113(.A(G217), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n299), .A2(new_n300), .A3(G953), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n188), .A2(G128), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n198), .A2(G143), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G134), .ZN(new_n306));
  INV_X1    g120(.A(G134), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n303), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(G116), .B(G122), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n220), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n237), .A2(G122), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(KEYINPUT14), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT94), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT14), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n317), .B1(new_n237), .B2(G122), .ZN(new_n318));
  AOI21_X1  g132(.A(KEYINPUT94), .B1(new_n318), .B2(new_n313), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n316), .B1(new_n319), .B2(new_n314), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n312), .B1(new_n320), .B2(G107), .ZN(new_n321));
  XNOR2_X1  g135(.A(new_n220), .B(new_n310), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n198), .A2(G143), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n323), .B1(KEYINPUT13), .B2(new_n304), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n323), .A2(KEYINPUT13), .ZN(new_n325));
  OAI21_X1  g139(.A(G134), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n322), .A2(new_n326), .A3(new_n308), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n302), .B1(new_n321), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n322), .A2(new_n326), .A3(new_n308), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n320), .A2(G107), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n329), .B(new_n301), .C1(new_n330), .C2(new_n312), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G902), .ZN(new_n333));
  AOI21_X1  g147(.A(KEYINPUT95), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT95), .ZN(new_n335));
  AOI211_X1 g149(.A(new_n335), .B(G902), .C1(new_n328), .C2(new_n331), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n298), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n332), .A2(new_n333), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n337), .B1(new_n339), .B2(new_n298), .ZN(new_n340));
  INV_X1    g154(.A(G953), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT67), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT67), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G953), .ZN(new_n344));
  INV_X1    g158(.A(G237), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n342), .A2(new_n344), .A3(G214), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n188), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT67), .B(G953), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n348), .A2(G143), .A3(G214), .A4(new_n345), .ZN(new_n349));
  NAND2_X1  g163(.A1(KEYINPUT18), .A2(G131), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n350), .B(KEYINPUT90), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n347), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT91), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n347), .A2(new_n349), .A3(KEYINPUT91), .A4(new_n351), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G125), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G140), .ZN(new_n358));
  INV_X1    g172(.A(G140), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G125), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(G146), .ZN(new_n362));
  NOR3_X1   g176(.A1(new_n359), .A2(KEYINPUT72), .A3(G125), .ZN(new_n363));
  XNOR2_X1  g177(.A(G125), .B(G140), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n363), .B1(new_n364), .B2(KEYINPUT72), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n362), .B1(new_n365), .B2(G146), .ZN(new_n366));
  INV_X1    g180(.A(G131), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n367), .B1(new_n347), .B2(new_n349), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n366), .B1(KEYINPUT18), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n356), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(KEYINPUT17), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n347), .A2(new_n349), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G131), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n347), .A2(new_n349), .A3(new_n367), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n371), .B1(new_n375), .B2(KEYINPUT17), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT73), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n360), .A2(KEYINPUT16), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT72), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n379), .A2(new_n357), .A3(G140), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n361), .B2(new_n379), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n378), .B1(new_n381), .B2(KEYINPUT16), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n377), .B1(new_n382), .B2(G146), .ZN(new_n383));
  INV_X1    g197(.A(new_n378), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT16), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n384), .B1(new_n365), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(KEYINPUT73), .A3(new_n190), .ZN(new_n387));
  OAI211_X1 g201(.A(G146), .B(new_n384), .C1(new_n365), .C2(new_n385), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n383), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n370), .B1(new_n376), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(G113), .B(G122), .ZN(new_n391));
  XNOR2_X1  g205(.A(KEYINPUT92), .B(G104), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n391), .B(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n393), .B(new_n370), .C1(new_n376), .C2(new_n389), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n333), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G475), .ZN(new_n399));
  OAI211_X1 g213(.A(KEYINPUT19), .B(new_n380), .C1(new_n361), .C2(new_n379), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT19), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n364), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(new_n190), .A3(new_n402), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n388), .A2(new_n403), .ZN(new_n404));
  AOI22_X1  g218(.A1(new_n356), .A2(new_n369), .B1(new_n404), .B2(new_n375), .ZN(new_n405));
  OAI21_X1  g219(.A(KEYINPUT93), .B1(new_n405), .B2(new_n393), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n404), .A2(new_n375), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n370), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT93), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(new_n394), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n406), .A2(new_n410), .A3(new_n396), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT20), .ZN(new_n412));
  NOR2_X1   g226(.A1(G475), .A2(G902), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n412), .B1(new_n411), .B2(new_n413), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n340), .B(new_n399), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(G234), .A2(G237), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n417), .A2(G952), .A3(new_n341), .ZN(new_n418));
  INV_X1    g232(.A(new_n348), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n419), .A2(G902), .A3(new_n417), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT21), .B(G898), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n418), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n416), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(G214), .B1(G237), .B2(G902), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n296), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n426));
  INV_X1    g240(.A(G137), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G134), .ZN(new_n428));
  NOR2_X1   g242(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n426), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n307), .A2(G137), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n427), .A2(KEYINPUT65), .A3(KEYINPUT11), .A4(G134), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n367), .A2(KEYINPUT66), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  AND4_X1   g248(.A1(new_n430), .A2(new_n431), .A3(new_n432), .A4(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n427), .A2(G134), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n307), .A2(G137), .ZN(new_n437));
  INV_X1    g251(.A(new_n426), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n434), .B1(new_n439), .B2(new_n430), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n194), .A2(new_n196), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(new_n199), .A3(new_n191), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT81), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT81), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n197), .A2(new_n445), .A3(new_n199), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n442), .A2(new_n191), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n189), .A2(G128), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n444), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(new_n258), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n258), .A2(new_n200), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n441), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT83), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT12), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT83), .B1(new_n454), .B2(KEYINPUT12), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n458), .B(new_n459), .C1(new_n457), .C2(new_n455), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT10), .ZN(new_n461));
  NOR3_X1   g275(.A1(new_n258), .A2(new_n200), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n462), .B1(new_n452), .B2(new_n461), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n234), .B(new_n207), .C1(new_n248), .C2(new_n250), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n463), .A2(new_n464), .A3(new_n441), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT82), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT82), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n463), .A2(new_n464), .A3(new_n467), .A4(new_n441), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n460), .A2(new_n469), .ZN(new_n470));
  XOR2_X1   g284(.A(G110), .B(G140), .Z(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(KEYINPUT77), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n348), .A2(G227), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n472), .B(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n474), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n469), .A2(KEYINPUT84), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n463), .A2(new_n464), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n478), .B1(new_n440), .B2(new_n435), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n474), .B1(new_n466), .B2(new_n468), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n481), .A2(KEYINPUT84), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n475), .B(G469), .C1(new_n480), .C2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G469), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n481), .A2(new_n460), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n476), .B1(new_n469), .B2(new_n479), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n484), .B(new_n333), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n484), .A2(new_n333), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n483), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT85), .ZN(new_n491));
  OAI21_X1  g305(.A(G221), .B1(new_n299), .B2(G902), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n491), .B1(new_n490), .B2(new_n492), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g309(.A1(new_n425), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n207), .B1(new_n435), .B2(new_n440), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n448), .A2(new_n206), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n443), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n439), .A2(new_n367), .A3(new_n430), .ZN(new_n500));
  OAI21_X1  g314(.A(G131), .B1(new_n437), .B2(new_n436), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n243), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n497), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT70), .B1(new_n505), .B2(KEYINPUT28), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n503), .B1(new_n497), .B2(new_n502), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT28), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT70), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT28), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n504), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n506), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n348), .A2(G210), .A3(new_n345), .ZN(new_n513));
  XOR2_X1   g327(.A(KEYINPUT26), .B(G101), .Z(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n516));
  XOR2_X1   g330(.A(new_n515), .B(new_n516), .Z(new_n517));
  NAND2_X1  g331(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT30), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n497), .A2(new_n502), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n519), .B1(new_n497), .B2(new_n502), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n243), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT69), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n515), .B(new_n516), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n522), .A2(new_n523), .A3(new_n524), .A4(new_n504), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT31), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n518), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(G472), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n529), .A2(KEYINPUT32), .A3(new_n530), .A4(new_n333), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT71), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n529), .A2(new_n530), .A3(new_n333), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT32), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n497), .A2(new_n502), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT30), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n497), .A2(new_n502), .A3(new_n519), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n505), .B1(new_n539), .B2(new_n243), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n540), .A2(new_n523), .A3(KEYINPUT31), .A4(new_n524), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n525), .A2(new_n526), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(G902), .B1(new_n543), .B2(new_n518), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT71), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n544), .A2(new_n545), .A3(KEYINPUT32), .A4(new_n530), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n508), .A2(new_n511), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n547), .A2(KEYINPUT29), .A3(new_n524), .A4(new_n506), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n512), .A2(new_n517), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT29), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n550), .B1(new_n540), .B2(new_n524), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n548), .B(new_n333), .C1(new_n549), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(G472), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n532), .A2(new_n535), .A3(new_n546), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n198), .A2(G119), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n235), .A2(G128), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT24), .B(G110), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT23), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n198), .A2(KEYINPUT23), .A3(G119), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(new_n562), .A3(new_n556), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n559), .B1(new_n563), .B2(G110), .ZN(new_n564));
  XOR2_X1   g378(.A(new_n564), .B(KEYINPUT75), .Z(new_n565));
  OAI211_X1 g379(.A(new_n565), .B(new_n388), .C1(G146), .C2(new_n361), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT74), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n557), .A2(new_n558), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n568), .B1(G110), .B2(new_n563), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n389), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n567), .B1(new_n389), .B2(new_n569), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n566), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n348), .A2(G221), .A3(G234), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT22), .B(G137), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n575), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n566), .B(new_n577), .C1(new_n570), .C2(new_n571), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(KEYINPUT25), .B1(new_n579), .B2(new_n333), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT25), .ZN(new_n581));
  AOI211_X1 g395(.A(new_n581), .B(G902), .C1(new_n576), .C2(new_n578), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n300), .B1(G234), .B2(new_n333), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT76), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n579), .A2(new_n333), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n585), .B1(new_n586), .B2(new_n584), .ZN(new_n587));
  INV_X1    g401(.A(new_n584), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n579), .A2(KEYINPUT76), .A3(new_n333), .A4(new_n588), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n583), .A2(new_n584), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n554), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n496), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(G101), .ZN(G3));
  NAND2_X1  g407(.A1(new_n490), .A2(new_n492), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT85), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n587), .A2(new_n589), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n584), .B1(new_n580), .B2(new_n582), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n529), .A2(new_n333), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G472), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n533), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n595), .A2(new_n596), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n424), .ZN(new_n605));
  INV_X1    g419(.A(new_n289), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n606), .B1(new_n273), .B2(new_n282), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n605), .B1(new_n607), .B2(new_n292), .ZN(new_n608));
  INV_X1    g422(.A(new_n422), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n399), .B1(new_n414), .B2(new_n415), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n297), .A2(G902), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT96), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n328), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT33), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n328), .A2(new_n331), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n614), .A2(new_n615), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n611), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OR3_X1    g433(.A1(new_n334), .A2(new_n336), .A3(G478), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n610), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n608), .A2(new_n609), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n604), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT34), .B(G104), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  OAI21_X1  g441(.A(new_n338), .B1(KEYINPUT15), .B2(new_n297), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n337), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n629), .B(new_n399), .C1(new_n415), .C2(new_n414), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT97), .B1(new_n630), .B2(new_n422), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n411), .A2(new_n413), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(KEYINPUT20), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n634));
  AOI22_X1  g448(.A1(new_n633), .A2(new_n634), .B1(G475), .B2(new_n398), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT97), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n635), .A2(new_n636), .A3(new_n609), .A4(new_n629), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n608), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n638), .A2(new_n608), .A3(KEYINPUT98), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n604), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT35), .B(G107), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  NOR2_X1   g459(.A1(new_n577), .A2(KEYINPUT36), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n572), .B(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(new_n333), .A3(new_n588), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n598), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(new_n602), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n496), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT99), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  NAND2_X1  g469(.A1(new_n633), .A2(new_n634), .ZN(new_n656));
  INV_X1    g470(.A(G900), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n418), .B1(new_n420), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n656), .A2(new_n399), .A3(new_n629), .A4(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n598), .B2(new_n648), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n554), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n662), .A2(new_n595), .A3(new_n596), .A4(new_n608), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  XNOR2_X1  g478(.A(new_n296), .B(KEYINPUT38), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n517), .B1(new_n505), .B2(new_n507), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n666), .A2(KEYINPUT100), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n540), .A2(new_n524), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n666), .A2(KEYINPUT100), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(G902), .B1(new_n670), .B2(KEYINPUT101), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n671), .B1(KEYINPUT101), .B2(new_n670), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(G472), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n673), .A2(new_n532), .A3(new_n546), .A4(new_n535), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT102), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n610), .A2(new_n629), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n649), .A2(new_n605), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n665), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n658), .B(KEYINPUT39), .Z(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n493), .A2(new_n494), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(KEYINPUT40), .ZN(new_n683));
  OR2_X1    g497(.A1(new_n682), .A2(KEYINPUT40), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n679), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(new_n188), .ZN(G45));
  NAND3_X1  g500(.A1(new_n610), .A2(new_n621), .A3(new_n659), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n598), .B2(new_n648), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n554), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n689), .A2(new_n595), .A3(new_n596), .A4(new_n608), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G146), .ZN(G48));
  NAND2_X1  g505(.A1(new_n469), .A2(new_n479), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n474), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n481), .A2(new_n460), .ZN(new_n694));
  AOI21_X1  g508(.A(G902), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(KEYINPUT103), .A2(G469), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI22_X1  g511(.A1(new_n692), .A2(new_n474), .B1(new_n481), .B2(new_n460), .ZN(new_n698));
  OAI211_X1 g512(.A(KEYINPUT103), .B(G469), .C1(new_n698), .C2(G902), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n697), .A2(new_n699), .A3(new_n492), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(new_n554), .A3(new_n590), .ZN(new_n701));
  OR3_X1    g515(.A1(new_n701), .A2(new_n624), .A3(KEYINPUT104), .ZN(new_n702));
  OAI21_X1  g516(.A(KEYINPUT104), .B1(new_n701), .B2(new_n624), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(KEYINPUT41), .B(G113), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G15));
  AOI21_X1  g520(.A(new_n701), .B1(new_n641), .B2(new_n642), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n237), .ZN(G18));
  AND2_X1   g522(.A1(new_n649), .A2(new_n423), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n709), .A2(new_n554), .A3(new_n608), .A4(new_n700), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G119), .ZN(G21));
  NAND3_X1  g525(.A1(new_n600), .A2(KEYINPUT106), .A3(G472), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n713), .B1(new_n544), .B2(new_n530), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n547), .A2(KEYINPUT105), .A3(new_n506), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n512), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n524), .B1(new_n715), .B2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n543), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n530), .B(new_n333), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n712), .A2(new_n714), .A3(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n599), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n697), .A2(new_n699), .A3(new_n492), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n422), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  AOI211_X1 g539(.A(new_n605), .B(new_n677), .C1(new_n607), .C2(new_n292), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  XOR2_X1   g542(.A(new_n728), .B(G122), .Z(G24));
  NOR3_X1   g543(.A1(new_n650), .A2(new_n721), .A3(new_n687), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n608), .A3(new_n700), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G125), .ZN(G27));
  AND2_X1   g546(.A1(new_n293), .A2(new_n295), .ZN(new_n733));
  INV_X1    g547(.A(new_n492), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n488), .B1(new_n695), .B2(new_n484), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n734), .B1(new_n735), .B2(new_n483), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n733), .A2(new_n736), .A3(new_n424), .A4(new_n291), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n535), .A2(new_n553), .A3(new_n531), .ZN(new_n738));
  INV_X1    g552(.A(new_n687), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n590), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  OAI21_X1  g554(.A(KEYINPUT42), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  AND4_X1   g555(.A1(new_n424), .A2(new_n291), .A3(new_n293), .A4(new_n295), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n687), .A2(KEYINPUT42), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n742), .A2(new_n591), .A3(new_n736), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n367), .ZN(G33));
  INV_X1    g560(.A(new_n660), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n742), .A2(new_n591), .A3(new_n736), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G134), .ZN(G36));
  NAND2_X1  g563(.A1(new_n635), .A2(new_n621), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT43), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n635), .A2(new_n753), .A3(new_n621), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n751), .A2(new_n752), .A3(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n752), .B1(new_n751), .B2(new_n754), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n602), .B(new_n649), .C1(new_n756), .C2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  AND3_X1   g573(.A1(new_n758), .A2(KEYINPUT110), .A3(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(KEYINPUT110), .B1(new_n758), .B2(new_n759), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n742), .B1(new_n758), .B2(new_n759), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XOR2_X1   g578(.A(KEYINPUT107), .B(KEYINPUT108), .Z(new_n765));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n475), .B1(new_n480), .B2(new_n482), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(KEYINPUT45), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n766), .B(G469), .C1(new_n768), .C2(G902), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n767), .A2(KEYINPUT45), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n767), .A2(KEYINPUT45), .ZN(new_n771));
  OAI21_X1  g585(.A(G469), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(KEYINPUT46), .A3(new_n489), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n769), .A2(new_n773), .A3(new_n487), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n492), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n765), .B1(new_n775), .B2(new_n681), .ZN(new_n776));
  INV_X1    g590(.A(new_n765), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n774), .A2(new_n492), .A3(new_n680), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n764), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G137), .ZN(G39));
  NAND4_X1  g595(.A1(new_n291), .A2(new_n424), .A3(new_n293), .A4(new_n295), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n782), .A2(new_n554), .A3(new_n590), .A4(new_n687), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n774), .A2(KEYINPUT47), .A3(new_n492), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT47), .B1(new_n774), .B2(new_n492), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n783), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  NAND2_X1  g602(.A1(new_n697), .A2(new_n699), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT49), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n492), .A2(new_n424), .ZN(new_n791));
  NOR4_X1   g605(.A1(new_n790), .A2(new_n599), .A3(new_n750), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n296), .A2(KEYINPUT38), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n296), .A2(KEYINPUT38), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n674), .B(KEYINPUT102), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n792), .A2(new_n793), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n751), .A2(new_n418), .A3(new_n754), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n797), .A2(new_n599), .A3(new_n721), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(new_n608), .A3(new_n700), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(G952), .A3(new_n341), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n782), .A2(new_n723), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n590), .A2(new_n418), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n795), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n800), .B1(new_n803), .B2(new_n623), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT48), .ZN(new_n805));
  INV_X1    g619(.A(new_n797), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n801), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT114), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n801), .A2(new_n809), .A3(new_n806), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n590), .A2(new_n738), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n805), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  AOI211_X1 g628(.A(KEYINPUT48), .B(new_n812), .C1(new_n808), .C2(new_n810), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n804), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n650), .A2(new_n721), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n811), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n723), .A2(new_n424), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n798), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n820), .A2(KEYINPUT50), .A3(new_n793), .A4(new_n794), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT50), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n798), .A2(new_n819), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n822), .B1(new_n665), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n621), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n803), .A2(new_n635), .A3(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n818), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT47), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n775), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n697), .A2(new_n699), .A3(new_n734), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n830), .A2(new_n784), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n742), .A3(new_n798), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n828), .A2(new_n833), .A3(KEYINPUT51), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT116), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n828), .A2(new_n833), .A3(KEYINPUT116), .A4(KEYINPUT51), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n816), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n798), .A2(new_n742), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n785), .A2(new_n786), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n840), .B1(new_n841), .B2(new_n831), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n818), .A2(new_n827), .A3(new_n825), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n839), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT115), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT115), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n846), .B(new_n839), .C1(new_n842), .C2(new_n843), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n838), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n849), .B1(new_n838), .B2(new_n848), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n649), .A2(new_n658), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n726), .A2(new_n674), .A3(new_n736), .A4(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n663), .A2(new_n690), .A3(new_n731), .A4(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT52), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT112), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n854), .A2(new_n855), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n854), .A2(KEYINPUT112), .A3(new_n855), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n710), .B1(new_n725), .B2(new_n727), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n707), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n622), .A2(new_n630), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n296), .A2(new_n609), .A3(new_n424), .A4(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n865), .A2(new_n604), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n425), .B(new_n495), .C1(new_n591), .C2(new_n651), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n863), .A2(new_n704), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT111), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(new_n416), .B2(new_n658), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n635), .A2(KEYINPUT111), .A3(new_n340), .A4(new_n659), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n554), .A2(new_n873), .A3(new_n649), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n874), .A2(new_n493), .A3(new_n494), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n782), .A2(new_n594), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n875), .A2(new_n742), .B1(new_n876), .B2(new_n730), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n877), .A2(new_n741), .A3(new_n744), .A4(new_n748), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n869), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n861), .A2(KEYINPUT53), .A3(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n881));
  INV_X1    g695(.A(new_n874), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n495), .A2(new_n882), .A3(new_n742), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n742), .A2(new_n736), .A3(new_n730), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n748), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(new_n745), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n866), .A2(new_n707), .A3(new_n862), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n886), .A2(new_n704), .A3(new_n887), .A4(new_n868), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n854), .B(KEYINPUT52), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n881), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT113), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n880), .A2(new_n890), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n861), .A2(new_n881), .A3(new_n879), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT53), .B1(new_n888), .B2(new_n889), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n894), .A2(new_n895), .A3(KEYINPUT54), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n880), .A2(new_n890), .A3(new_n892), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT113), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n850), .A2(new_n851), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(G952), .A2(G953), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n796), .B1(new_n901), .B2(new_n902), .ZN(G75));
  NOR2_X1   g717(.A1(new_n348), .A2(G952), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n284), .A2(new_n286), .A3(new_n211), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n273), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT55), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n333), .B1(new_n880), .B2(new_n890), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n606), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT56), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n907), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n908), .A2(new_n290), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n907), .A2(new_n910), .ZN(new_n913));
  AOI211_X1 g727(.A(new_n904), .B(new_n911), .C1(new_n912), .C2(new_n913), .ZN(G51));
  XNOR2_X1  g728(.A(new_n488), .B(KEYINPUT57), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n892), .B1(new_n880), .B2(new_n890), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n916), .A2(KEYINPUT118), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n898), .B1(new_n916), .B2(KEYINPUT118), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n486), .B2(new_n485), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n908), .A2(G469), .A3(new_n768), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n904), .B1(new_n920), .B2(new_n921), .ZN(G54));
  INV_X1    g736(.A(new_n904), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n908), .A2(KEYINPUT58), .A3(G475), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(new_n411), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n411), .B2(new_n924), .ZN(G60));
  XNOR2_X1  g740(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n927));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n929), .B1(new_n897), .B2(new_n899), .ZN(new_n930));
  OR2_X1    g744(.A1(new_n617), .A2(new_n618), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n923), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n931), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(new_n929), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(new_n917), .B2(new_n918), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT120), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI211_X1 g751(.A(KEYINPUT120), .B(new_n934), .C1(new_n917), .C2(new_n918), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n932), .B1(new_n937), .B2(new_n938), .ZN(G63));
  NAND2_X1  g753(.A1(new_n880), .A2(new_n890), .ZN(new_n940));
  NAND2_X1  g754(.A1(G217), .A2(G902), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT60), .Z(new_n942));
  NAND3_X1  g756(.A1(new_n940), .A2(new_n647), .A3(new_n942), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n940), .A2(new_n942), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n923), .B(new_n943), .C1(new_n944), .C2(new_n579), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g760(.A(G953), .B1(new_n421), .B2(new_n209), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT122), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT121), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n869), .B(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n948), .B1(new_n950), .B2(new_n419), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n267), .B(new_n272), .C1(G898), .C2(new_n348), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n951), .B(new_n952), .ZN(G69));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n419), .A2(new_n657), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT124), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n779), .A2(new_n726), .A3(new_n813), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n663), .A2(new_n690), .A3(new_n731), .ZN(new_n958));
  INV_X1    g772(.A(new_n748), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n745), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n780), .A2(new_n957), .A3(new_n787), .A4(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n956), .B1(new_n961), .B2(new_n348), .ZN(new_n962));
  AND4_X1   g776(.A1(new_n591), .A2(new_n682), .A3(new_n742), .A4(new_n864), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT62), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n685), .B2(new_n958), .ZN(new_n965));
  INV_X1    g779(.A(new_n958), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n684), .A2(new_n683), .ZN(new_n967));
  OAI211_X1 g781(.A(KEYINPUT62), .B(new_n966), .C1(new_n967), .C2(new_n679), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n963), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n841), .ZN(new_n970));
  AOI22_X1  g784(.A1(new_n970), .A2(new_n783), .B1(new_n764), .B2(new_n779), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n419), .B1(new_n969), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n400), .A2(new_n402), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n539), .B(new_n973), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n974), .A2(KEYINPUT123), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n962), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n974), .B1(new_n972), .B2(KEYINPUT123), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n348), .B1(G227), .B2(G900), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n954), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  AOI211_X1 g795(.A(KEYINPUT125), .B(new_n979), .C1(new_n976), .C2(new_n977), .ZN(new_n982));
  OAI22_X1  g796(.A1(new_n981), .A2(new_n982), .B1(new_n980), .B2(new_n978), .ZN(G72));
  NAND2_X1  g797(.A1(G472), .A2(G902), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT63), .Z(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT126), .Z(new_n986));
  INV_X1    g800(.A(new_n950), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n986), .B1(new_n961), .B2(new_n987), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n988), .A2(new_n517), .A3(new_n540), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n969), .A2(new_n950), .A3(new_n971), .ZN(new_n990));
  AOI211_X1 g804(.A(new_n517), .B(new_n540), .C1(new_n990), .C2(new_n986), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n540), .B(new_n524), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n985), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT127), .Z(new_n994));
  AND3_X1   g808(.A1(new_n894), .A2(new_n895), .A3(new_n994), .ZN(new_n995));
  NOR4_X1   g809(.A1(new_n989), .A2(new_n991), .A3(new_n904), .A4(new_n995), .ZN(G57));
endmodule


