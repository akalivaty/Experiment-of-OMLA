//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G125), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G140), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n192), .A2(new_n194), .A3(new_n195), .ZN(new_n196));
  OR2_X1    g010(.A1(new_n196), .A2(KEYINPUT78), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(KEYINPUT78), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT16), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(new_n191), .A3(G125), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n192), .A2(new_n194), .ZN(new_n202));
  OAI211_X1 g016(.A(G146), .B(new_n201), .C1(new_n202), .C2(new_n200), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n205));
  INV_X1    g019(.A(G119), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n206), .B2(G128), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(G128), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT23), .A3(G119), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G110), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT76), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(G119), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n208), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT24), .B(G110), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n212), .A2(KEYINPUT76), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT77), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g034(.A1(new_n212), .A2(KEYINPUT76), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT77), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n221), .A2(new_n222), .A3(new_n217), .A4(new_n213), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n204), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n201), .B1(new_n202), .B2(new_n200), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(new_n195), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n203), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n215), .A2(new_n216), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n229), .B1(G110), .B2(new_n211), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(KEYINPUT72), .B(G953), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(G221), .A3(G234), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT22), .B(G137), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n233), .B(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n225), .A2(new_n231), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n235), .ZN(new_n237));
  INV_X1    g051(.A(new_n231), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n237), .B1(new_n224), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n188), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n236), .A2(KEYINPUT25), .A3(new_n239), .A4(new_n188), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n190), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n236), .A2(new_n239), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n189), .A2(G902), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n245), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT32), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT74), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n254));
  INV_X1    g068(.A(G137), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n253), .A2(new_n254), .A3(new_n255), .A4(G134), .ZN(new_n256));
  INV_X1    g070(.A(G134), .ZN(new_n257));
  OAI22_X1  g071(.A1(new_n257), .A2(G137), .B1(KEYINPUT66), .B2(KEYINPUT11), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G131), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n257), .A2(G137), .B1(KEYINPUT66), .B2(KEYINPUT11), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n257), .A2(G137), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n255), .A2(G134), .ZN(new_n264));
  OAI21_X1  g078(.A(G131), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G143), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT64), .B1(new_n267), .B2(G146), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT64), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(new_n195), .A3(G143), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n267), .A2(G146), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n268), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n267), .A2(G146), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT1), .ZN(new_n274));
  OAI21_X1  g088(.A(G128), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(G143), .B(G146), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n272), .A2(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n266), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n259), .A2(new_n261), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G131), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n262), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n195), .A2(G143), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n283), .A2(new_n271), .A3(KEYINPUT0), .A4(G128), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT65), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT65), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n276), .A2(new_n286), .A3(KEYINPUT0), .A4(G128), .ZN(new_n287));
  XOR2_X1   g101(.A(KEYINPUT0), .B(G128), .Z(new_n288));
  AOI22_X1  g102(.A1(new_n285), .A2(new_n287), .B1(new_n272), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n279), .B1(new_n282), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT71), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT70), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n292), .B1(new_n206), .B2(G116), .ZN(new_n293));
  INV_X1    g107(.A(G116), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(KEYINPUT70), .A3(G119), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n206), .A2(G116), .ZN(new_n297));
  INV_X1    g111(.A(G113), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT2), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT2), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G113), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n296), .A2(new_n297), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n302), .B1(new_n296), .B2(new_n297), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n291), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n294), .A2(KEYINPUT70), .A3(G119), .ZN(new_n306));
  AOI21_X1  g120(.A(KEYINPUT70), .B1(new_n294), .B2(G119), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n297), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n302), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n296), .A2(new_n297), .A3(new_n302), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(KEYINPUT71), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n305), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n290), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT28), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n313), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n272), .A2(new_n275), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n277), .A2(new_n283), .A3(new_n271), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n262), .A2(KEYINPUT67), .A3(new_n265), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT67), .B1(new_n262), .B2(new_n265), .ZN(new_n323));
  OAI211_X1 g137(.A(KEYINPUT68), .B(new_n321), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n282), .A2(new_n289), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT67), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n266), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n262), .A2(KEYINPUT67), .A3(new_n265), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT68), .B1(new_n330), .B2(new_n321), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n318), .B1(new_n326), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT73), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n333), .B1(new_n290), .B2(new_n313), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n315), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n333), .B(new_n318), .C1(new_n326), .C2(new_n331), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n317), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G237), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n232), .A2(G210), .A3(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(KEYINPUT27), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT26), .B(G101), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n340), .B(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n252), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n324), .A2(new_n325), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n330), .A2(new_n321), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT68), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n313), .B1(new_n344), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n334), .ZN(new_n349));
  OAI211_X1 g163(.A(KEYINPUT28), .B(new_n336), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n316), .ZN(new_n351));
  INV_X1    g165(.A(new_n342), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(KEYINPUT74), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n343), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT30), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(new_n326), .B2(new_n331), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT69), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n290), .A2(KEYINPUT30), .ZN(new_n359));
  OAI211_X1 g173(.A(KEYINPUT69), .B(new_n355), .C1(new_n326), .C2(new_n331), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n358), .A2(new_n318), .A3(new_n359), .A4(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(new_n342), .A3(new_n314), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT31), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n361), .A2(KEYINPUT31), .A3(new_n342), .A4(new_n314), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n354), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(G472), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n188), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n251), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n368), .A2(new_n251), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n343), .A2(new_n353), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n364), .A2(new_n365), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT29), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n361), .A2(new_n352), .A3(new_n314), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n352), .B1(new_n350), .B2(new_n316), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OR2_X1    g192(.A1(new_n290), .A2(new_n313), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n315), .B1(new_n379), .B2(new_n314), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT75), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n316), .A2(KEYINPUT75), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n382), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n352), .A2(new_n375), .ZN(new_n385));
  AOI21_X1  g199(.A(G902), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n367), .B1(new_n378), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n374), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n250), .B1(new_n369), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(G214), .B1(G237), .B2(G902), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(KEYINPUT81), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(G110), .B(G122), .ZN(new_n393));
  INV_X1    g207(.A(G104), .ZN(new_n394));
  OAI21_X1  g208(.A(KEYINPUT3), .B1(new_n394), .B2(G107), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n396));
  INV_X1    g210(.A(G107), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(G104), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(G107), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n395), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n400), .A2(new_n401), .A3(G101), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(G101), .ZN(new_n403));
  INV_X1    g217(.A(G101), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n395), .A2(new_n398), .A3(new_n404), .A4(new_n399), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(KEYINPUT4), .A3(new_n405), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n305), .A2(new_n312), .A3(new_n402), .A4(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n296), .A2(KEYINPUT5), .A3(new_n297), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n408), .B(G113), .C1(KEYINPUT5), .C2(new_n297), .ZN(new_n409));
  OAI21_X1  g223(.A(KEYINPUT79), .B1(new_n394), .B2(G107), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT79), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(new_n397), .A3(G104), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n412), .A3(new_n399), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G101), .ZN(new_n414));
  AND2_X1   g228(.A1(new_n414), .A2(new_n405), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n409), .A2(new_n415), .A3(new_n311), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n393), .B1(new_n407), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT6), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT6), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n407), .A2(new_n393), .A3(new_n416), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT82), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT82), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n407), .A2(new_n422), .A3(new_n393), .A4(new_n416), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n419), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n418), .B1(new_n424), .B2(new_n417), .ZN(new_n425));
  OR3_X1    g239(.A1(new_n321), .A2(KEYINPUT83), .A3(G125), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT83), .B1(new_n321), .B2(G125), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n289), .A2(new_n193), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G224), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(G953), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n431), .B(KEYINPUT84), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n429), .B(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n425), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G210), .B1(G237), .B2(G902), .ZN(new_n435));
  XOR2_X1   g249(.A(new_n393), .B(KEYINPUT8), .Z(new_n436));
  NAND2_X1  g250(.A1(new_n409), .A2(new_n311), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n414), .A2(new_n405), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n436), .B1(new_n439), .B2(new_n416), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT7), .B1(new_n430), .B2(G953), .ZN(new_n441));
  OR2_X1    g255(.A1(new_n429), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n429), .A2(new_n441), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n440), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n421), .A2(new_n423), .ZN(new_n445));
  AOI21_X1  g259(.A(G902), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n434), .A2(new_n435), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n435), .B1(new_n434), .B2(new_n446), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n392), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT85), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n434), .A2(new_n446), .ZN(new_n452));
  INV_X1    g266(.A(new_n435), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n434), .A2(new_n435), .A3(new_n446), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(KEYINPUT85), .A3(new_n392), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT9), .B(G234), .ZN(new_n458));
  OAI21_X1  g272(.A(G221), .B1(new_n458), .B2(G902), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G469), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n415), .A2(KEYINPUT10), .A3(new_n321), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n289), .A2(new_n402), .A3(new_n406), .ZN(new_n463));
  INV_X1    g277(.A(new_n282), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n209), .B1(new_n283), .B2(KEYINPUT1), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n320), .B1(new_n465), .B2(new_n276), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n414), .A3(new_n405), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT10), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n462), .A2(new_n463), .A3(new_n464), .A4(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n232), .A2(G227), .ZN(new_n471));
  XOR2_X1   g285(.A(G110), .B(G140), .Z(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT12), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT80), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n438), .A2(new_n477), .A3(new_n278), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n477), .B1(new_n438), .B2(new_n278), .ZN(new_n479));
  INV_X1    g293(.A(new_n467), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n476), .B1(new_n481), .B2(new_n464), .ZN(new_n482));
  INV_X1    g296(.A(new_n479), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n438), .A2(new_n477), .A3(new_n278), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n467), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(KEYINPUT12), .A3(new_n282), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n475), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n462), .A2(new_n463), .A3(new_n469), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n282), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n474), .B1(new_n489), .B2(new_n470), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n461), .B(new_n188), .C1(new_n487), .C2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n461), .A2(new_n188), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n475), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n489), .ZN(new_n496));
  INV_X1    g310(.A(new_n470), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n497), .B1(new_n482), .B2(new_n486), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n496), .B(G469), .C1(new_n498), .C2(new_n474), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n460), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n451), .A2(new_n457), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(G953), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT72), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT72), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G953), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n503), .A2(new_n505), .A3(G214), .A4(new_n338), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n267), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n232), .A2(G143), .A3(G214), .A4(new_n338), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(G131), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT17), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n507), .A2(new_n508), .A3(new_n260), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT89), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT88), .ZN(new_n516));
  AOI211_X1 g330(.A(new_n511), .B(new_n260), .C1(new_n507), .C2(new_n508), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n516), .B1(new_n517), .B2(new_n228), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n509), .A2(KEYINPUT17), .A3(G131), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n519), .A2(KEYINPUT88), .A3(new_n203), .A4(new_n227), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n510), .A2(KEYINPUT89), .A3(new_n511), .A4(new_n512), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n515), .A2(new_n518), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n509), .A2(KEYINPUT18), .A3(G131), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n509), .B1(KEYINPUT18), .B2(G131), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n197), .A2(new_n198), .B1(G146), .B2(new_n202), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(G113), .B(G122), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT87), .B(G104), .ZN(new_n529));
  XOR2_X1   g343(.A(new_n528), .B(new_n529), .Z(new_n530));
  NAND3_X1  g344(.A1(new_n522), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n530), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n202), .B(KEYINPUT19), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n203), .B1(new_n533), .B2(G146), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n534), .B1(new_n510), .B2(new_n512), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n532), .B1(new_n526), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT20), .ZN(new_n538));
  NOR2_X1   g352(.A1(G475), .A2(G902), .ZN(new_n539));
  XOR2_X1   g353(.A(new_n539), .B(KEYINPUT90), .Z(new_n540));
  NAND3_X1  g354(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT91), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT91), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n537), .A2(new_n543), .A3(new_n538), .A4(new_n540), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n537), .A2(new_n540), .ZN(new_n545));
  XOR2_X1   g359(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n542), .A2(new_n544), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n531), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n530), .B1(new_n522), .B2(new_n527), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n188), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(G475), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT92), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n549), .A2(KEYINPUT92), .A3(new_n553), .ZN(new_n557));
  INV_X1    g371(.A(new_n232), .ZN(new_n558));
  NAND2_X1  g372(.A1(G234), .A2(G237), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n558), .A2(G902), .A3(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT21), .B(G898), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n559), .A2(G952), .A3(new_n502), .ZN(new_n563));
  OR2_X1    g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(G128), .B(G143), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT13), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n209), .A2(KEYINPUT13), .A3(G143), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(new_n257), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n565), .A2(new_n257), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT94), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n566), .A2(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n565), .A2(KEYINPUT94), .A3(new_n257), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n294), .A2(G122), .ZN(new_n573));
  INV_X1    g387(.A(G122), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G116), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT93), .ZN(new_n577));
  XNOR2_X1  g391(.A(G116), .B(G122), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT93), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n577), .A2(new_n580), .A3(G107), .ZN(new_n581));
  AOI21_X1  g395(.A(G107), .B1(new_n577), .B2(new_n580), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n571), .B(new_n572), .C1(new_n581), .C2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n576), .A2(KEYINPUT93), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n578), .A2(new_n579), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n397), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n565), .B(new_n257), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT14), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n578), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT95), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n574), .A2(G116), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n397), .B1(new_n591), .B2(KEYINPUT14), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n589), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n590), .B1(new_n589), .B2(new_n592), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n586), .B(new_n587), .C1(new_n593), .C2(new_n594), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n458), .A2(new_n187), .A3(G953), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n583), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT96), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n583), .A2(new_n595), .ZN(new_n600));
  INV_X1    g414(.A(new_n596), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g416(.A1(new_n583), .A2(new_n595), .A3(KEYINPUT96), .A4(new_n596), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n599), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(G478), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n605), .A2(KEYINPUT15), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n604), .A2(new_n188), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n606), .B1(new_n604), .B2(new_n188), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n556), .A2(new_n557), .A3(new_n564), .A4(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n501), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n389), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(G101), .ZN(G3));
  NAND2_X1  g427(.A1(new_n372), .A2(new_n373), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n367), .B1(new_n614), .B2(new_n188), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n368), .B1(new_n372), .B2(new_n373), .ZN(new_n616));
  INV_X1    g430(.A(new_n500), .ZN(new_n617));
  NOR4_X1   g431(.A1(new_n615), .A2(new_n616), .A3(new_n250), .A4(new_n617), .ZN(new_n618));
  OR2_X1    g432(.A1(new_n604), .A2(KEYINPUT33), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT97), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n602), .B1(new_n620), .B2(new_n597), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n597), .A2(new_n620), .ZN(new_n622));
  OAI21_X1  g436(.A(KEYINPUT33), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n605), .A2(G902), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n604), .A2(new_n188), .ZN(new_n626));
  AOI22_X1  g440(.A1(new_n624), .A2(new_n625), .B1(new_n605), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n557), .ZN(new_n629));
  AOI21_X1  g443(.A(KEYINPUT92), .B1(new_n549), .B2(new_n553), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n628), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n391), .B1(new_n454), .B2(new_n455), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n564), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n618), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT34), .B(G104), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  INV_X1    g451(.A(KEYINPUT98), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n552), .A2(new_n638), .A3(G475), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n638), .B1(new_n552), .B2(G475), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n537), .A2(new_n540), .A3(new_n546), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n609), .B1(new_n548), .B2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(new_n564), .B(KEYINPUT99), .Z(new_n644));
  AND4_X1   g458(.A1(new_n632), .A2(new_n641), .A3(new_n643), .A4(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n618), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT35), .B(G107), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  NOR2_X1   g462(.A1(new_n615), .A2(new_n616), .ZN(new_n649));
  OR4_X1    g463(.A1(KEYINPUT36), .A2(new_n224), .A3(new_n238), .A4(new_n237), .ZN(new_n650));
  OAI22_X1  g464(.A1(new_n224), .A2(new_n238), .B1(KEYINPUT36), .B2(new_n237), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n650), .A2(new_n248), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n244), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n611), .A2(new_n649), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  NAND2_X1  g471(.A1(new_n553), .A2(KEYINPUT98), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n552), .A2(new_n638), .A3(G475), .ZN(new_n659));
  INV_X1    g473(.A(G900), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n563), .B1(new_n560), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n643), .A2(new_n658), .A3(new_n659), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT100), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT100), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n641), .A2(new_n665), .A3(new_n643), .A4(new_n662), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n664), .A2(new_n666), .A3(new_n632), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n664), .A2(new_n666), .A3(KEYINPUT101), .A4(new_n632), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n654), .A2(new_n500), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n369), .B2(new_n388), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G128), .ZN(G30));
  NAND2_X1  g489(.A1(new_n379), .A2(new_n314), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n352), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n362), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT102), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n188), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n678), .A2(KEYINPUT102), .ZN(new_n681));
  OAI21_X1  g495(.A(G472), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n614), .A2(new_n370), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n682), .B(new_n683), .C1(KEYINPUT32), .C2(new_n616), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n629), .A2(new_n630), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n456), .B(KEYINPUT38), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n609), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n653), .A2(new_n689), .A3(new_n392), .ZN(new_n690));
  NOR4_X1   g504(.A1(new_n685), .A2(new_n686), .A3(new_n688), .A4(new_n690), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n691), .A2(KEYINPUT103), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(KEYINPUT103), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n661), .B(KEYINPUT39), .Z(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n617), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT40), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n692), .A2(new_n693), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G143), .ZN(G45));
  OAI211_X1 g513(.A(new_n628), .B(new_n662), .C1(new_n629), .C2(new_n630), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n700), .A2(new_n449), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n673), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G146), .ZN(G48));
  NAND2_X1  g517(.A1(new_n378), .A2(new_n386), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G472), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n683), .B(new_n705), .C1(KEYINPUT32), .C2(new_n616), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n482), .A2(new_n486), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n490), .B1(new_n707), .B2(new_n495), .ZN(new_n708));
  OAI21_X1  g522(.A(G469), .B1(new_n708), .B2(G902), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n709), .A2(new_n459), .A3(new_n491), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n250), .A2(new_n711), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n706), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n634), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  NAND2_X1  g530(.A1(new_n713), .A2(new_n645), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G116), .ZN(G18));
  OAI211_X1 g532(.A(new_n710), .B(new_n392), .C1(new_n447), .C2(new_n448), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(KEYINPUT104), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n456), .A2(new_n721), .A3(new_n392), .A4(new_n710), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n720), .A2(new_n654), .A3(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n610), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n723), .A2(new_n706), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  OR2_X1    g540(.A1(new_n384), .A2(new_n342), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n368), .B1(new_n373), .B2(new_n727), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n615), .A2(new_n250), .A3(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n456), .A2(new_n689), .A3(new_n392), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n710), .A2(new_n644), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n686), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G122), .ZN(G24));
  NOR2_X1   g548(.A1(new_n615), .A2(new_n728), .ZN(new_n735));
  INV_X1    g549(.A(new_n700), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n723), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G125), .ZN(G27));
  OAI21_X1  g552(.A(KEYINPUT107), .B1(KEYINPUT106), .B2(KEYINPUT42), .ZN(new_n739));
  INV_X1    g553(.A(new_n250), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n683), .A2(new_n705), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n616), .A2(KEYINPUT32), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n740), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n627), .B1(new_n556), .B2(new_n557), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n454), .A2(new_n392), .A3(new_n455), .ZN(new_n745));
  INV_X1    g559(.A(new_n493), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n491), .B(new_n746), .C1(new_n499), .C2(new_n747), .ZN(new_n748));
  AND2_X1   g562(.A1(new_n499), .A2(new_n747), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n459), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n744), .A2(new_n662), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n739), .B1(new_n743), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n739), .B1(KEYINPUT107), .B2(KEYINPUT42), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n389), .A2(new_n736), .A3(new_n751), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G131), .ZN(G33));
  AND3_X1   g571(.A1(new_n751), .A2(new_n666), .A3(new_n664), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n706), .A2(new_n758), .A3(new_n740), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G134), .ZN(G36));
  OAI21_X1  g574(.A(new_n496), .B1(new_n498), .B2(new_n474), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XOR2_X1   g577(.A(new_n763), .B(KEYINPUT108), .Z(new_n764));
  AOI21_X1  g578(.A(new_n461), .B1(new_n761), .B2(new_n762), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n493), .ZN(new_n767));
  OR3_X1    g581(.A1(new_n767), .A2(KEYINPUT109), .A3(KEYINPUT46), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT109), .B1(new_n767), .B2(KEYINPUT46), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n492), .B1(new_n767), .B2(KEYINPUT46), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n459), .ZN(new_n772));
  XOR2_X1   g586(.A(new_n745), .B(KEYINPUT110), .Z(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n772), .A2(new_n695), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n556), .A2(new_n557), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n627), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT43), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n649), .A2(new_n653), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n780), .A2(KEYINPUT44), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(KEYINPUT44), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n775), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  NOR4_X1   g598(.A1(new_n706), .A2(new_n740), .A3(new_n700), .A4(new_n745), .ZN(new_n785));
  AND3_X1   g599(.A1(new_n771), .A2(KEYINPUT47), .A3(new_n459), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT47), .B1(new_n771), .B2(new_n459), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  NAND4_X1  g607(.A1(new_n740), .A2(new_n628), .A3(new_n392), .A4(new_n459), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n709), .A2(new_n491), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT49), .Z(new_n796));
  NOR4_X1   g610(.A1(new_n687), .A2(new_n794), .A3(new_n796), .A4(new_n776), .ZN(new_n797));
  AOI21_X1  g611(.A(G953), .B1(new_n797), .B2(new_n685), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n748), .A2(new_n749), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n459), .A3(new_n653), .A4(new_n662), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n686), .A2(new_n801), .A3(new_n730), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n673), .A2(new_n701), .B1(new_n684), .B2(new_n802), .ZN(new_n803));
  AND4_X1   g617(.A1(new_n799), .A2(new_n803), .A3(new_n674), .A4(new_n737), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n720), .A2(new_n654), .A3(new_n722), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n805), .A2(new_n700), .ZN(new_n806));
  AOI22_X1  g620(.A1(new_n673), .A2(new_n671), .B1(new_n806), .B2(new_n735), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n799), .B1(new_n807), .B2(new_n803), .ZN(new_n808));
  OAI21_X1  g622(.A(KEYINPUT113), .B1(new_n804), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n451), .A2(new_n457), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(KEYINPUT112), .A3(new_n744), .A4(new_n644), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT112), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n451), .A2(new_n457), .A3(new_n644), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n812), .B1(new_n813), .B2(new_n631), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n629), .A2(new_n630), .A3(new_n609), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n810), .A2(new_n644), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n811), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(new_n618), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n501), .A2(new_n610), .A3(new_n653), .ZN(new_n819));
  AOI22_X1  g633(.A1(new_n649), .A2(new_n819), .B1(new_n389), .B2(new_n611), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n706), .B(new_n712), .C1(new_n634), .C2(new_n645), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n610), .B1(new_n369), .B2(new_n388), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n723), .A2(new_n822), .B1(new_n729), .B2(new_n732), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n818), .A2(new_n820), .A3(new_n821), .A4(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n735), .A2(new_n736), .A3(new_n654), .A4(new_n751), .ZN(new_n825));
  INV_X1    g639(.A(new_n672), .ZN(new_n826));
  INV_X1    g640(.A(new_n745), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n548), .A2(new_n642), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n609), .A2(new_n641), .A3(new_n828), .A4(new_n662), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n706), .A2(new_n826), .A3(new_n827), .A4(new_n829), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n825), .A2(new_n830), .A3(new_n759), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(new_n756), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n824), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n684), .A2(new_n802), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n674), .A2(new_n702), .A3(new_n737), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT52), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT113), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n807), .A2(new_n799), .A3(new_n803), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n809), .A2(new_n833), .A3(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n804), .A2(new_n808), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n833), .A2(new_n843), .A3(KEYINPUT53), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n845), .A2(KEYINPUT54), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n833), .A2(new_n843), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n841), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n848), .B1(new_n841), .B2(new_n840), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT54), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n778), .A2(new_n563), .A3(new_n729), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(new_n391), .A3(new_n688), .A4(new_n710), .ZN(new_n854));
  XOR2_X1   g668(.A(new_n854), .B(KEYINPUT50), .Z(new_n855));
  NOR2_X1   g669(.A1(new_n745), .A2(new_n711), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n685), .A2(new_n740), .A3(new_n563), .A4(new_n856), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n857), .A2(new_n776), .A3(new_n628), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n778), .A2(new_n563), .A3(new_n856), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n615), .A2(new_n653), .A3(new_n728), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n855), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT114), .ZN(new_n864));
  INV_X1    g678(.A(new_n853), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n865), .A2(new_n774), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  AOI211_X1 g681(.A(new_n787), .B(new_n786), .C1(new_n460), .C2(new_n795), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n864), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n863), .A2(KEYINPUT114), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n852), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n863), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n868), .A2(KEYINPUT115), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n866), .B1(new_n868), .B2(KEYINPUT115), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n872), .B(KEYINPUT51), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n853), .A2(new_n720), .A3(new_n722), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n876), .B1(new_n631), .B2(new_n857), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT116), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n878), .B(KEYINPUT48), .C1(new_n860), .C2(new_n389), .ZN(new_n879));
  XOR2_X1   g693(.A(KEYINPUT116), .B(KEYINPUT48), .Z(new_n880));
  NOR3_X1   g694(.A1(new_n859), .A2(new_n743), .A3(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n877), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  AND4_X1   g696(.A1(new_n851), .A2(new_n871), .A3(new_n875), .A4(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(G952), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n798), .B1(new_n883), .B2(new_n884), .ZN(G75));
  NOR2_X1   g699(.A1(new_n232), .A2(G952), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n188), .B1(new_n842), .B2(new_n844), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT56), .B1(new_n887), .B2(G210), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n425), .B(new_n433), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT55), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n886), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n891), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n888), .A2(KEYINPUT117), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT117), .B1(new_n888), .B2(new_n893), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT118), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n892), .B(new_n898), .C1(new_n894), .C2(new_n895), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n897), .A2(new_n899), .ZN(G51));
  XNOR2_X1  g714(.A(new_n845), .B(KEYINPUT54), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n493), .B(KEYINPUT57), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n708), .B(KEYINPUT119), .Z(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n887), .A2(new_n766), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n886), .B1(new_n905), .B2(new_n906), .ZN(G54));
  INV_X1    g721(.A(new_n886), .ZN(new_n908));
  AND3_X1   g722(.A1(new_n887), .A2(KEYINPUT58), .A3(G475), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n908), .B1(new_n909), .B2(new_n537), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n910), .B1(new_n537), .B2(new_n909), .ZN(G60));
  NAND2_X1  g725(.A1(new_n846), .A2(new_n850), .ZN(new_n912));
  NAND2_X1  g726(.A1(G478), .A2(G902), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT59), .Z(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n624), .B1(new_n912), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n901), .A2(new_n624), .A3(new_n915), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n917), .A2(KEYINPUT120), .A3(new_n908), .A4(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT120), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n918), .A2(new_n908), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n920), .B1(new_n921), .B2(new_n916), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n919), .A2(new_n922), .ZN(G63));
  INV_X1    g737(.A(KEYINPUT122), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n650), .A2(new_n651), .ZN(new_n925));
  NAND2_X1  g739(.A1(G217), .A2(G902), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT60), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n837), .B1(new_n836), .B2(new_n838), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n821), .A2(new_n733), .A3(new_n725), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n612), .A2(new_n655), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n932), .A2(new_n756), .A3(new_n818), .A4(new_n831), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n929), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT53), .B1(new_n934), .B2(new_n839), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n833), .A2(new_n843), .A3(KEYINPUT53), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n925), .B(new_n928), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(KEYINPUT61), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n927), .B1(new_n842), .B2(new_n844), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n908), .B1(new_n939), .B2(new_n247), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n924), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(new_n939), .B2(new_n925), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n936), .B1(new_n841), .B2(new_n840), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n246), .B1(new_n944), .B2(new_n927), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n943), .A2(new_n945), .A3(KEYINPUT122), .A4(new_n908), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n941), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT121), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n937), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n939), .A2(KEYINPUT121), .A3(new_n925), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n949), .A2(new_n950), .A3(new_n945), .A4(new_n908), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n942), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n947), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT123), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT123), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n947), .A2(new_n952), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n954), .A2(new_n956), .ZN(G66));
  OAI21_X1  g771(.A(G953), .B1(new_n561), .B2(new_n430), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT124), .ZN(new_n959));
  INV_X1    g773(.A(new_n824), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n959), .B1(new_n960), .B2(new_n558), .ZN(new_n961));
  INV_X1    g775(.A(new_n425), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(G898), .B2(new_n232), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n961), .B(new_n963), .ZN(G69));
  NAND3_X1  g778(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(new_n533), .Z(new_n966));
  INV_X1    g780(.A(G227), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n558), .A2(G900), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n807), .A2(new_n702), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n698), .A2(new_n969), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n970), .A2(KEYINPUT62), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(KEYINPUT62), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n617), .A2(new_n745), .A3(new_n695), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n389), .B(new_n973), .C1(new_n744), .C2(new_n815), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n783), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n792), .A2(new_n971), .A3(new_n972), .A4(new_n975), .ZN(new_n976));
  OAI221_X1 g790(.A(new_n966), .B1(new_n967), .B2(new_n968), .C1(new_n976), .C2(new_n558), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n772), .A2(new_n695), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n686), .A2(new_n730), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n758), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n756), .B1(new_n980), .B2(new_n743), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n790), .B2(new_n791), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT125), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n783), .A2(new_n983), .A3(new_n969), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n983), .B1(new_n783), .B2(new_n969), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT126), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n982), .B(KEYINPUT126), .C1(new_n984), .C2(new_n985), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n558), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(new_n966), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n991), .B1(G227), .B2(new_n968), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n977), .B1(new_n990), .B2(new_n992), .ZN(G72));
  NAND2_X1  g807(.A1(G472), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT63), .Z(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n976), .B2(new_n824), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n361), .A2(new_n314), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n996), .A2(new_n342), .A3(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n376), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n997), .A2(new_n342), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n999), .A2(new_n995), .A3(new_n1000), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT127), .Z(new_n1002));
  AOI21_X1  g816(.A(new_n886), .B1(new_n849), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n998), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n988), .A2(new_n960), .A3(new_n989), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n995), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1004), .B1(new_n1006), .B2(new_n376), .ZN(G57));
endmodule


