//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:26 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1190, new_n1191, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  OAI21_X1  g0008(.A(G50), .B1(G58), .B2(G68), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G1), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n212), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT0), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G226), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n221), .B1(new_n201), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(KEYINPUT64), .B(G77), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(KEYINPUT65), .B(G244), .Z(new_n226));
  AOI21_X1  g0026(.A(new_n223), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n217), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n214), .B(new_n220), .C1(new_n233), .C2(KEYINPUT1), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G226), .B(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n201), .A2(G68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n203), .A2(G50), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n247), .B(new_n252), .Z(G351));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G1), .A3(G13), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G41), .ZN(new_n257));
  INV_X1    g0057(.A(G45), .ZN(new_n258));
  AOI21_X1  g0058(.A(G1), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G226), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n259), .A2(new_n255), .A3(G274), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT3), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(G1698), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G222), .ZN(new_n270));
  INV_X1    g0070(.A(G223), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT3), .B(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G1698), .ZN(new_n273));
  OAI221_X1 g0073(.A(new_n270), .B1(new_n271), .B2(new_n273), .C1(new_n224), .C2(new_n272), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n263), .B1(new_n274), .B2(new_n256), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT73), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(new_n276), .A3(G190), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n276), .B1(new_n275), .B2(G190), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n275), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G200), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n211), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n212), .A2(G33), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n287), .A2(new_n289), .B1(G20), .B2(new_n204), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n212), .A2(new_n264), .A3(KEYINPUT68), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT68), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(G20), .B2(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G150), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n285), .B1(new_n290), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G13), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n297), .A2(new_n212), .A3(G1), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(new_n284), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n215), .A2(G20), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(G50), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n298), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n301), .B1(G50), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n296), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT9), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n304), .A2(KEYINPUT9), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n282), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT10), .B1(new_n280), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n305), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(KEYINPUT10), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT72), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n282), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n281), .A2(KEYINPUT72), .A3(G200), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n308), .B1(new_n314), .B2(new_n280), .ZN(new_n315));
  INV_X1    g0115(.A(G179), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n275), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n304), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n317), .B(new_n318), .C1(G169), .C2(new_n275), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT74), .ZN(new_n321));
  INV_X1    g0121(.A(G274), .ZN(new_n322));
  INV_X1    g0122(.A(new_n211), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(new_n254), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n260), .A2(G238), .B1(new_n324), .B2(new_n259), .ZN(new_n325));
  INV_X1    g0125(.A(G1698), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n265), .A2(new_n267), .A3(G226), .A4(new_n326), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n265), .A2(new_n267), .A3(G232), .A4(G1698), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G33), .A2(G97), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n327), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n256), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n321), .B1(new_n332), .B2(KEYINPUT13), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT13), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(new_n325), .B2(new_n331), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n325), .A2(new_n331), .A3(KEYINPUT74), .A4(new_n334), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n333), .A2(new_n336), .A3(G190), .A4(new_n337), .ZN(new_n338));
  AND3_X1   g0138(.A1(new_n325), .A2(new_n331), .A3(new_n334), .ZN(new_n339));
  OAI21_X1  g0139(.A(G200), .B1(new_n339), .B2(new_n335), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n298), .A2(new_n203), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n341), .B(KEYINPUT12), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n299), .A2(G68), .A3(new_n300), .ZN(new_n343));
  INV_X1    g0143(.A(new_n294), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n344), .A2(new_n201), .ZN(new_n345));
  INV_X1    g0145(.A(G77), .ZN(new_n346));
  OAI22_X1  g0146(.A1(new_n288), .A2(new_n346), .B1(new_n212), .B2(G68), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n284), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT11), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n342), .B(new_n343), .C1(new_n348), .C2(new_n349), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n348), .A2(new_n349), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n338), .A2(new_n340), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  AND2_X1   g0154(.A1(KEYINPUT75), .A2(G169), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(new_n339), .B2(new_n335), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(KEYINPUT14), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n333), .A2(new_n336), .A3(G179), .A4(new_n337), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT14), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n359), .B(new_n355), .C1(new_n339), .C2(new_n335), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT76), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n357), .A2(new_n358), .A3(KEYINPUT76), .A4(new_n360), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n352), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT15), .B(G87), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT69), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(new_n368), .A3(new_n289), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n287), .A2(new_n294), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n225), .A2(G20), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT69), .B1(new_n366), .B2(new_n288), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n369), .A2(new_n370), .A3(new_n371), .A4(new_n372), .ZN(new_n373));
  AOI22_X1  g0173(.A1(new_n373), .A2(new_n284), .B1(new_n224), .B2(new_n298), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n299), .A2(G77), .A3(new_n300), .ZN(new_n375));
  XNOR2_X1  g0175(.A(new_n375), .B(KEYINPUT70), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(G200), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n269), .A2(G232), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n272), .A2(G238), .A3(G1698), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n268), .A2(G107), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n256), .ZN(new_n383));
  AOI22_X1  g0183(.A1(new_n260), .A2(new_n226), .B1(new_n324), .B2(new_n259), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n378), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n377), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT71), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n383), .A2(G190), .A3(new_n384), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT71), .B1(new_n377), .B2(new_n385), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n383), .A2(new_n384), .ZN(new_n392));
  INV_X1    g0192(.A(G169), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n383), .A2(new_n316), .A3(new_n384), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(new_n377), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  NOR4_X1   g0197(.A1(new_n320), .A2(new_n354), .A3(new_n365), .A4(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT18), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT80), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT7), .B1(new_n268), .B2(new_n212), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT7), .ZN(new_n402));
  AOI211_X1 g0202(.A(new_n402), .B(G20), .C1(new_n265), .C2(new_n267), .ZN(new_n403));
  OAI21_X1  g0203(.A(G68), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g0204(.A(G58), .B(G68), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n294), .A2(G159), .B1(new_n405), .B2(G20), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(KEYINPUT16), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT16), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n402), .B1(new_n272), .B2(G20), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n266), .A2(G33), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n411));
  OAI211_X1 g0211(.A(KEYINPUT7), .B(new_n212), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n203), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n405), .A2(G20), .ZN(new_n414));
  INV_X1    g0214(.A(G159), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n414), .B1(new_n344), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n408), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n407), .A2(new_n417), .A3(new_n284), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n286), .B1(new_n215), .B2(G20), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n419), .A2(new_n299), .B1(new_n298), .B2(new_n286), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n418), .A2(KEYINPUT77), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT77), .B1(new_n418), .B2(new_n420), .ZN(new_n422));
  NOR2_X1   g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n215), .B1(G41), .B2(G45), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n255), .A2(G232), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT78), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT78), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n255), .A2(new_n424), .A3(new_n427), .A4(G232), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(new_n262), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n271), .A2(new_n326), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n222), .A2(G1698), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n265), .A2(new_n430), .A3(new_n267), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(G33), .A2(G87), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n255), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n393), .B1(new_n429), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n434), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n428), .A2(new_n262), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n436), .A2(new_n437), .A3(new_n316), .A4(new_n426), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT79), .ZN(new_n439));
  AND3_X1   g0239(.A1(new_n435), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n439), .B1(new_n435), .B2(new_n438), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n400), .B1(new_n423), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n418), .A2(new_n420), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT77), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n418), .A2(KEYINPUT77), .A3(new_n420), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n446), .A2(new_n442), .A3(new_n400), .A4(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n399), .B1(new_n443), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT83), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT17), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT81), .ZN(new_n453));
  INV_X1    g0253(.A(G190), .ZN(new_n454));
  NOR2_X1   g0254(.A1(G223), .A2(G1698), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n455), .B1(new_n222), .B2(G1698), .ZN(new_n456));
  AOI22_X1  g0256(.A1(new_n456), .A2(new_n272), .B1(G33), .B2(G87), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n454), .B1(new_n457), .B2(new_n255), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n453), .B1(new_n458), .B2(new_n429), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n378), .B1(new_n429), .B2(new_n434), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n432), .A2(new_n433), .ZN(new_n461));
  AOI21_X1  g0261(.A(G190), .B1(new_n461), .B2(new_n256), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n462), .A2(KEYINPUT81), .A3(new_n426), .A4(new_n437), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n459), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(KEYINPUT82), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT82), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n459), .A2(new_n463), .A3(new_n466), .A4(new_n460), .ZN(new_n467));
  AOI211_X1 g0267(.A(new_n452), .B(new_n444), .C1(new_n465), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n465), .A2(new_n467), .ZN(new_n469));
  INV_X1    g0269(.A(new_n444), .ZN(new_n470));
  AOI21_X1  g0270(.A(KEYINPUT17), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n451), .B1(new_n468), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n469), .A2(new_n470), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n452), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n469), .A2(KEYINPUT17), .A3(new_n470), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n474), .A2(KEYINPUT83), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n446), .A2(new_n442), .A3(new_n447), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT80), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n478), .A2(KEYINPUT18), .A3(new_n448), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n450), .A2(new_n472), .A3(new_n476), .A4(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n398), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G97), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n298), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n215), .A2(G33), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n299), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(KEYINPUT84), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT84), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n299), .A2(new_n489), .A3(new_n486), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT6), .ZN(new_n492));
  INV_X1    g0292(.A(G107), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n484), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n492), .B1(new_n494), .B2(new_n206), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(KEYINPUT6), .A3(G97), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n497), .A2(G20), .B1(G77), .B2(new_n294), .ZN(new_n498));
  OAI21_X1  g0298(.A(G107), .B1(new_n401), .B2(new_n403), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  OAI221_X1 g0300(.A(new_n485), .B1(new_n484), .B2(new_n491), .C1(new_n500), .C2(new_n285), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT86), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT5), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n502), .B1(new_n503), .B2(G41), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n257), .A2(KEYINPUT86), .A3(KEYINPUT5), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n258), .A2(G1), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n507), .B(KEYINPUT85), .C1(KEYINPUT5), .C2(new_n257), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n215), .B(G45), .C1(new_n257), .C2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT85), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n506), .A2(new_n508), .A3(new_n511), .A4(new_n324), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n504), .A2(new_n505), .ZN(new_n513));
  OAI211_X1 g0313(.A(G257), .B(new_n255), .C1(new_n513), .C2(new_n509), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT87), .ZN(new_n516));
  XNOR2_X1  g0316(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n272), .A2(G250), .A3(G1698), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G283), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n272), .A2(G244), .A3(new_n326), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT4), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n518), .B(new_n519), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT4), .B1(new_n269), .B2(G244), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n256), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n517), .A2(new_n316), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n515), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n393), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n501), .A2(new_n525), .A3(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n515), .A2(new_n516), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT87), .B1(new_n512), .B2(new_n514), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n524), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT88), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n378), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n533), .B2(new_n532), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n527), .A2(new_n454), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n501), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n529), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n491), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G107), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n298), .A2(new_n493), .ZN(new_n541));
  XOR2_X1   g0341(.A(new_n541), .B(KEYINPUT25), .Z(new_n542));
  AND2_X1   g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(G33), .A2(G116), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n544), .A2(G20), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT23), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n212), .B2(G107), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n493), .A2(KEYINPUT23), .A3(G20), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n272), .A2(new_n212), .A3(G87), .ZN(new_n550));
  XOR2_X1   g0350(.A(KEYINPUT90), .B(KEYINPUT22), .Z(new_n551));
  AND2_X1   g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n550), .A2(new_n551), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n549), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT24), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT24), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n556), .B(new_n549), .C1(new_n552), .C2(new_n553), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n284), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n272), .A2(G257), .A3(G1698), .ZN(new_n560));
  NAND2_X1  g0360(.A1(G33), .A2(G294), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n265), .A2(new_n267), .A3(G250), .A4(new_n326), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n562), .A2(KEYINPUT91), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n562), .A2(KEYINPUT91), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n560), .B(new_n561), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n256), .ZN(new_n566));
  INV_X1    g0366(.A(new_n509), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n256), .B1(new_n506), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G264), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n566), .A2(new_n512), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(G200), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n565), .A2(new_n256), .B1(G264), .B2(new_n568), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n572), .A2(G190), .A3(new_n512), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n543), .A2(new_n559), .A3(new_n571), .A4(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n507), .A2(new_n322), .ZN(new_n575));
  INV_X1    g0375(.A(G250), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n258), .B2(G1), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n255), .A3(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n272), .A2(G238), .A3(new_n326), .ZN(new_n580));
  INV_X1    g0380(.A(G244), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n580), .B(new_n544), .C1(new_n273), .C2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n579), .B1(new_n582), .B2(new_n256), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n316), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n491), .A2(new_n366), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n366), .A2(new_n298), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n272), .A2(new_n212), .A3(G68), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT19), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n212), .B1(new_n329), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(G87), .B2(new_n207), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n588), .B1(new_n288), .B2(new_n484), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n587), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n586), .B1(new_n592), .B2(new_n285), .ZN(new_n593));
  OAI221_X1 g0393(.A(new_n584), .B1(G169), .B2(new_n583), .C1(new_n585), .C2(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n593), .B1(new_n539), .B2(G87), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n582), .A2(new_n256), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n578), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(G200), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n595), .B(new_n598), .C1(new_n454), .C2(new_n597), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n574), .A2(new_n594), .A3(new_n599), .ZN(new_n600));
  MUX2_X1   g0400(.A(new_n302), .B(new_n487), .S(G116), .Z(new_n601));
  OAI211_X1 g0401(.A(new_n519), .B(new_n212), .C1(G33), .C2(new_n484), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n602), .B(new_n284), .C1(new_n212), .C2(G116), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT20), .ZN(new_n604));
  XNOR2_X1  g0404(.A(new_n603), .B(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n393), .B1(new_n601), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n568), .A2(KEYINPUT89), .A3(G270), .ZN(new_n607));
  OAI211_X1 g0407(.A(G270), .B(new_n255), .C1(new_n513), .C2(new_n509), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT89), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n272), .A2(G257), .A3(new_n326), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n268), .A2(G303), .ZN(new_n613));
  INV_X1    g0413(.A(G264), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n612), .B(new_n613), .C1(new_n273), .C2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n256), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n611), .A2(new_n512), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n606), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT21), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT21), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n606), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n570), .A2(new_n393), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n572), .A2(new_n316), .A3(new_n512), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n540), .A2(new_n542), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n285), .B1(new_n555), .B2(new_n557), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n601), .A2(new_n605), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n628), .B1(new_n617), .B2(G200), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n454), .B2(new_n617), .ZN(new_n630));
  INV_X1    g0430(.A(new_n512), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n607), .B2(new_n610), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n316), .B1(new_n615), .B2(new_n256), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n628), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AND4_X1   g0434(.A1(new_n622), .A2(new_n627), .A3(new_n630), .A4(new_n634), .ZN(new_n635));
  AND4_X1   g0435(.A1(new_n483), .A2(new_n538), .A3(new_n600), .A4(new_n635), .ZN(G372));
  INV_X1    g0436(.A(new_n319), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n442), .A2(new_n444), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT18), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n442), .A2(new_n399), .A3(new_n444), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n396), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n365), .B1(new_n353), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n476), .A2(new_n472), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n641), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n637), .B1(new_n645), .B2(new_n315), .ZN(new_n646));
  INV_X1    g0446(.A(new_n594), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n599), .A2(new_n594), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n648), .A2(KEYINPUT26), .A3(new_n529), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n599), .A2(new_n594), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n501), .A2(new_n525), .A3(new_n528), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n650), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n647), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n622), .A2(new_n627), .A3(new_n634), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n538), .A2(new_n600), .A3(new_n655), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n646), .B1(new_n482), .B2(new_n657), .ZN(G369));
  NAND3_X1  g0458(.A1(new_n215), .A2(new_n212), .A3(G13), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(new_n661), .A3(G213), .ZN(new_n662));
  INV_X1    g0462(.A(G343), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n630), .B1(new_n628), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n622), .A2(new_n634), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n628), .A2(new_n664), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT92), .ZN(new_n669));
  XOR2_X1   g0469(.A(new_n667), .B(new_n669), .Z(new_n670));
  NOR2_X1   g0470(.A1(new_n627), .A2(new_n664), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n664), .B1(new_n625), .B2(new_n626), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n574), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n671), .B1(new_n627), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n670), .A2(G330), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n664), .B1(new_n622), .B2(new_n634), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n671), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g0478(.A(new_n678), .B(KEYINPUT93), .Z(G399));
  INV_X1    g0479(.A(new_n218), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G41), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G1), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n209), .B2(new_n682), .ZN(new_n685));
  XOR2_X1   g0485(.A(new_n685), .B(KEYINPUT28), .Z(new_n686));
  AOI21_X1  g0486(.A(new_n664), .B1(new_n654), .B2(new_n656), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT29), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI211_X1 g0489(.A(KEYINPUT29), .B(new_n664), .C1(new_n654), .C2(new_n656), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n664), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT94), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n572), .A2(new_n632), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n524), .A2(new_n633), .A3(new_n583), .A4(new_n526), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n597), .A2(new_n316), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n517), .B2(new_n524), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n572), .A2(new_n512), .B1(new_n632), .B2(new_n616), .ZN(new_n699));
  AOI22_X1  g0499(.A1(new_n696), .A2(KEYINPUT30), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT30), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n693), .B(new_n701), .C1(new_n694), .C2(new_n695), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n692), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n703), .A2(KEYINPUT31), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n635), .A2(new_n538), .A3(new_n600), .A4(new_n692), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n703), .A2(KEYINPUT31), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G330), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n691), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n686), .B1(new_n709), .B2(new_n215), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT95), .ZN(G364));
  NAND2_X1  g0511(.A1(new_n670), .A2(G330), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n297), .A2(G20), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n215), .B1(new_n713), .B2(G45), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n681), .A2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n712), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n670), .A2(G330), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G13), .A2(G33), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G20), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n670), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n211), .B1(G20), .B2(new_n393), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n680), .A2(new_n268), .ZN(new_n726));
  INV_X1    g0526(.A(G116), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n726), .A2(G355), .B1(new_n727), .B2(new_n680), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n680), .A2(new_n272), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(G45), .B2(new_n209), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n252), .A2(new_n258), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n728), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  AOI211_X1 g0532(.A(new_n722), .B(new_n725), .C1(new_n732), .C2(KEYINPUT96), .ZN(new_n733));
  OR2_X1    g0533(.A1(new_n732), .A2(KEYINPUT96), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n717), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n212), .A2(G190), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n378), .A2(G179), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G87), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n212), .A2(new_n454), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n737), .ZN(new_n741));
  OAI221_X1 g0541(.A(new_n272), .B1(new_n738), .B2(new_n493), .C1(new_n739), .C2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(G179), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n736), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  XNOR2_X1  g0545(.A(KEYINPUT98), .B(G159), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT32), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n212), .B1(new_n743), .B2(G190), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n484), .ZN(new_n751));
  NAND3_X1  g0551(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G190), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n203), .ZN(new_n755));
  OR4_X1    g0555(.A1(new_n742), .A2(new_n749), .A3(new_n751), .A4(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n316), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n740), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n736), .A2(new_n757), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n759), .A2(G58), .B1(new_n761), .B2(new_n225), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n752), .A2(new_n454), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n762), .B1(new_n201), .B2(new_n764), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT97), .Z(new_n766));
  INV_X1    g0566(.A(new_n741), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n272), .B1(new_n767), .B2(G303), .ZN(new_n768));
  INV_X1    g0568(.A(new_n750), .ZN(new_n769));
  XNOR2_X1  g0569(.A(KEYINPUT33), .B(G317), .ZN(new_n770));
  AOI22_X1  g0570(.A1(new_n769), .A2(G294), .B1(new_n753), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n763), .A2(G326), .ZN(new_n772));
  AND3_X1   g0572(.A1(new_n768), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n738), .ZN(new_n774));
  AOI22_X1  g0574(.A1(G322), .A2(new_n759), .B1(new_n774), .B2(G283), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n761), .A2(G311), .B1(new_n745), .B2(G329), .ZN(new_n776));
  AND3_X1   g0576(.A1(new_n773), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n756), .A2(new_n766), .B1(KEYINPUT99), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n778), .B1(KEYINPUT99), .B2(new_n777), .ZN(new_n779));
  INV_X1    g0579(.A(new_n725), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n735), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n718), .A2(new_n719), .B1(new_n724), .B2(new_n781), .ZN(G396));
  INV_X1    g0582(.A(KEYINPUT101), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n396), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g0584(.A1(new_n394), .A2(KEYINPUT101), .A3(new_n377), .A4(new_n395), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n377), .A2(new_n664), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n391), .A2(new_n784), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n642), .A2(new_n664), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n687), .A2(new_n790), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n791), .A2(KEYINPUT102), .ZN(new_n792));
  AND3_X1   g0592(.A1(new_n391), .A2(new_n784), .A3(new_n785), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n687), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n791), .A2(KEYINPUT102), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n792), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n716), .B1(new_n796), .B2(new_n708), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n708), .B2(new_n796), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n759), .A2(G143), .B1(new_n761), .B2(new_n747), .ZN(new_n799));
  INV_X1    g0599(.A(G150), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n799), .B1(new_n800), .B2(new_n754), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(G137), .B2(new_n763), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n802), .A2(KEYINPUT34), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(KEYINPUT34), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n272), .B1(new_n738), .B2(new_n203), .ZN(new_n805));
  INV_X1    g0605(.A(G132), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n741), .A2(new_n201), .B1(new_n744), .B2(new_n806), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n805), .B(new_n807), .C1(G58), .C2(new_n769), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n803), .A2(new_n804), .A3(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n761), .A2(G116), .B1(G283), .B2(new_n753), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT100), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n738), .A2(new_n739), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n741), .A2(new_n493), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n812), .B(new_n813), .C1(G294), .C2(new_n759), .ZN(new_n814));
  INV_X1    g0614(.A(G311), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n268), .B1(new_n744), .B2(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n751), .B(new_n816), .C1(G303), .C2(new_n763), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n811), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n780), .B1(new_n809), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n725), .A2(new_n720), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n717), .B(new_n819), .C1(new_n346), .C2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(new_n790), .B2(new_n721), .ZN(new_n822));
  AND2_X1   g0622(.A1(new_n798), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(G384));
  OR2_X1    g0624(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n497), .A2(KEYINPUT35), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n825), .A2(G116), .A3(new_n213), .A4(new_n826), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT36), .Z(new_n828));
  OAI211_X1 g0628(.A(new_n225), .B(new_n210), .C1(new_n202), .C2(new_n203), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n215), .B(G13), .C1(new_n829), .C2(new_n248), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT38), .ZN(new_n832));
  AND4_X1   g0632(.A1(new_n474), .A2(new_n640), .A3(new_n475), .A4(new_n639), .ZN(new_n833));
  INV_X1    g0633(.A(new_n662), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n446), .A2(new_n447), .A3(new_n834), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n473), .A2(new_n835), .A3(new_n638), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n423), .B1(new_n442), .B2(new_n834), .ZN(new_n837));
  AOI21_X1  g0637(.A(KEYINPUT37), .B1(new_n469), .B2(new_n470), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n836), .A2(KEYINPUT37), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n833), .A2(new_n835), .B1(new_n839), .B2(KEYINPUT104), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n839), .A2(KEYINPUT104), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n832), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n444), .A2(new_n834), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n480), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n473), .A2(new_n638), .A3(new_n843), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n846), .A2(KEYINPUT37), .B1(new_n837), .B2(new_n838), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n845), .A2(KEYINPUT38), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n842), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g0650(.A(KEYINPUT105), .B(KEYINPUT39), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT103), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n478), .A2(KEYINPUT18), .A3(new_n448), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT18), .B1(new_n478), .B2(new_n448), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AND2_X1   g0657(.A1(new_n476), .A2(new_n472), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n843), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n832), .B1(new_n859), .B2(new_n847), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n849), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n854), .B1(new_n861), .B2(KEYINPUT39), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT38), .B1(new_n845), .B2(new_n848), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n832), .B(new_n847), .C1(new_n480), .C2(new_n844), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n854), .B(KEYINPUT39), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n853), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n365), .A2(new_n692), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n641), .A2(new_n834), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n784), .A2(new_n785), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n687), .A2(new_n793), .B1(new_n692), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n363), .A2(new_n364), .ZN(new_n874));
  INV_X1    g0674(.A(new_n352), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n875), .A2(new_n664), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n876), .A2(new_n353), .A3(new_n877), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n875), .B(new_n664), .C1(new_n874), .C2(new_n354), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n873), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n871), .B1(new_n861), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n870), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n481), .B(new_n398), .C1(new_n689), .C2(new_n690), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n646), .ZN(new_n886));
  XNOR2_X1  g0686(.A(new_n884), .B(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n789), .B1(new_n878), .B2(new_n879), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT31), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n703), .B2(KEYINPUT106), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT106), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n891), .B(new_n692), .C1(new_n700), .C2(new_n702), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n705), .B(new_n706), .C1(new_n890), .C2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT40), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n888), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n864), .B2(new_n863), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n888), .A2(new_n893), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(new_n842), .B2(new_n849), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n896), .B1(new_n898), .B2(new_n894), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n899), .A2(new_n483), .A3(new_n893), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(G330), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n899), .B1(new_n483), .B2(new_n893), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n887), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n904), .B1(new_n215), .B2(new_n713), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n887), .A2(new_n903), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n831), .B1(new_n905), .B2(new_n906), .ZN(G367));
  OR2_X1    g0707(.A1(new_n595), .A2(new_n692), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n648), .A2(new_n908), .ZN(new_n909));
  OR2_X1    g0709(.A1(new_n908), .A2(new_n594), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n722), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n722), .A2(new_n725), .ZN(new_n914));
  INV_X1    g0714(.A(new_n729), .ZN(new_n915));
  OAI221_X1 g0715(.A(new_n914), .B1(new_n218), .B2(new_n366), .C1(new_n915), .C2(new_n243), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n716), .ZN(new_n917));
  OAI22_X1  g0717(.A1(new_n758), .A2(new_n800), .B1(new_n760), .B2(new_n201), .ZN(new_n918));
  INV_X1    g0718(.A(G143), .ZN(new_n919));
  OAI221_X1 g0719(.A(new_n272), .B1(new_n738), .B2(new_n224), .C1(new_n764), .C2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(KEYINPUT108), .B(G137), .ZN(new_n921));
  OAI22_X1  g0721(.A1(new_n741), .A2(new_n202), .B1(new_n744), .B2(new_n921), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n754), .A2(new_n746), .B1(new_n203), .B2(new_n750), .ZN(new_n923));
  OR4_X1    g0723(.A1(new_n918), .A2(new_n920), .A3(new_n922), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n767), .A2(G116), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT46), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n738), .A2(new_n484), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n927), .A2(new_n272), .ZN(new_n928));
  AOI22_X1  g0728(.A1(G303), .A2(new_n759), .B1(new_n745), .B2(G317), .ZN(new_n929));
  AOI22_X1  g0729(.A1(G294), .A2(new_n753), .B1(new_n763), .B2(G311), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n926), .A2(new_n928), .A3(new_n929), .A4(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(G283), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n760), .A2(new_n932), .B1(new_n750), .B2(new_n493), .ZN(new_n933));
  XOR2_X1   g0733(.A(new_n933), .B(KEYINPUT107), .Z(new_n934));
  OAI21_X1  g0734(.A(new_n924), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT47), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n917), .B1(new_n936), .B2(new_n725), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n913), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n501), .A2(new_n664), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n538), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n529), .A2(new_n664), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n677), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT45), .Z(new_n944));
  NOR2_X1   g0744(.A1(new_n677), .A2(new_n942), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(KEYINPUT44), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n944), .A2(new_n675), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n675), .B1(new_n944), .B2(new_n946), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n709), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n674), .B(new_n676), .Z(new_n951));
  XNOR2_X1  g0751(.A(new_n712), .B(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n949), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n950), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n681), .B(KEYINPUT41), .Z(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n715), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n535), .A2(new_n537), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(new_n627), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n664), .B1(new_n959), .B2(new_n652), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n942), .A2(new_n674), .A3(new_n676), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n960), .B1(new_n961), .B2(KEYINPUT42), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(KEYINPUT42), .B2(new_n961), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT43), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n963), .B1(new_n964), .B2(new_n912), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n912), .A2(new_n964), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n965), .B(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n942), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n675), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n967), .B(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n938), .B1(new_n957), .B2(new_n970), .ZN(G387));
  NAND2_X1  g0771(.A1(new_n952), .A2(new_n715), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n268), .B(new_n927), .C1(new_n287), .C2(new_n753), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n763), .A2(G159), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT110), .Z(new_n975));
  OAI22_X1  g0775(.A1(new_n201), .A2(new_n758), .B1(new_n741), .B2(new_n224), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n760), .A2(new_n203), .B1(new_n744), .B2(new_n800), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n769), .A2(new_n367), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n973), .A2(new_n975), .A3(new_n978), .A4(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n272), .B1(new_n745), .B2(G326), .ZN(new_n981));
  INV_X1    g0781(.A(G294), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n741), .A2(new_n982), .B1(new_n750), .B2(new_n932), .ZN(new_n983));
  AOI22_X1  g0783(.A1(G317), .A2(new_n759), .B1(new_n761), .B2(G303), .ZN(new_n984));
  XNOR2_X1  g0784(.A(KEYINPUT111), .B(G322), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n984), .B1(new_n764), .B2(new_n985), .C1(new_n815), .C2(new_n754), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT48), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n983), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n987), .B2(new_n986), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT49), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n981), .B1(new_n727), .B2(new_n738), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n989), .A2(new_n990), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n980), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n725), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n683), .B(new_n258), .C1(new_n203), .C2(new_n346), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT109), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(KEYINPUT50), .B1(new_n286), .B2(G50), .ZN(new_n998));
  OR3_X1    g0798(.A1(new_n286), .A2(KEYINPUT50), .A3(G50), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n995), .A2(new_n996), .ZN(new_n1001));
  OAI221_X1 g0801(.A(new_n729), .B1(new_n1000), .B2(new_n1001), .C1(new_n240), .C2(new_n258), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n726), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1002), .B1(G107), .B2(new_n218), .C1(new_n683), .C2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n717), .B1(new_n1004), .B2(new_n914), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n994), .B(new_n1005), .C1(new_n674), .C2(new_n723), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n952), .A2(new_n950), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n681), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n952), .A2(new_n950), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n972), .B(new_n1006), .C1(new_n1008), .C2(new_n1009), .ZN(G393));
  OAI21_X1  g0810(.A(new_n1007), .B1(new_n947), .B2(new_n948), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n953), .A2(new_n681), .A3(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n759), .A2(G311), .B1(G317), .B2(new_n763), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT52), .Z(new_n1014));
  OAI22_X1  g0814(.A1(new_n760), .A2(new_n982), .B1(new_n744), .B2(new_n985), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n1015), .B1(G283), .B2(new_n767), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n750), .A2(new_n727), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n268), .B1(new_n738), .B2(new_n493), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1017), .B(new_n1018), .C1(G303), .C2(new_n753), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1014), .A2(new_n1016), .A3(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n759), .A2(G159), .B1(G150), .B2(new_n763), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT51), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n741), .A2(new_n203), .B1(new_n744), .B2(new_n919), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT112), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n268), .B(new_n812), .C1(new_n287), .C2(new_n761), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n750), .A2(new_n346), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n753), .B2(G50), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1024), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1020), .B1(new_n1022), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n725), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n729), .A2(new_n247), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1031), .B(new_n914), .C1(new_n484), .C2(new_n218), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1030), .A2(new_n716), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n968), .B2(new_n722), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n949), .B2(new_n715), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1012), .A2(new_n1035), .ZN(G390));
  OAI21_X1  g0836(.A(new_n868), .B1(new_n873), .B2(new_n881), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n853), .B(new_n1037), .C1(new_n862), .C2(new_n866), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n707), .A2(G330), .A3(new_n790), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1039), .A2(new_n881), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n868), .B(KEYINPUT113), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n882), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n850), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1038), .A2(new_n1041), .A3(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(KEYINPUT39), .B1(new_n863), .B2(new_n864), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(KEYINPUT103), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n852), .B1(new_n1047), .B2(new_n865), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n1048), .A2(new_n1037), .B1(new_n850), .B2(new_n1043), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n888), .A2(new_n893), .A3(G330), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1045), .B(new_n715), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n820), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n716), .B1(new_n287), .B2(new_n1052), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT117), .Z(new_n1054));
  OAI22_X1  g0854(.A1(new_n758), .A2(new_n727), .B1(new_n760), .B2(new_n484), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n272), .B(new_n1055), .C1(G87), .C2(new_n767), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n764), .A2(new_n932), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1026), .B(new_n1057), .C1(G107), .C2(new_n753), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n738), .A2(new_n203), .B1(new_n744), .B2(new_n982), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT118), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1056), .A2(new_n1058), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n754), .A2(new_n921), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(KEYINPUT54), .B(G143), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n268), .B(new_n1064), .C1(new_n761), .C2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n769), .A2(G159), .B1(G128), .B2(new_n763), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n741), .A2(new_n800), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT53), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n758), .A2(new_n806), .B1(new_n738), .B2(new_n201), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(G125), .B2(new_n745), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1063), .A2(new_n1073), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1074), .A2(KEYINPUT119), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(KEYINPUT119), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n725), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1054), .B1(new_n1075), .B2(new_n1077), .C1(new_n867), .C2(new_n721), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1051), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1039), .A2(new_n881), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n873), .B1(new_n1080), .B2(new_n1050), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n873), .B1(new_n1039), .B2(new_n881), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n893), .A2(G330), .A3(new_n790), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n881), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1082), .B1(new_n1085), .B2(KEYINPUT115), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT115), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1081), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n398), .A2(new_n893), .A3(new_n481), .A4(G330), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n885), .A2(new_n646), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT114), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n885), .A2(new_n1090), .A3(KEYINPUT114), .A4(new_n646), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1089), .A2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1045), .B(new_n1096), .C1(new_n1049), .C2(new_n1050), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT116), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1097), .A2(new_n1098), .A3(new_n681), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1045), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1096), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1097), .A2(new_n681), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(KEYINPUT116), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1079), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(G378));
  NOR2_X1   g0907(.A1(new_n1048), .A2(new_n868), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n883), .ZN(new_n1109));
  XOR2_X1   g0909(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT123), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n320), .B(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n304), .A2(new_n662), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1113), .B(KEYINPUT55), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT121), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1112), .B(new_n1115), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n899), .A2(G330), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1116), .B1(new_n899), .B2(G330), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n1108), .A2(new_n1109), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n899), .A2(G330), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1116), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n899), .A2(G330), .A3(new_n1116), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n870), .A2(new_n1122), .A3(new_n883), .A4(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1119), .A2(new_n1124), .A3(new_n715), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n268), .A2(new_n257), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1126), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1126), .B1(G283), .B2(new_n745), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1128), .B1(new_n202), .B2(new_n738), .C1(new_n224), .C2(new_n741), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT120), .Z(new_n1130));
  OAI22_X1  g0930(.A1(new_n758), .A2(new_n493), .B1(new_n760), .B2(new_n366), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(G68), .B2(new_n769), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(G97), .A2(new_n753), .B1(new_n763), .B2(G116), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1130), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT58), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1127), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n754), .A2(new_n806), .B1(new_n750), .B2(new_n800), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(G128), .A2(new_n759), .B1(new_n767), .B2(new_n1066), .ZN(new_n1138));
  INV_X1    g0938(.A(G137), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1138), .B1(new_n1139), .B2(new_n760), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1137), .B(new_n1140), .C1(G125), .C2(new_n763), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1142), .A2(KEYINPUT59), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1142), .A2(KEYINPUT59), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n745), .A2(G124), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n264), .B(new_n257), .C1(new_n738), .C2(new_n746), .ZN(new_n1146));
  NOR4_X1   g0946(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .A4(new_n1146), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1136), .B(new_n1147), .C1(new_n1135), .C2(new_n1134), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n716), .B1(G50), .B2(new_n1052), .C1(new_n1148), .C2(new_n780), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n1116), .B2(new_n720), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT124), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1125), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1095), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1097), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1119), .A2(new_n1124), .A3(KEYINPUT57), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n681), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1097), .A2(new_n1153), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n1119), .A2(new_n1124), .ZN(new_n1158));
  AOI21_X1  g0958(.A(KEYINPUT57), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1152), .B1(new_n1156), .B2(new_n1159), .ZN(G375));
  NAND2_X1  g0960(.A1(new_n1089), .A2(new_n1095), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1101), .A2(new_n956), .A3(new_n1161), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n880), .A2(new_n721), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT125), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n717), .B1(new_n203), .B2(new_n820), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n758), .A2(new_n932), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n346), .A2(new_n738), .B1(new_n760), .B2(new_n493), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n1166), .B(new_n1167), .C1(G97), .C2(new_n767), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G116), .A2(new_n753), .B1(new_n763), .B2(G294), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n272), .B1(new_n745), .B2(G303), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1169), .A2(new_n979), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n741), .A2(new_n415), .ZN(new_n1173));
  OAI22_X1  g0973(.A1(new_n758), .A2(new_n921), .B1(new_n760), .B2(new_n800), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(G128), .C2(new_n745), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n268), .B1(new_n774), .B2(G58), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n1066), .A2(new_n753), .B1(G132), .B2(new_n763), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1176), .B(new_n1177), .C1(new_n201), .C2(new_n750), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1168), .A2(new_n1172), .B1(new_n1175), .B2(new_n1179), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1164), .B(new_n1165), .C1(new_n780), .C2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n1089), .B2(new_n714), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1162), .A2(new_n1183), .ZN(G381));
  INV_X1    g0984(.A(G387), .ZN(new_n1185));
  INV_X1    g0985(.A(G390), .ZN(new_n1186));
  NOR3_X1   g0986(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  OR4_X1    g0988(.A1(G378), .A2(G375), .A3(new_n1188), .A4(G381), .ZN(G407));
  NAND2_X1  g0989(.A1(new_n663), .A2(G213), .ZN(new_n1190));
  OR3_X1    g0990(.A1(G378), .A2(G375), .A3(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(G407), .A2(new_n1191), .A3(G213), .ZN(G409));
  NAND3_X1  g0992(.A1(new_n1157), .A2(new_n1158), .A3(new_n956), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n1152), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1105), .A2(new_n1102), .A3(new_n1099), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1079), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(G375), .B2(new_n1106), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1089), .A2(new_n1095), .A3(KEYINPUT60), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1199), .A2(new_n681), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT60), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1161), .B1(new_n1096), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1203), .A2(G384), .A3(new_n1183), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(G384), .B1(new_n1203), .B2(new_n1183), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1198), .A2(new_n1190), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(KEYINPUT62), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1198), .A2(new_n1190), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n663), .A2(G213), .A3(G2897), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1207), .B(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT61), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT62), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1198), .A2(new_n1216), .A3(new_n1190), .A4(new_n1207), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1209), .A2(new_n1214), .A3(new_n1215), .A4(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1185), .A2(G390), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(G387), .A2(new_n1186), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(KEYINPUT126), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(G393), .B(G396), .ZN(new_n1222));
  AND4_X1   g1022(.A1(new_n1219), .A2(new_n1221), .A3(new_n1220), .A4(new_n1222), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1221), .A2(new_n1222), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1218), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT61), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1225), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT63), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1208), .A2(new_n1229), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1198), .A2(KEYINPUT63), .A3(new_n1190), .A4(new_n1207), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1227), .A2(new_n1228), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1226), .A2(new_n1232), .ZN(G405));
  AND2_X1   g1033(.A1(G375), .A2(new_n1106), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(G375), .A2(new_n1106), .ZN(new_n1235));
  OR3_X1    g1035(.A1(new_n1234), .A2(new_n1235), .A3(new_n1207), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1207), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1236), .A2(new_n1225), .A3(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1225), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(G402));
endmodule


