//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n838, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n949, new_n950;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  AOI21_X1  g004(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n206));
  OR2_X1    g005(.A1(new_n206), .A2(KEYINPUT72), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(KEYINPUT72), .ZN(new_n208));
  XNOR2_X1  g007(.A(G197gat), .B(G204gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(G211gat), .B(G218gat), .Z(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214));
  INV_X1    g013(.A(G183gat), .ZN(new_n215));
  INV_X1    g014(.A(G190gat), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT67), .B(G183gat), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT68), .ZN(new_n221));
  OR3_X1    g020(.A1(new_n220), .A2(new_n221), .A3(G190gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n221), .B1(new_n220), .B2(G190gat), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n219), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n225));
  NOR2_X1   g024(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT66), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n230));
  OAI221_X1 g029(.A(new_n230), .B1(G169gat), .B2(G176gat), .C1(new_n225), .C2(new_n226), .ZN(new_n231));
  INV_X1    g030(.A(G169gat), .ZN(new_n232));
  INV_X1    g031(.A(G176gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n234), .B1(KEYINPUT23), .B2(new_n228), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n229), .A2(KEYINPUT25), .A3(new_n231), .A4(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT64), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n237), .ZN(new_n238));
  NAND4_X1  g037(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n215), .A2(new_n216), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n217), .A2(new_n238), .A3(new_n239), .A4(new_n240), .ZN(new_n241));
  AND4_X1   g040(.A1(new_n229), .A2(new_n241), .A3(new_n231), .A4(new_n235), .ZN(new_n242));
  OAI22_X1  g041(.A1(new_n224), .A2(new_n236), .B1(new_n242), .B2(KEYINPUT25), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT27), .B(G183gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(KEYINPUT28), .A3(new_n216), .ZN(new_n245));
  NOR2_X1   g044(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n246), .B1(new_n220), .B2(KEYINPUT27), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n247), .A2(G190gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n245), .B1(new_n248), .B2(KEYINPUT28), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n215), .A2(new_n216), .ZN(new_n250));
  NOR3_X1   g049(.A1(new_n234), .A2(KEYINPUT26), .A3(new_n228), .ZN(new_n251));
  AOI211_X1 g050(.A(new_n250), .B(new_n251), .C1(KEYINPUT26), .C2(new_n228), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n243), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(G226gat), .A3(G233gat), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT29), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n254), .A2(new_n257), .B1(G226gat), .B2(G233gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n213), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G226gat), .A2(G233gat), .ZN(new_n260));
  INV_X1    g059(.A(new_n254), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n260), .B1(new_n261), .B2(KEYINPUT29), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n262), .A2(new_n212), .A3(new_n255), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT37), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n205), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n264), .A2(KEYINPUT37), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT38), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G1gat), .B(G29gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT0), .ZN(new_n271));
  XOR2_X1   g070(.A(G57gat), .B(G85gat), .Z(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT84), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G127gat), .B(G134gat), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n276), .A2(KEYINPUT69), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(KEYINPUT69), .ZN(new_n278));
  INV_X1    g077(.A(G113gat), .ZN(new_n279));
  INV_X1    g078(.A(G120gat), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT1), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G113gat), .A2(G120gat), .ZN(new_n282));
  AND2_X1   g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n277), .A2(new_n278), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n281), .A2(new_n282), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n285), .A2(KEYINPUT69), .A3(new_n276), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G148gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G141gat), .ZN(new_n289));
  INV_X1    g088(.A(G141gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G148gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT76), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n289), .A2(new_n291), .B1(new_n292), .B2(KEYINPUT2), .ZN(new_n293));
  NAND2_X1  g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT76), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n292), .A2(G155gat), .A3(G162gat), .ZN(new_n296));
  INV_X1    g095(.A(G155gat), .ZN(new_n297));
  INV_X1    g096(.A(G162gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n295), .A2(new_n296), .A3(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n293), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n294), .B1(new_n299), .B2(KEYINPUT2), .ZN(new_n302));
  OR3_X1    g101(.A1(new_n290), .A2(KEYINPUT77), .A3(G148gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n289), .A2(KEYINPUT77), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n303), .A2(new_n304), .A3(new_n291), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n301), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n287), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT4), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n287), .A2(new_n306), .A3(KEYINPUT4), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G225gat), .A2(G233gat), .ZN(new_n312));
  XOR2_X1   g111(.A(KEYINPUT78), .B(KEYINPUT3), .Z(new_n313));
  NAND2_X1  g112(.A1(new_n306), .A2(new_n313), .ZN(new_n314));
  OR2_X1    g113(.A1(new_n293), .A2(new_n300), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n305), .A2(new_n302), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT3), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n284), .A2(new_n286), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n314), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n321));
  NAND4_X1  g120(.A1(new_n311), .A2(new_n312), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n317), .A2(new_n286), .A3(new_n284), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n312), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n321), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n320), .A2(new_n309), .A3(new_n310), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n326), .B1(new_n327), .B2(new_n325), .ZN(new_n328));
  AND3_X1   g127(.A1(new_n322), .A2(new_n328), .A3(KEYINPUT85), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT85), .B1(new_n322), .B2(new_n328), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n275), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n322), .A2(new_n328), .A3(new_n273), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT6), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n273), .B1(new_n322), .B2(new_n328), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n331), .A2(new_n334), .B1(KEYINPUT6), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n259), .A2(new_n263), .A3(new_n204), .ZN(new_n337));
  AND2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n204), .B(KEYINPUT73), .Z(new_n339));
  NOR3_X1   g138(.A1(new_n268), .A2(KEYINPUT38), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n263), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n341), .A2(KEYINPUT86), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n259), .B1(new_n341), .B2(KEYINPUT86), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT37), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT87), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n340), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n345), .B1(new_n340), .B2(new_n344), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n269), .B(new_n338), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  XOR2_X1   g147(.A(G78gat), .B(G106gat), .Z(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT31), .B(G50gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT83), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n314), .A2(new_n257), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n213), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n306), .A2(KEYINPUT29), .ZN(new_n356));
  AOI22_X1  g155(.A1(new_n356), .A2(new_n212), .B1(KEYINPUT3), .B2(new_n317), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n355), .B1(new_n357), .B2(KEYINPUT82), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n356), .A2(new_n212), .ZN(new_n359));
  AND3_X1   g158(.A1(new_n359), .A2(KEYINPUT82), .A3(new_n318), .ZN(new_n360));
  OAI211_X1 g159(.A(G228gat), .B(G233gat), .C1(new_n358), .C2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(G22gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n313), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n317), .A2(new_n363), .B1(G228gat), .B2(G233gat), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n355), .A2(new_n359), .A3(new_n364), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n361), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n362), .B1(new_n361), .B2(new_n365), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n353), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n361), .A2(new_n365), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(G22gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n361), .A2(new_n362), .A3(new_n365), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n351), .B(new_n352), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n327), .A2(new_n325), .ZN(new_n376));
  OAI211_X1 g175(.A(new_n376), .B(KEYINPUT39), .C1(new_n325), .C2(new_n324), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n377), .B(new_n274), .C1(KEYINPUT39), .C2(new_n376), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n378), .B(KEYINPUT40), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n379), .A2(new_n331), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n259), .A2(new_n263), .A3(new_n204), .ZN(new_n381));
  INV_X1    g180(.A(new_n339), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n381), .A2(KEYINPUT30), .B1(new_n264), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT74), .B(KEYINPUT30), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n337), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT75), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT75), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n337), .A2(new_n387), .A3(new_n384), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n383), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n375), .B1(new_n380), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n348), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n335), .A2(KEYINPUT6), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n333), .B(new_n332), .C1(new_n335), .C2(KEYINPUT80), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n335), .A2(KEYINPUT80), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n395), .A2(new_n383), .A3(new_n388), .A4(new_n386), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT81), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT30), .ZN(new_n399));
  OAI22_X1  g198(.A1(new_n265), .A2(new_n339), .B1(new_n337), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n387), .B1(new_n337), .B2(new_n384), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n402), .A2(KEYINPUT81), .A3(new_n388), .A4(new_n395), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n375), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n254), .A2(new_n287), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n243), .A2(new_n253), .A3(new_n319), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT34), .ZN(new_n409));
  NAND2_X1  g208(.A1(G227gat), .A2(G233gat), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n409), .B1(new_n408), .B2(new_n410), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n406), .A2(G227gat), .A3(G233gat), .A4(new_n407), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT70), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT32), .ZN(new_n417));
  XNOR2_X1  g216(.A(G15gat), .B(G43gat), .ZN(new_n418));
  XNOR2_X1  g217(.A(G71gat), .B(G99gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n417), .B1(new_n421), .B2(KEYINPUT33), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n415), .A2(new_n416), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n416), .B1(new_n415), .B2(new_n422), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n417), .A2(KEYINPUT33), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n420), .B1(new_n415), .B2(new_n427), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n414), .B(KEYINPUT71), .C1(new_n426), .C2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n425), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n423), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT71), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n432), .B1(new_n412), .B2(new_n413), .ZN(new_n433));
  INV_X1    g232(.A(new_n413), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n434), .A2(KEYINPUT71), .A3(new_n411), .ZN(new_n435));
  INV_X1    g234(.A(new_n428), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n431), .A2(new_n433), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n429), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT36), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n391), .A2(new_n405), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  AOI221_X4 g240(.A(KEYINPUT89), .B1(new_n368), .B2(new_n373), .C1(new_n429), .C2(new_n437), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT89), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n443), .B1(new_n438), .B2(new_n374), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT35), .B1(new_n445), .B2(new_n404), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT90), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n389), .A2(new_n336), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT88), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n438), .A2(new_n374), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n451), .A2(KEYINPUT35), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n446), .A2(new_n447), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  OAI211_X1 g252(.A(KEYINPUT90), .B(KEYINPUT35), .C1(new_n445), .C2(new_n404), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n441), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(G50gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(G43gat), .ZN(new_n457));
  INV_X1    g256(.A(G43gat), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(G50gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT91), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT91), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n457), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n461), .A2(KEYINPUT15), .A3(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT92), .B1(new_n456), .B2(G43gat), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT92), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n466), .A2(new_n458), .A3(G50gat), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n467), .A3(new_n457), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT15), .ZN(new_n469));
  INV_X1    g268(.A(G36gat), .ZN(new_n470));
  AND2_X1   g269(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n471));
  NOR2_X1   g270(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(G29gat), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n474), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n468), .A2(new_n469), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n464), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n473), .A2(new_n475), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n478), .A2(new_n461), .A3(KEYINPUT15), .A4(new_n463), .ZN(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT17), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(G15gat), .B(G22gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n482), .A2(G1gat), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT93), .ZN(new_n484));
  OAI21_X1  g283(.A(G8gat), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(G1gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT16), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(G1gat), .B2(new_n482), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n485), .B(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT17), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n479), .B(new_n491), .C1(new_n464), .C2(new_n476), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n481), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(G229gat), .A2(G233gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n477), .A2(new_n480), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n489), .B(G8gat), .C1(new_n484), .C2(new_n483), .ZN(new_n496));
  INV_X1    g295(.A(new_n483), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n485), .A2(new_n497), .A3(new_n488), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n493), .A2(new_n494), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT18), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n495), .B(new_n499), .ZN(new_n504));
  XOR2_X1   g303(.A(KEYINPUT94), .B(KEYINPUT13), .Z(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(new_n494), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n493), .A2(KEYINPUT18), .A3(new_n494), .A4(new_n500), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n503), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G113gat), .B(G141gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(G197gat), .ZN(new_n511));
  XOR2_X1   g310(.A(KEYINPUT11), .B(G169gat), .Z(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(KEYINPUT12), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n509), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n503), .A2(new_n507), .A3(new_n514), .A4(new_n508), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(G190gat), .B(G218gat), .Z(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(G99gat), .A2(G106gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT8), .ZN(new_n523));
  NAND2_X1  g322(.A1(G85gat), .A2(G92gat), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(G85gat), .ZN(new_n527));
  INV_X1    g326(.A(G92gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n523), .A2(new_n526), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G99gat), .B(G106gat), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AND3_X1   g333(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI22_X1  g336(.A1(KEYINPUT8), .A2(new_n522), .B1(new_n527), .B2(new_n528), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n532), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g339(.A1(G232gat), .A2(G233gat), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n495), .A2(new_n540), .B1(KEYINPUT41), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n540), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n481), .A2(new_n492), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n521), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n541), .A2(KEYINPUT41), .ZN(new_n547));
  XNOR2_X1  g346(.A(G134gat), .B(G162gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(KEYINPUT97), .B(KEYINPUT98), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n542), .A2(new_n544), .A3(new_n521), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n546), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n551), .ZN(new_n554));
  INV_X1    g353(.A(new_n552), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n554), .B1(new_n555), .B2(new_n545), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G71gat), .B(G78gat), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n560));
  AND2_X1   g359(.A1(G57gat), .A2(G64gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(G57gat), .A2(G64gat), .ZN(new_n562));
  NOR3_X1   g361(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n559), .B1(new_n563), .B2(KEYINPUT95), .ZN(new_n564));
  NAND2_X1  g363(.A1(G71gat), .A2(G78gat), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OR2_X1    g366(.A1(G57gat), .A2(G64gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(G57gat), .A2(G64gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT95), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(new_n571), .A3(new_n558), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n564), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n499), .B1(KEYINPUT21), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT21), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n564), .A2(new_n576), .A3(new_n572), .ZN(new_n577));
  XNOR2_X1  g376(.A(G127gat), .B(G155gat), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n577), .B(new_n578), .Z(new_n579));
  NAND2_X1  g378(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n579), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n574), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT96), .ZN(new_n585));
  XOR2_X1   g384(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G183gat), .B(G211gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n583), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n580), .A2(new_n582), .A3(new_n589), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT99), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n537), .A2(new_n532), .A3(new_n538), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n531), .A2(new_n533), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n570), .A2(new_n571), .A3(new_n558), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n558), .B1(new_n570), .B2(new_n571), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n595), .B(new_n596), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT10), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n594), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI211_X1 g400(.A(new_n564), .B(new_n572), .C1(new_n534), .C2(new_n539), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n599), .A2(new_n602), .A3(new_n600), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n540), .A2(new_n573), .A3(KEYINPUT99), .A4(KEYINPUT10), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n601), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G230gat), .A2(G233gat), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n606), .B(KEYINPUT100), .Z(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n599), .A2(new_n602), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n607), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G120gat), .B(G148gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(G176gat), .B(G204gat), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n613), .B(new_n614), .Z(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n609), .A2(new_n611), .A3(new_n615), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  AND3_X1   g419(.A1(new_n557), .A2(new_n593), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NOR3_X1   g421(.A1(new_n455), .A2(new_n519), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT101), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n395), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n395), .A2(new_n624), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n623), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g428(.A1(new_n450), .A2(new_n452), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT35), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n451), .A2(KEYINPUT89), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n438), .A2(new_n443), .A3(new_n374), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(new_n398), .A2(new_n403), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n631), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n630), .B1(new_n636), .B2(KEYINPUT90), .ZN(new_n637));
  INV_X1    g436(.A(new_n454), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n440), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n639), .A2(new_n518), .A3(new_n389), .A4(new_n621), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT102), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n446), .A2(new_n447), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n643), .A2(new_n454), .A3(new_n630), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n519), .B1(new_n644), .B2(new_n440), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n645), .A2(KEYINPUT102), .A3(new_n389), .A4(new_n621), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  XOR2_X1   g446(.A(KEYINPUT16), .B(G8gat), .Z(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT42), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n642), .A2(G8gat), .A3(new_n646), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n623), .A2(KEYINPUT42), .A3(new_n389), .A4(new_n648), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n651), .A2(new_n654), .A3(KEYINPUT103), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT103), .ZN(new_n656));
  AOI21_X1  g455(.A(KEYINPUT42), .B1(new_n647), .B2(new_n648), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n652), .A2(new_n653), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n655), .A2(new_n659), .ZN(G1325gat));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n621), .ZN(new_n661));
  OAI21_X1  g460(.A(G15gat), .B1(new_n661), .B2(new_n439), .ZN(new_n662));
  INV_X1    g461(.A(G15gat), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n623), .A2(new_n663), .A3(new_n438), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(KEYINPUT104), .Z(G1326gat));
  OAI21_X1  g465(.A(KEYINPUT105), .B1(new_n661), .B2(new_n374), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n623), .A2(new_n668), .A3(new_n375), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT43), .B(G22gat), .ZN(new_n671));
  XOR2_X1   g470(.A(new_n670), .B(new_n671), .Z(G1327gat));
  NOR2_X1   g471(.A1(new_n593), .A2(new_n619), .ZN(new_n673));
  INV_X1    g472(.A(new_n557), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT106), .ZN(new_n676));
  NOR3_X1   g475(.A1(new_n455), .A2(new_n519), .A3(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n677), .A2(new_n474), .A3(new_n627), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT45), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n680), .B1(new_n455), .B2(new_n557), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n639), .A2(KEYINPUT44), .A3(new_n674), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n516), .A2(KEYINPUT107), .A3(new_n517), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT107), .B1(new_n516), .B2(new_n517), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g485(.A1(new_n686), .A2(new_n673), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n683), .A2(new_n627), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n679), .B1(new_n474), .B2(new_n688), .ZN(G1328gat));
  NAND3_X1  g488(.A1(new_n677), .A2(new_n470), .A3(new_n389), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT46), .Z(new_n691));
  AND3_X1   g490(.A1(new_n683), .A2(new_n389), .A3(new_n687), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n691), .B1(new_n470), .B2(new_n692), .ZN(G1329gat));
  INV_X1    g492(.A(new_n439), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n681), .A2(new_n682), .A3(new_n694), .A4(new_n687), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(G43gat), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT108), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT47), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n677), .A2(new_n458), .A3(new_n438), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n696), .B(new_n699), .C1(new_n697), .C2(KEYINPUT47), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(G1330gat));
  NAND3_X1  g502(.A1(new_n677), .A2(new_n456), .A3(new_n375), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n681), .A2(new_n682), .A3(new_n375), .A4(new_n687), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT110), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(G50gat), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n705), .A2(new_n706), .ZN(new_n709));
  OAI211_X1 g508(.A(KEYINPUT48), .B(new_n704), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n705), .A2(G50gat), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n711), .A2(KEYINPUT109), .A3(new_n704), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT48), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n705), .A2(new_n714), .A3(G50gat), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n710), .A2(new_n716), .ZN(G1331gat));
  NAND3_X1  g516(.A1(new_n557), .A2(new_n593), .A3(new_n619), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n455), .A2(new_n686), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n627), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g520(.A1(new_n389), .A2(KEYINPUT111), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n389), .A2(KEYINPUT111), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT49), .ZN(new_n725));
  INV_X1    g524(.A(G64gat), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  XOR2_X1   g526(.A(new_n727), .B(KEYINPUT112), .Z(new_n728));
  NAND2_X1  g527(.A1(new_n719), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n725), .A2(new_n726), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1333gat));
  INV_X1    g530(.A(G71gat), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n719), .A2(new_n732), .A3(new_n438), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n719), .A2(new_n694), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n733), .B1(new_n734), .B2(new_n732), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT50), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1334gat));
  NAND2_X1  g536(.A1(new_n719), .A2(new_n375), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(G78gat), .ZN(G1335gat));
  INV_X1    g538(.A(new_n686), .ZN(new_n740));
  INV_X1    g539(.A(new_n593), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT113), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n620), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n681), .A2(new_n682), .A3(new_n627), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(KEYINPUT114), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G85gat), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n745), .A2(KEYINPUT114), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n455), .A2(new_n557), .ZN(new_n749));
  INV_X1    g548(.A(new_n743), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n749), .A2(KEYINPUT115), .A3(KEYINPUT51), .A4(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n639), .A2(new_n674), .A3(new_n750), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n639), .A2(KEYINPUT51), .A3(new_n674), .A4(new_n750), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT115), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n751), .A2(new_n754), .A3(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n627), .A2(new_n527), .A3(new_n619), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n747), .A2(new_n748), .B1(new_n759), .B2(new_n760), .ZN(G1336gat));
  NAND4_X1  g560(.A1(new_n681), .A2(new_n682), .A3(new_n724), .A4(new_n744), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT116), .ZN(new_n763));
  OR2_X1    g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n528), .B1(new_n762), .B2(new_n763), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n724), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n767), .A2(G92gat), .A3(new_n620), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT52), .B1(new_n758), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT51), .B1(new_n749), .B2(new_n750), .ZN(new_n771));
  INV_X1    g570(.A(new_n755), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n768), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n681), .A2(new_n682), .A3(new_n389), .A4(new_n744), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G92gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT52), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n770), .A2(new_n777), .ZN(G1337gat));
  AND3_X1   g577(.A1(new_n683), .A2(new_n694), .A3(new_n744), .ZN(new_n779));
  INV_X1    g578(.A(G99gat), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n438), .A2(new_n780), .A3(new_n619), .ZN(new_n781));
  OAI22_X1  g580(.A1(new_n779), .A2(new_n780), .B1(new_n759), .B2(new_n781), .ZN(G1338gat));
  NOR3_X1   g581(.A1(new_n374), .A2(G106gat), .A3(new_n620), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n758), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n681), .A2(new_n682), .A3(new_n375), .A4(new_n744), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G106gat), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n784), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n783), .B(KEYINPUT117), .Z(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(new_n771), .B2(new_n772), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n790), .A2(new_n787), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n788), .B1(new_n785), .B2(new_n791), .ZN(G1339gat));
  OAI21_X1  g591(.A(KEYINPUT118), .B1(new_n622), .B2(new_n686), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n621), .B(new_n794), .C1(new_n685), .C2(new_n684), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n605), .A2(new_n797), .A3(new_n608), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n798), .A2(KEYINPUT55), .A3(new_n616), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n601), .A2(new_n603), .A3(new_n607), .A4(new_n604), .ZN(new_n800));
  AND4_X1   g599(.A1(KEYINPUT119), .A2(new_n609), .A3(KEYINPUT54), .A4(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n797), .B1(new_n605), .B2(new_n608), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT119), .B1(new_n802), .B2(new_n800), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n799), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n798), .A2(new_n616), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n609), .A2(KEYINPUT54), .A3(new_n800), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT119), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n802), .A2(KEYINPUT119), .A3(new_n800), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n805), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n618), .B(new_n804), .C1(new_n810), .C2(KEYINPUT55), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n504), .A2(new_n506), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n494), .B1(new_n493), .B2(new_n500), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n513), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n517), .ZN(new_n815));
  OR3_X1    g614(.A1(new_n811), .A2(new_n557), .A3(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n619), .A2(new_n517), .A3(new_n814), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT120), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n619), .A2(new_n814), .A3(new_n517), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n811), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n821), .B1(new_n686), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n816), .B1(new_n823), .B2(new_n674), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n796), .B1(new_n824), .B2(new_n741), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(new_n375), .ZN(new_n826));
  NAND4_X1  g625(.A1(new_n826), .A2(new_n438), .A3(new_n627), .A4(new_n767), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n827), .A2(new_n279), .A3(new_n519), .ZN(new_n828));
  INV_X1    g627(.A(new_n627), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n634), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(new_n724), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n686), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n828), .B1(new_n279), .B2(new_n833), .ZN(G1340gat));
  NOR3_X1   g633(.A1(new_n827), .A2(new_n280), .A3(new_n620), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n619), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n835), .B1(new_n280), .B2(new_n836), .ZN(G1341gat));
  INV_X1    g636(.A(G127gat), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n832), .A2(new_n838), .A3(new_n593), .ZN(new_n839));
  OAI21_X1  g638(.A(G127gat), .B1(new_n827), .B2(new_n741), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(G1342gat));
  NAND3_X1  g640(.A1(new_n402), .A2(new_n388), .A3(new_n674), .ZN(new_n842));
  OR3_X1    g641(.A1(new_n831), .A2(G134gat), .A3(new_n842), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n844));
  OAI21_X1  g643(.A(G134gat), .B1(new_n827), .B2(new_n557), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(KEYINPUT56), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(G1343gat));
  NOR4_X1   g646(.A1(new_n825), .A2(new_n694), .A3(new_n829), .A4(new_n374), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(new_n767), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n849), .A2(G141gat), .A3(new_n519), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(KEYINPUT58), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n694), .A2(new_n829), .A3(new_n724), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT122), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n374), .A2(new_n854), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n811), .A2(new_n557), .A3(new_n815), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n817), .B1(new_n811), .B2(new_n519), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n557), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n805), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n861), .B1(new_n801), .B2(new_n803), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT55), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n864), .A2(new_n518), .A3(new_n618), .A4(new_n804), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n674), .B1(new_n865), .B2(new_n817), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT121), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n593), .B1(new_n860), .B2(new_n867), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n853), .B(new_n855), .C1(new_n868), .C2(new_n796), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n854), .B1(new_n825), .B2(new_n374), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n867), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n816), .B1(new_n866), .B2(KEYINPUT121), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n741), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(new_n796), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n853), .B1(new_n876), .B2(new_n855), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n852), .B1(new_n871), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(G141gat), .B1(new_n878), .B2(new_n519), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n851), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT123), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g681(.A(KEYINPUT123), .B(new_n852), .C1(new_n871), .C2(new_n877), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n882), .A2(new_n686), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n850), .B1(new_n884), .B2(G141gat), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT58), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n880), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT124), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n889), .B(new_n880), .C1(new_n885), .C2(new_n886), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(G1344gat));
  AND2_X1   g690(.A1(new_n882), .A2(new_n883), .ZN(new_n892));
  AOI211_X1 g691(.A(KEYINPUT59), .B(new_n288), .C1(new_n892), .C2(new_n619), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT57), .B1(new_n825), .B2(new_n374), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n593), .B1(new_n858), .B2(new_n816), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n622), .A2(new_n518), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n854), .B(new_n375), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n895), .A2(new_n852), .A3(new_n619), .A4(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n894), .B1(new_n899), .B2(G148gat), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n619), .A2(new_n288), .ZN(new_n901));
  OAI22_X1  g700(.A1(new_n893), .A2(new_n900), .B1(new_n849), .B2(new_n901), .ZN(G1345gat));
  AOI21_X1  g701(.A(new_n297), .B1(new_n892), .B2(new_n593), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n849), .A2(G155gat), .A3(new_n741), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n903), .A2(new_n904), .ZN(G1346gat));
  NOR2_X1   g704(.A1(new_n842), .A2(G162gat), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n848), .A2(new_n906), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n892), .A2(new_n674), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(new_n298), .ZN(G1347gat));
  AOI21_X1  g708(.A(new_n627), .B1(new_n388), .B2(new_n402), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n826), .A2(new_n438), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(G169gat), .B1(new_n911), .B2(new_n519), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT125), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n825), .A2(new_n627), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n634), .A3(new_n724), .ZN(new_n915));
  INV_X1    g714(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n232), .A3(new_n686), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n913), .A2(new_n917), .ZN(G1348gat));
  OAI21_X1  g717(.A(G176gat), .B1(new_n911), .B2(new_n620), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n619), .A2(new_n233), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n919), .B1(new_n915), .B2(new_n920), .ZN(G1349gat));
  NAND3_X1  g720(.A1(new_n916), .A2(new_n244), .A3(new_n593), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n220), .B1(new_n911), .B2(new_n741), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g725(.A(G190gat), .B1(new_n911), .B2(new_n557), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT61), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n916), .A2(new_n216), .A3(new_n674), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1351gat));
  NAND3_X1  g729(.A1(new_n724), .A2(new_n439), .A3(new_n375), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n931), .A2(new_n627), .A3(new_n825), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n933), .A2(new_n740), .ZN(new_n934));
  NAND4_X1  g733(.A1(new_n895), .A2(new_n439), .A3(new_n898), .A4(new_n910), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n518), .A2(G197gat), .ZN(new_n936));
  OAI22_X1  g735(.A1(new_n934), .A2(G197gat), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(G1352gat));
  OR3_X1    g737(.A1(new_n933), .A2(G204gat), .A3(new_n620), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n939), .A2(KEYINPUT62), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT127), .ZN(new_n941));
  OAI21_X1  g740(.A(G204gat), .B1(new_n935), .B2(new_n620), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n939), .A2(KEYINPUT62), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(G1353gat));
  OAI21_X1  g743(.A(G211gat), .B1(new_n935), .B2(new_n741), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT63), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n933), .A2(G211gat), .A3(new_n741), .ZN(new_n947));
  OR2_X1    g746(.A1(new_n946), .A2(new_n947), .ZN(G1354gat));
  OAI21_X1  g747(.A(G218gat), .B1(new_n935), .B2(new_n557), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n557), .A2(G218gat), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n933), .B2(new_n950), .ZN(G1355gat));
endmodule


