//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n209, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1270, new_n1271, new_n1272,
    new_n1274, new_n1275, new_n1276, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(KEYINPUT64), .A3(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  AOI21_X1  g0004(.A(KEYINPUT64), .B1(new_n201), .B2(new_n202), .ZN(new_n205));
  NOR3_X1   g0005(.A1(new_n204), .A2(G77), .A3(new_n205), .ZN(G353));
  INV_X1    g0006(.A(G97), .ZN(new_n207));
  INV_X1    g0007(.A(G107), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(G355));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G20), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G68), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  OAI221_X1 g0023(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  INV_X1    g0025(.A(G58), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  INV_X1    g0027(.A(G257), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n225), .B1(new_n226), .B2(new_n227), .C1(new_n207), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n211), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n214), .B1(new_n217), .B2(new_n218), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT65), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n227), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n236), .B(new_n240), .Z(G358));
  XNOR2_X1  g0041(.A(G87), .B(G97), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT82), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT3), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n252), .A2(G33), .ZN(new_n253));
  OAI21_X1  g0053(.A(G303), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n256));
  NAND4_X1  g0056(.A1(new_n255), .A2(new_n256), .A3(G264), .A4(G1698), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n255), .A2(new_n256), .A3(G257), .A4(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n254), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G1), .A3(G13), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G45), .ZN(new_n266));
  OR2_X1    g0066(.A1(KEYINPUT5), .A2(G41), .ZN(new_n267));
  NAND2_X1  g0067(.A1(KEYINPUT5), .A2(G41), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n270), .B1(new_n216), .B2(new_n261), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g0072(.A(KEYINPUT5), .B(G41), .ZN(new_n273));
  INV_X1    g0073(.A(new_n266), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n262), .ZN(new_n276));
  INV_X1    g0076(.A(G270), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n272), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n249), .B1(new_n264), .B2(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n269), .A2(new_n263), .ZN(new_n280));
  AOI22_X1  g0080(.A1(new_n280), .A2(G270), .B1(new_n271), .B2(new_n269), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n260), .A2(new_n263), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(KEYINPUT82), .A3(new_n282), .ZN(new_n283));
  NAND4_X1  g0083(.A1(new_n279), .A2(KEYINPUT21), .A3(G169), .A4(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n281), .A2(G179), .A3(new_n282), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  INV_X1    g0087(.A(G116), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n287), .A2(new_n215), .B1(G20), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n207), .A2(KEYINPUT79), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT79), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G97), .ZN(new_n292));
  AOI21_X1  g0092(.A(G33), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G283), .ZN(new_n294));
  INV_X1    g0094(.A(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(KEYINPUT20), .B(new_n289), .C1(new_n293), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(KEYINPUT83), .ZN(new_n298));
  XNOR2_X1  g0098(.A(KEYINPUT79), .B(G97), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n295), .B(new_n294), .C1(new_n299), .C2(G33), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT83), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n300), .A2(new_n301), .A3(KEYINPUT20), .A4(new_n289), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT20), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n290), .A2(new_n292), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n296), .B1(new_n304), .B2(new_n250), .ZN(new_n305));
  INV_X1    g0105(.A(new_n289), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n298), .A2(new_n302), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G13), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(G1), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G20), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n288), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n287), .A2(new_n215), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n314), .B(new_n311), .C1(G1), .C2(new_n250), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n312), .B1(new_n316), .B2(new_n288), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n308), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT84), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n308), .A2(new_n317), .A3(KEYINPUT84), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n286), .A2(new_n322), .A3(KEYINPUT85), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT85), .B1(new_n286), .B2(new_n322), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n279), .A2(G169), .A3(new_n283), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n326), .B1(new_n320), .B2(new_n321), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT86), .B1(new_n327), .B2(KEYINPUT21), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT86), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT21), .ZN(new_n330));
  INV_X1    g0130(.A(new_n321), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT84), .B1(new_n308), .B2(new_n317), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n329), .B(new_n330), .C1(new_n333), .C2(new_n326), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n328), .A2(new_n334), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n279), .A2(new_n283), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G200), .ZN(new_n337));
  INV_X1    g0137(.A(G190), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n333), .B(new_n337), .C1(new_n338), .C2(new_n336), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n325), .A2(new_n335), .A3(new_n339), .ZN(new_n340));
  NOR3_X1   g0140(.A1(new_n309), .A2(new_n295), .A3(G1), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n341), .A2(KEYINPUT25), .A3(new_n208), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(KEYINPUT25), .B1(new_n341), .B2(new_n208), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n315), .A2(new_n208), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n255), .A2(new_n256), .A3(new_n295), .A4(G87), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT87), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT22), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT3), .B(G33), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n351), .A2(new_n295), .A3(G87), .A4(new_n348), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT24), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G33), .A2(G116), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n355), .A2(G20), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT23), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n295), .B2(G107), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n208), .A2(KEYINPUT23), .A3(G20), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n356), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n353), .A2(new_n354), .A3(new_n360), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n354), .B1(new_n353), .B2(new_n360), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n313), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT88), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT88), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n366), .B(new_n313), .C1(new_n362), .C2(new_n363), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n345), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n351), .A2(G257), .A3(G1698), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n351), .A2(G250), .A3(new_n258), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G294), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n263), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT89), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n372), .A2(KEYINPUT89), .A3(new_n263), .ZN(new_n376));
  INV_X1    g0176(.A(new_n272), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(G264), .B2(new_n280), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n280), .A2(G264), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n373), .A2(new_n380), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n381), .A2(new_n377), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n379), .A2(G169), .B1(new_n382), .B2(G179), .ZN(new_n383));
  OR2_X1    g0183(.A1(new_n368), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(G179), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n377), .B1(G257), .B2(new_n280), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n255), .A2(new_n256), .A3(G250), .A4(G1698), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n294), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n255), .A2(new_n256), .A3(G244), .A4(new_n258), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT4), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT4), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n351), .A2(new_n391), .A3(G244), .A4(new_n258), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n388), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n263), .B1(new_n393), .B2(KEYINPUT80), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n390), .A2(new_n392), .ZN(new_n395));
  INV_X1    g0195(.A(new_n388), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT80), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n385), .B(new_n386), .C1(new_n394), .C2(new_n399), .ZN(new_n400));
  XOR2_X1   g0200(.A(G97), .B(G107), .Z(new_n401));
  NAND2_X1  g0201(.A1(new_n208), .A2(KEYINPUT6), .ZN(new_n402));
  OAI22_X1  g0202(.A1(new_n401), .A2(KEYINPUT6), .B1(new_n299), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G20), .ZN(new_n404));
  NOR2_X1   g0204(.A1(G20), .A2(G33), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G77), .ZN(new_n406));
  XOR2_X1   g0206(.A(new_n406), .B(KEYINPUT78), .Z(new_n407));
  NAND2_X1  g0207(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT72), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n250), .B2(KEYINPUT3), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n252), .A2(KEYINPUT72), .A3(G33), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n256), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT7), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n413), .A2(G20), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n413), .B1(new_n351), .B2(G20), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n208), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n313), .B1(new_n408), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n341), .A2(new_n207), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n315), .B2(new_n207), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n386), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n262), .B1(new_n397), .B2(new_n398), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n393), .A2(KEYINPUT80), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n400), .B(new_n422), .C1(new_n426), .C2(G169), .ZN(new_n427));
  OAI211_X1 g0227(.A(G190), .B(new_n386), .C1(new_n394), .C2(new_n399), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n415), .A2(new_n416), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n404), .B(new_n407), .C1(new_n429), .C2(new_n208), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n420), .B1(new_n430), .B2(new_n313), .ZN(new_n431));
  INV_X1    g0231(.A(G200), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n428), .B(new_n431), .C1(new_n426), .C2(new_n432), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n432), .B1(new_n381), .B2(new_n377), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(new_n379), .B2(G190), .ZN(new_n436));
  INV_X1    g0236(.A(new_n345), .ZN(new_n437));
  INV_X1    g0237(.A(new_n363), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n361), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n366), .B1(new_n439), .B2(new_n313), .ZN(new_n440));
  INV_X1    g0240(.A(new_n367), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n436), .B(new_n437), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  XNOR2_X1  g0242(.A(KEYINPUT15), .B(G87), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(new_n311), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n299), .A2(new_n222), .A3(new_n208), .ZN(new_n446));
  NAND2_X1  g0246(.A1(G33), .A2(G97), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT19), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n295), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n351), .A2(new_n295), .A3(G68), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n250), .A2(G20), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n448), .B1(new_n299), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n450), .A2(new_n451), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n445), .B1(new_n455), .B2(new_n313), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n316), .A2(new_n444), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n351), .A2(G244), .A3(G1698), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n351), .A2(new_n258), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n459), .B(new_n355), .C1(new_n460), .C2(new_n221), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n263), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n263), .A2(new_n223), .A3(new_n274), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n463), .B1(new_n271), .B2(new_n274), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(G179), .ZN(new_n466));
  AOI21_X1  g0266(.A(G169), .B1(new_n462), .B2(new_n464), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n458), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n465), .A2(new_n338), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n455), .A2(new_n313), .ZN(new_n470));
  INV_X1    g0270(.A(new_n445), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n316), .A2(G87), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n432), .B1(new_n462), .B2(new_n464), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n469), .B1(new_n475), .B2(KEYINPUT81), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT81), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n473), .B2(new_n474), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n468), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n384), .A2(new_n434), .A3(new_n442), .A4(new_n479), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n263), .B1(new_n351), .B2(G77), .ZN(new_n481));
  XNOR2_X1  g0281(.A(KEYINPUT66), .B(G223), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G1698), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(G222), .B2(G1698), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n481), .B1(new_n484), .B2(new_n351), .ZN(new_n485));
  INV_X1    g0285(.A(G41), .ZN(new_n486));
  INV_X1    g0286(.A(G45), .ZN(new_n487));
  AOI21_X1  g0287(.A(G1), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(new_n262), .A3(G274), .ZN(new_n489));
  INV_X1    g0289(.A(G226), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n262), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n489), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n485), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(G169), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n341), .A2(new_n202), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n341), .A2(new_n313), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n265), .A2(G20), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n497), .A2(G50), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n205), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n295), .B1(new_n500), .B2(new_n203), .ZN(new_n501));
  XNOR2_X1  g0301(.A(KEYINPUT8), .B(G58), .ZN(new_n502));
  INV_X1    g0302(.A(G150), .ZN(new_n503));
  INV_X1    g0303(.A(new_n405), .ZN(new_n504));
  OAI22_X1  g0304(.A1(new_n502), .A2(new_n453), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n313), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT67), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n496), .B(new_n499), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(new_n502), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n509), .A2(new_n452), .B1(G150), .B2(new_n405), .ZN(new_n510));
  OAI21_X1  g0310(.A(G20), .B1(new_n204), .B2(new_n205), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n314), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(KEYINPUT67), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  AOI211_X1 g0314(.A(new_n495), .B(new_n514), .C1(new_n385), .C2(new_n494), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n494), .A2(new_n432), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n485), .A2(new_n338), .A3(new_n493), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT10), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT9), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n499), .A2(new_n496), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n512), .B2(KEYINPUT67), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n506), .A2(new_n507), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR3_X1   g0324(.A1(new_n508), .A2(new_n513), .A3(KEYINPUT9), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n518), .B(new_n519), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n518), .B1(new_n525), .B2(new_n524), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT10), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n515), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n341), .A2(new_n220), .ZN(new_n530));
  XNOR2_X1  g0330(.A(new_n530), .B(KEYINPUT12), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n405), .A2(G50), .B1(G20), .B2(new_n220), .ZN(new_n532));
  INV_X1    g0332(.A(G77), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n532), .B1(new_n453), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(KEYINPUT11), .A3(new_n313), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n497), .A2(G68), .A3(new_n498), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n531), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT11), .B1(new_n534), .B2(new_n313), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT14), .ZN(new_n541));
  OAI22_X1  g0341(.A1(new_n489), .A2(KEYINPUT71), .B1(new_n492), .B2(new_n221), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT71), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(new_n271), .B2(new_n488), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT13), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT70), .ZN(new_n547));
  NOR2_X1   g0347(.A1(G226), .A2(G1698), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n227), .A2(G1698), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n549), .A2(new_n255), .A3(new_n256), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n447), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n547), .B1(new_n552), .B2(new_n263), .ZN(new_n553));
  AOI211_X1 g0353(.A(KEYINPUT70), .B(new_n262), .C1(new_n551), .C2(new_n447), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n545), .B(new_n546), .C1(new_n553), .C2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n548), .B1(new_n227), .B2(G1698), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n557), .A2(new_n351), .B1(G33), .B2(G97), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT70), .B1(new_n558), .B2(new_n262), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n552), .A2(new_n547), .A3(new_n263), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n546), .B1(new_n561), .B2(new_n545), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n541), .B(G169), .C1(new_n556), .C2(new_n562), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n545), .B1(new_n553), .B2(new_n554), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT13), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n565), .A2(G179), .A3(new_n555), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n555), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n541), .B1(new_n568), .B2(G169), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n540), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n556), .A2(new_n562), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n540), .B1(new_n571), .B2(G190), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n432), .B2(new_n571), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n351), .A2(G238), .A3(G1698), .ZN(new_n574));
  OAI221_X1 g0374(.A(new_n574), .B1(new_n208), .B2(new_n351), .C1(new_n460), .C2(new_n227), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n263), .ZN(new_n576));
  INV_X1    g0376(.A(new_n492), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n577), .A2(G244), .B1(new_n488), .B2(new_n271), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(G169), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT68), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n311), .B2(G77), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n341), .A2(KEYINPUT68), .A3(new_n533), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n533), .B1(new_n265), .B2(G20), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n582), .A2(new_n583), .B1(new_n497), .B2(new_n584), .ZN(new_n585));
  OAI22_X1  g0385(.A1(new_n502), .A2(new_n504), .B1(new_n295), .B2(new_n533), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n443), .A2(new_n453), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n313), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT69), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n585), .A2(new_n588), .A3(KEYINPUT69), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n579), .A2(new_n580), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n576), .A2(new_n385), .A3(new_n578), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n579), .A2(G200), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n576), .A2(G190), .A3(new_n578), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n596), .A2(new_n591), .A3(new_n592), .A4(new_n597), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n529), .A2(new_n570), .A3(new_n573), .A4(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT74), .ZN(new_n601));
  OR2_X1    g0401(.A1(G223), .A2(G1698), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n490), .A2(G1698), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n255), .A2(new_n602), .A3(new_n256), .A4(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(G33), .A2(G87), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n263), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n262), .A2(G232), .A3(new_n491), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n489), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n580), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n262), .B1(new_n604), .B2(new_n605), .ZN(new_n612));
  NOR3_X1   g0412(.A1(new_n612), .A2(new_n609), .A3(new_n385), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT16), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n220), .B1(new_n415), .B2(new_n416), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n226), .A2(new_n220), .ZN(new_n617));
  OAI21_X1  g0417(.A(G20), .B1(new_n617), .B2(new_n201), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n405), .A2(G159), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n615), .B1(new_n616), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n255), .A2(new_n256), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT7), .B1(new_n622), .B2(new_n295), .ZN(new_n623));
  AOI211_X1 g0423(.A(new_n413), .B(G20), .C1(new_n255), .C2(new_n256), .ZN(new_n624));
  OAI21_X1  g0424(.A(G68), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n620), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n625), .A2(KEYINPUT16), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n621), .A2(new_n627), .A3(new_n313), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n502), .B1(new_n265), .B2(G20), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n629), .A2(new_n497), .B1(new_n341), .B2(new_n502), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n614), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n601), .B1(new_n631), .B2(KEYINPUT18), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT18), .ZN(new_n633));
  INV_X1    g0433(.A(new_n630), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n622), .A2(KEYINPUT7), .A3(new_n295), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n416), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n620), .B1(new_n636), .B2(G68), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n314), .B1(new_n637), .B2(KEYINPUT16), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n634), .B1(new_n638), .B2(new_n621), .ZN(new_n639));
  OAI211_X1 g0439(.A(KEYINPUT74), .B(new_n633), .C1(new_n639), .C2(new_n614), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n632), .A2(new_n640), .ZN(new_n641));
  NOR4_X1   g0441(.A1(new_n639), .A2(KEYINPUT73), .A3(new_n633), .A4(new_n614), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT73), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n643), .B1(new_n631), .B2(KEYINPUT18), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT76), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n607), .A2(new_n610), .A3(new_n338), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n432), .B1(new_n612), .B2(new_n609), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n628), .A2(new_n646), .A3(new_n630), .A4(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT75), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n628), .A2(KEYINPUT75), .A3(new_n630), .A4(new_n649), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(KEYINPUT17), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n650), .A2(new_n651), .A3(KEYINPUT17), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n641), .A2(new_n645), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  OR3_X1    g0458(.A1(new_n600), .A2(new_n658), .A3(KEYINPUT77), .ZN(new_n659));
  OAI21_X1  g0459(.A(KEYINPUT77), .B1(new_n600), .B2(new_n658), .ZN(new_n660));
  AOI211_X1 g0460(.A(new_n340), .B(new_n480), .C1(new_n659), .C2(new_n660), .ZN(G372));
  NAND2_X1  g0461(.A1(new_n659), .A2(new_n660), .ZN(new_n662));
  INV_X1    g0462(.A(new_n442), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n427), .A2(new_n433), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n466), .A2(new_n467), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n456), .A2(new_n457), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n469), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n475), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n663), .A2(new_n664), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n286), .A2(new_n322), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n335), .A2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n384), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n427), .ZN(new_n676));
  XNOR2_X1  g0476(.A(KEYINPUT90), .B(KEYINPUT26), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n479), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT26), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n670), .B2(new_n427), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n468), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n675), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n662), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n631), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n633), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n631), .A2(KEYINPUT18), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT91), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n593), .A2(new_n689), .A3(new_n594), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n689), .B1(new_n593), .B2(new_n594), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT14), .B1(new_n571), .B2(new_n580), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(new_n566), .A3(new_n563), .ZN(new_n695));
  AOI22_X1  g0495(.A1(new_n693), .A2(new_n573), .B1(new_n695), .B2(new_n540), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n655), .A2(new_n656), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n688), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n528), .A2(new_n526), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n515), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n684), .A2(new_n701), .ZN(G369));
  INV_X1    g0502(.A(G330), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n310), .A2(new_n295), .ZN(new_n704));
  OR2_X1    g0504(.A1(new_n704), .A2(KEYINPUT27), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(KEYINPUT27), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n705), .A2(new_n706), .A3(G213), .ZN(new_n707));
  INV_X1    g0507(.A(G343), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n333), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g0511(.A1(new_n340), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n673), .A2(new_n711), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n703), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n442), .B1(new_n383), .B2(new_n368), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n368), .A2(new_n710), .ZN(new_n716));
  OAI22_X1  g0516(.A1(new_n715), .A2(new_n716), .B1(new_n384), .B2(new_n710), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n384), .A2(new_n709), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n325), .A2(new_n335), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n709), .ZN(new_n721));
  INV_X1    g0521(.A(new_n715), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n718), .A2(new_n723), .ZN(G399));
  NOR2_X1   g0524(.A1(new_n446), .A2(G116), .ZN(new_n725));
  INV_X1    g0525(.A(new_n212), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G41), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n725), .A2(new_n728), .A3(G1), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n729), .B1(new_n218), .B2(new_n728), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT28), .ZN(new_n731));
  INV_X1    g0531(.A(new_n474), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n732), .A2(KEYINPUT81), .A3(new_n456), .A4(new_n472), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n733), .A2(new_n478), .A3(new_n668), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(new_n667), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n715), .A2(new_n664), .A3(new_n735), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n720), .A2(new_n736), .A3(new_n339), .A4(new_n710), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n465), .A2(new_n285), .A3(new_n381), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(new_n426), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT30), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n738), .A2(new_n426), .A3(KEYINPUT30), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n373), .A2(new_n272), .A3(new_n380), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n336), .A2(new_n385), .A3(new_n743), .A4(new_n465), .ZN(new_n744));
  OAI211_X1 g0544(.A(new_n741), .B(new_n742), .C1(new_n744), .C2(new_n426), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n745), .A2(KEYINPUT31), .A3(new_n709), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT31), .B1(new_n745), .B2(new_n709), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n703), .B1(new_n737), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n325), .A2(new_n335), .A3(new_n384), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT92), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n325), .A2(new_n335), .A3(KEYINPUT92), .A4(new_n384), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n753), .A2(new_n671), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n677), .B1(new_n735), .B2(new_n427), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n676), .A2(KEYINPUT26), .A3(new_n667), .A4(new_n669), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n468), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n759), .A2(KEYINPUT29), .A3(new_n710), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n709), .B1(new_n675), .B2(new_n682), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n761), .A2(KEYINPUT29), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n750), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n731), .B1(new_n763), .B2(G1), .ZN(G364));
  NOR2_X1   g0564(.A1(new_n309), .A2(G20), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n265), .B1(new_n765), .B2(G45), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n727), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n714), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n712), .A2(new_n703), .A3(new_n713), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G13), .A2(G33), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n712), .A2(new_n713), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n215), .B1(G20), .B2(new_n580), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n247), .A2(G45), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT93), .Z(new_n780));
  NOR2_X1   g0580(.A1(new_n726), .A2(new_n351), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n780), .B(new_n781), .C1(G45), .C2(new_n218), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n726), .A2(new_n622), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n783), .A2(G355), .B1(new_n288), .B2(new_n726), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n778), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n776), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n295), .A2(G179), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n787), .A2(G190), .A3(G200), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n222), .ZN(new_n789));
  NOR2_X1   g0589(.A1(G190), .A2(G200), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G159), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(KEYINPUT32), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n338), .A2(G179), .A3(G200), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n295), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n789), .B(new_n794), .C1(G97), .C2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n787), .A2(new_n338), .A3(G200), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n799), .A2(KEYINPUT94), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(KEYINPUT94), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G107), .ZN(new_n804));
  NAND2_X1  g0604(.A1(G20), .A2(G179), .ZN(new_n805));
  NOR3_X1   g0605(.A1(new_n805), .A2(new_n338), .A3(new_n432), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n805), .A2(new_n432), .A3(G190), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n807), .A2(new_n202), .B1(new_n809), .B2(new_n220), .ZN(new_n810));
  INV_X1    g0610(.A(new_n805), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n790), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n810), .B1(G77), .B2(new_n813), .ZN(new_n814));
  NOR3_X1   g0614(.A1(new_n805), .A2(new_n338), .A3(G200), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n351), .B1(new_n816), .B2(new_n226), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(KEYINPUT32), .B2(new_n793), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n798), .A2(new_n804), .A3(new_n814), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n803), .A2(G283), .ZN(new_n820));
  INV_X1    g0620(.A(G311), .ZN(new_n821));
  INV_X1    g0621(.A(G294), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n622), .B1(new_n812), .B2(new_n821), .C1(new_n796), .C2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n788), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n823), .B1(G303), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(KEYINPUT33), .B(G317), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n808), .A2(new_n826), .B1(new_n806), .B2(G326), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n792), .A2(G329), .B1(new_n815), .B2(G322), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n820), .A2(new_n825), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n786), .B1(new_n819), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n768), .ZN(new_n831));
  NOR3_X1   g0631(.A1(new_n785), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n775), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n771), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(G396));
  AOI21_X1  g0635(.A(new_n710), .B1(new_n591), .B2(new_n592), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  AND3_X1   g0637(.A1(new_n595), .A2(new_n598), .A3(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n692), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n840), .A2(new_n690), .A3(new_n836), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n761), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n434), .A2(new_n442), .A3(new_n667), .A4(new_n669), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n328), .A2(new_n334), .B1(new_n322), .B2(new_n286), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n844), .B1(new_n384), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n679), .A2(new_n681), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n667), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n710), .B(new_n842), .C1(new_n846), .C2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n843), .A2(new_n750), .A3(new_n849), .ZN(new_n850));
  NOR3_X1   g0650(.A1(new_n340), .A2(new_n480), .A3(new_n709), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n745), .A2(new_n709), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT31), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n746), .ZN(new_n855));
  OAI21_X1  g0655(.A(G330), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n849), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n761), .A2(new_n842), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n856), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n850), .A2(new_n859), .A3(new_n831), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n776), .A2(new_n772), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT95), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n831), .B1(new_n863), .B2(new_n533), .ZN(new_n864));
  INV_X1    g0664(.A(G283), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n809), .A2(new_n865), .B1(new_n812), .B2(new_n288), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT96), .ZN(new_n867));
  INV_X1    g0667(.A(G303), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n866), .A2(new_n867), .B1(new_n868), .B2(new_n807), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n867), .B2(new_n866), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT97), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n803), .A2(G87), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n622), .B1(new_n816), .B2(new_n822), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(G311), .B2(new_n792), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n797), .A2(G97), .B1(new_n824), .B2(G107), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n871), .A2(new_n872), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n813), .A2(G159), .B1(G150), .B2(new_n808), .ZN(new_n877));
  INV_X1    g0677(.A(G137), .ZN(new_n878));
  XOR2_X1   g0678(.A(KEYINPUT98), .B(G143), .Z(new_n879));
  OAI221_X1 g0679(.A(new_n877), .B1(new_n878), .B2(new_n807), .C1(new_n816), .C2(new_n879), .ZN(new_n880));
  XOR2_X1   g0680(.A(KEYINPUT99), .B(KEYINPUT34), .Z(new_n881));
  XNOR2_X1  g0681(.A(new_n880), .B(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n803), .A2(G68), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n788), .A2(new_n202), .ZN(new_n884));
  INV_X1    g0684(.A(G132), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n351), .B1(new_n791), .B2(new_n885), .ZN(new_n886));
  AOI211_X1 g0686(.A(new_n884), .B(new_n886), .C1(G58), .C2(new_n797), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n882), .A2(new_n883), .A3(new_n887), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n876), .A2(new_n888), .ZN(new_n889));
  OAI221_X1 g0689(.A(new_n864), .B1(new_n889), .B2(new_n786), .C1(new_n842), .C2(new_n773), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n860), .A2(new_n890), .ZN(G384));
  AOI211_X1 g0691(.A(new_n288), .B(new_n217), .C1(new_n403), .C2(KEYINPUT35), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(KEYINPUT35), .B2(new_n403), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n893), .B(KEYINPUT36), .ZN(new_n894));
  OAI21_X1  g0694(.A(G77), .B1(new_n226), .B2(new_n220), .ZN(new_n895));
  OAI22_X1  g0695(.A1(new_n895), .A2(new_n218), .B1(G50), .B2(new_n220), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(G1), .A3(new_n309), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT100), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n628), .A2(new_n630), .A3(new_n649), .ZN(new_n900));
  OR2_X1    g0700(.A1(new_n637), .A2(KEYINPUT16), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n634), .B1(new_n901), .B2(new_n638), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n900), .B1(new_n902), .B2(new_n707), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n614), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT37), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n628), .A2(new_n630), .ZN(new_n906));
  INV_X1    g0706(.A(new_n707), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT37), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n685), .A2(new_n908), .A3(new_n909), .A4(new_n900), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n902), .A2(new_n707), .ZN(new_n912));
  OAI211_X1 g0712(.A(KEYINPUT38), .B(new_n911), .C1(new_n657), .C2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT38), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n900), .B1(new_n639), .B2(new_n614), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n639), .A2(new_n707), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT37), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(KEYINPUT101), .A3(new_n910), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT101), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n919), .B(KEYINPUT37), .C1(new_n915), .C2(new_n916), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n908), .B1(new_n697), .B2(new_n688), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n914), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT102), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n913), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n924), .B1(new_n913), .B2(new_n923), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n838), .B1(new_n693), .B2(new_n836), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n540), .A2(new_n709), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n570), .A2(new_n573), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n571), .A2(new_n432), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n539), .B1(new_n568), .B2(new_n338), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n540), .B(new_n709), .C1(new_n695), .C2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n928), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n935), .B(KEYINPUT40), .C1(new_n851), .C2(new_n855), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT40), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n687), .A2(KEYINPUT73), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n631), .A2(new_n643), .A3(KEYINPUT18), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n939), .A2(new_n632), .A3(new_n640), .A4(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n912), .B1(new_n941), .B2(new_n697), .ZN(new_n942));
  INV_X1    g0742(.A(new_n911), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n914), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n913), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n737), .A2(new_n749), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n945), .A2(new_n946), .A3(new_n935), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n927), .A2(new_n937), .B1(new_n938), .B2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n662), .A2(new_n946), .ZN(new_n950));
  OAI21_X1  g0750(.A(G330), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n950), .B2(new_n949), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT39), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n918), .A2(new_n920), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n697), .A2(new_n688), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n916), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT38), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n942), .A2(new_n943), .A3(new_n914), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n953), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n695), .A2(new_n540), .A3(new_n710), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n959), .B(new_n961), .C1(new_n953), .C2(new_n945), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n595), .A2(new_n709), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n849), .A2(new_n964), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n570), .A2(new_n573), .A3(new_n929), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n929), .B1(new_n570), .B2(new_n573), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n965), .A2(new_n945), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n686), .A2(new_n687), .A3(new_n707), .ZN(new_n971));
  AND3_X1   g0771(.A1(new_n962), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n760), .A2(new_n762), .A3(new_n662), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n701), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n972), .B(new_n974), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n952), .A2(new_n975), .B1(new_n265), .B2(new_n765), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n952), .A2(new_n975), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n899), .B1(new_n976), .B2(new_n977), .ZN(G367));
  NOR2_X1   g0778(.A1(new_n796), .A2(new_n220), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n351), .B1(new_n816), .B2(new_n503), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n979), .B(new_n980), .C1(G58), .C2(new_n824), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n803), .A2(G77), .ZN(new_n982));
  INV_X1    g0782(.A(new_n879), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n983), .A2(new_n806), .B1(G159), .B2(new_n808), .ZN(new_n984));
  AOI22_X1  g0784(.A1(G137), .A2(new_n792), .B1(new_n813), .B2(G50), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n981), .A2(new_n982), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n622), .B1(new_n812), .B2(new_n865), .ZN(new_n987));
  INV_X1    g0787(.A(G317), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n809), .A2(new_n822), .B1(new_n988), .B2(new_n791), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n987), .B(new_n989), .C1(G107), .C2(new_n797), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT46), .ZN(new_n991));
  AOI21_X1  g0791(.A(KEYINPUT110), .B1(new_n824), .B2(G116), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI22_X1  g0793(.A1(G311), .A2(new_n806), .B1(new_n815), .B2(G303), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT109), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n992), .A2(new_n991), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n995), .B(new_n996), .C1(new_n299), .C2(new_n802), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n986), .B1(new_n993), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT111), .Z(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT47), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(new_n786), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n777), .B1(new_n212), .B2(new_n443), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1002), .B1(new_n236), .B2(new_n781), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT108), .Z(new_n1004));
  NOR3_X1   g0804(.A1(new_n1001), .A2(new_n831), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n473), .A2(new_n709), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT103), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1007), .A2(new_n468), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n670), .B2(new_n1007), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n1005), .A2(KEYINPUT112), .B1(new_n774), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(KEYINPUT112), .B2(new_n1005), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n727), .B(new_n1013), .Z(new_n1014));
  INV_X1    g0814(.A(new_n718), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n434), .B1(new_n431), .B2(new_n710), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n676), .A2(new_n709), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n723), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT45), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n723), .A2(KEYINPUT45), .A3(new_n1018), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g0823(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  OR3_X1    g0825(.A1(new_n723), .A2(new_n1018), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1025), .B1(new_n723), .B2(new_n1018), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1015), .B1(new_n1023), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n721), .A2(new_n722), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n717), .B2(new_n721), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(new_n714), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n1032), .A2(new_n763), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1034), .A2(new_n718), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1029), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1014), .B1(new_n1036), .B2(new_n763), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n766), .B(KEYINPUT107), .Z(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1018), .ZN(new_n1041));
  OR3_X1    g0841(.A1(new_n718), .A2(KEYINPUT104), .A3(new_n1041), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1009), .A2(KEYINPUT43), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(KEYINPUT104), .B1(new_n718), .B2(new_n1041), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1042), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n721), .A2(new_n722), .A3(new_n1018), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n427), .B1(new_n1016), .B2(new_n384), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1048), .A2(KEYINPUT42), .B1(new_n710), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(KEYINPUT42), .B2(new_n1048), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1009), .A2(KEYINPUT43), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1044), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1054));
  OR3_X1    g0854(.A1(new_n1047), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1053), .B1(new_n1047), .B2(new_n1054), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1012), .B1(new_n1040), .B2(new_n1057), .ZN(G387));
  OAI21_X1  g0858(.A(new_n781), .B1(new_n240), .B2(new_n487), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n783), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1059), .B1(new_n725), .B2(new_n1060), .ZN(new_n1061));
  OR3_X1    g0861(.A1(new_n502), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1062));
  AOI21_X1  g0862(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1063));
  OAI21_X1  g0863(.A(KEYINPUT50), .B1(new_n502), .B2(G50), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n725), .A2(new_n1062), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n1061), .A2(new_n1065), .B1(new_n208), .B2(new_n726), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n768), .B1(new_n1066), .B2(new_n778), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n816), .A2(new_n988), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n809), .A2(new_n821), .B1(new_n812), .B2(new_n868), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1068), .B(new_n1069), .C1(G322), .C2(new_n806), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n1070), .A2(KEYINPUT48), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1070), .A2(KEYINPUT48), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n796), .A2(new_n865), .B1(new_n788), .B2(new_n822), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n1071), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1074), .A2(KEYINPUT49), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(KEYINPUT49), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n803), .A2(G116), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n351), .B1(new_n792), .B2(G326), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n622), .B1(new_n792), .B2(G150), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1080), .B1(new_n533), .B2(new_n788), .C1(new_n802), .C2(new_n207), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT113), .Z(new_n1082));
  NAND2_X1  g0882(.A1(new_n797), .A2(new_n444), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n509), .A2(new_n808), .B1(new_n815), .B2(G50), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n813), .A2(G68), .B1(new_n806), .B2(G159), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n786), .B1(new_n1079), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n717), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1067), .B(new_n1087), .C1(new_n1088), .C2(new_n774), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(new_n1032), .B2(new_n1039), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1032), .A2(new_n763), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n727), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1032), .A2(new_n763), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1090), .B1(new_n1092), .B2(new_n1093), .ZN(G393));
  AND2_X1   g0894(.A1(new_n1036), .A2(new_n727), .ZN(new_n1095));
  AND2_X1   g0895(.A1(new_n1029), .A2(new_n1035), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1095), .B1(new_n1033), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1041), .A2(new_n774), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n777), .B1(new_n212), .B2(new_n299), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(new_n244), .B2(new_n781), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(G317), .A2(new_n806), .B1(new_n815), .B2(G311), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT52), .Z(new_n1102));
  OAI21_X1  g0902(.A(new_n622), .B1(new_n812), .B2(new_n822), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n809), .A2(new_n868), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n1103), .B(new_n1104), .C1(G322), .C2(new_n792), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n797), .A2(G116), .B1(new_n824), .B2(G283), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1102), .A2(new_n804), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G150), .A2(new_n806), .B1(new_n815), .B2(G159), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT51), .Z(new_n1109));
  AOI22_X1  g0909(.A1(new_n792), .A2(new_n983), .B1(new_n824), .B2(G68), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(KEYINPUT114), .ZN(new_n1111));
  OR2_X1    g0911(.A1(new_n1110), .A2(KEYINPUT114), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1109), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n797), .A2(G77), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n808), .A2(G50), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n622), .B1(new_n813), .B2(new_n509), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n872), .A2(new_n1114), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1107), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n831), .B(new_n1100), .C1(new_n1118), .C2(new_n776), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1096), .A2(new_n1039), .B1(new_n1098), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1097), .A2(new_n1120), .ZN(G390));
  AOI21_X1  g0921(.A(new_n968), .B1(new_n849), .B2(new_n964), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n945), .A2(new_n953), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT39), .B1(new_n913), .B2(new_n923), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1122), .A2(new_n961), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n759), .A2(new_n710), .A3(new_n842), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n968), .B1(new_n1126), .B2(new_n964), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n927), .A2(new_n960), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1125), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n750), .A2(new_n842), .A3(new_n969), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1129), .B1(KEYINPUT115), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n662), .A2(new_n750), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n973), .A2(new_n701), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1130), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n969), .B1(new_n750), .B2(new_n842), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n965), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n709), .B1(new_n755), .B2(new_n758), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n963), .B1(new_n1137), .B2(new_n842), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n968), .B1(new_n856), .B2(new_n928), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1138), .A2(new_n1130), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1133), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1130), .A2(KEYINPUT115), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1125), .B(new_n1143), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1131), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1144), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n960), .B(new_n927), .C1(new_n1138), .C2(new_n968), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1143), .B1(new_n1147), .B2(new_n1125), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1141), .B1(new_n1146), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1145), .A2(new_n727), .A3(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n768), .B1(new_n862), .B2(new_n509), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1152), .A2(new_n773), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n809), .A2(new_n878), .ZN(new_n1154));
  INV_X1    g0954(.A(G128), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n807), .A2(new_n1155), .B1(new_n816), .B2(new_n885), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1154), .B(new_n1156), .C1(G125), .C2(new_n792), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n803), .A2(G50), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT54), .B(G143), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n351), .B1(new_n812), .B2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(G159), .B2(new_n797), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n788), .A2(new_n503), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(new_n1162), .B(KEYINPUT53), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1157), .A2(new_n1158), .A3(new_n1161), .A4(new_n1163), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n813), .A2(new_n304), .B1(G283), .B2(new_n806), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n208), .B2(new_n809), .ZN(new_n1166));
  XOR2_X1   g0966(.A(new_n1166), .B(KEYINPUT116), .Z(new_n1167));
  AOI22_X1  g0967(.A1(new_n792), .A2(G294), .B1(new_n815), .B2(G116), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1167), .A2(new_n883), .A3(new_n1114), .A4(new_n1168), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n789), .A2(new_n351), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT117), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1164), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1151), .B(new_n1153), .C1(new_n776), .C2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1131), .A2(new_n1144), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1173), .B1(new_n1174), .B2(new_n1039), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1150), .A2(new_n1175), .ZN(G378));
  INV_X1    g0976(.A(KEYINPUT121), .ZN(new_n1177));
  OAI21_X1  g0977(.A(KEYINPUT102), .B1(new_n957), .B2(new_n958), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n842), .B1(new_n966), .B2(new_n967), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(new_n737), .B2(new_n749), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n913), .A2(new_n923), .A3(new_n924), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1178), .A2(new_n1180), .A3(KEYINPUT40), .A4(new_n1181), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n944), .A2(new_n913), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n935), .B1(new_n851), .B2(new_n855), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n938), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1182), .A2(G330), .A3(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n514), .A2(new_n707), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n529), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n529), .A2(new_n1188), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1192), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1186), .A2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1195), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1182), .A2(new_n1197), .A3(G330), .A4(new_n1185), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1196), .A2(new_n972), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n972), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1177), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n972), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1197), .B1(new_n948), .B2(G330), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1198), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1202), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1196), .A2(new_n972), .A3(new_n1198), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1205), .A2(KEYINPUT121), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1201), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1133), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1149), .A2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(KEYINPUT57), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1136), .A2(new_n1140), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1133), .B1(new_n1174), .B2(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(KEYINPUT57), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n727), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1211), .A2(new_n1215), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n351), .A2(G41), .ZN(new_n1217));
  AOI211_X1 g1017(.A(G50), .B(new_n1217), .C1(new_n250), .C2(new_n486), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n792), .A2(G283), .B1(new_n808), .B2(G97), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n443), .B2(new_n812), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n807), .A2(new_n288), .B1(new_n816), .B2(new_n208), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1220), .A2(new_n979), .A3(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1217), .B1(new_n533), .B2(new_n788), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT118), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n803), .A2(G58), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1222), .A2(new_n1224), .A3(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT58), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1218), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n797), .A2(G150), .B1(G125), .B2(new_n806), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT120), .Z(new_n1230));
  AOI22_X1  g1030(.A1(new_n813), .A2(G137), .B1(G132), .B2(new_n808), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1231), .B1(new_n1155), .B2(new_n816), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT119), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n788), .A2(new_n1159), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1232), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  OAI211_X1 g1035(.A(new_n1230), .B(new_n1235), .C1(new_n1233), .C2(new_n1234), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT59), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n803), .A2(G159), .ZN(new_n1238));
  AOI211_X1 g1038(.A(G33), .B(G41), .C1(new_n792), .C2(G124), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1236), .A2(KEYINPUT59), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1228), .B1(new_n1227), .B2(new_n1226), .C1(new_n1240), .C2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n776), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n831), .B1(new_n202), .B2(new_n861), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1243), .B(new_n1244), .C1(new_n1197), .C2(new_n773), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n1208), .B2(new_n1039), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1216), .A2(new_n1247), .ZN(G375));
  OAI21_X1  g1048(.A(new_n768), .B1(new_n862), .B2(G68), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n969), .A2(new_n773), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n351), .B1(new_n791), .B2(new_n1155), .C1(new_n796), .C2(new_n202), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(G159), .B2(new_n824), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n807), .A2(new_n885), .B1(new_n809), .B2(new_n1159), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n816), .A2(new_n878), .B1(new_n812), .B2(new_n503), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1225), .A2(new_n1252), .A3(new_n1255), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n816), .A2(new_n865), .B1(new_n812), .B2(new_n208), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1257), .B1(G116), .B2(new_n808), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n351), .B1(new_n806), .B2(G294), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n982), .A2(new_n1083), .A3(new_n1258), .A4(new_n1259), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n788), .A2(new_n207), .B1(new_n791), .B2(new_n868), .ZN(new_n1261));
  XOR2_X1   g1061(.A(new_n1261), .B(KEYINPUT122), .Z(new_n1262));
  OAI21_X1  g1062(.A(new_n1256), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1263));
  AOI211_X1 g1063(.A(new_n1249), .B(new_n1250), .C1(new_n776), .C2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n1212), .B2(new_n1039), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1014), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1142), .A2(new_n1266), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1209), .A2(new_n1212), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1265), .B1(new_n1267), .B2(new_n1268), .ZN(G381));
  OR4_X1    g1069(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1270), .A2(G387), .A3(G381), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1150), .A2(new_n1175), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1271), .A2(new_n1272), .A3(new_n1216), .A4(new_n1247), .ZN(G407));
  NAND2_X1  g1073(.A1(new_n708), .A2(G213), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1272), .A2(new_n1275), .ZN(new_n1276));
  OAI211_X1 g1076(.A(G407), .B(G213), .C1(G375), .C2(new_n1276), .ZN(G409));
  INV_X1    g1077(.A(G390), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(G393), .B(G396), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(G387), .B2(KEYINPUT126), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1055), .B(new_n1056), .C1(new_n1037), .C2(new_n1039), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1279), .B1(new_n1282), .B2(new_n1012), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1278), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(G387), .A2(new_n1280), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT126), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1286), .B1(new_n1282), .B2(new_n1012), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1285), .B(G390), .C1(new_n1280), .C2(new_n1287), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1284), .A2(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(G378), .B(new_n1247), .C1(new_n1211), .C2(new_n1215), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1199), .A2(new_n1200), .A3(new_n1177), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT121), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1292));
  OAI211_X1 g1092(.A(new_n1266), .B(new_n1210), .C1(new_n1291), .C2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1246), .B1(new_n1294), .B2(new_n1039), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1272), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1290), .A2(new_n1297), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1133), .A2(new_n1136), .A3(KEYINPUT60), .A4(new_n1140), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT123), .ZN(new_n1300));
  AOI22_X1  g1100(.A1(new_n1139), .A2(new_n1130), .B1(new_n849), .B2(new_n964), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1301), .B1(new_n1302), .B2(new_n1138), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT123), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1303), .A2(new_n1304), .A3(KEYINPUT60), .A4(new_n1133), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT60), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1306), .B1(new_n1209), .B2(new_n1212), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n728), .B1(new_n1209), .B2(new_n1212), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1300), .A2(new_n1305), .A3(new_n1307), .A4(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n860), .A2(KEYINPUT124), .A3(new_n890), .ZN(new_n1310));
  AND2_X1   g1110(.A1(new_n1265), .A2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1309), .A2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT124), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(G384), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1312), .A2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1309), .A2(new_n1311), .A3(new_n1314), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  AND4_X1   g1118(.A1(KEYINPUT63), .A2(new_n1298), .A3(new_n1274), .A4(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1275), .B1(new_n1290), .B2(new_n1297), .ZN(new_n1320));
  AOI21_X1  g1120(.A(KEYINPUT63), .B1(new_n1320), .B2(new_n1318), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1319), .A2(new_n1321), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1309), .A2(new_n1311), .A3(new_n1314), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1314), .B1(new_n1309), .B2(new_n1311), .ZN(new_n1324));
  INV_X1    g1124(.A(G2897), .ZN(new_n1325));
  OAI22_X1  g1125(.A1(new_n1323), .A2(new_n1324), .B1(new_n1325), .B2(new_n1274), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1274), .A2(new_n1325), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1316), .A2(new_n1327), .A3(new_n1317), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1326), .A2(new_n1328), .ZN(new_n1329));
  AOI22_X1  g1129(.A1(new_n1298), .A2(new_n1274), .B1(new_n1329), .B2(KEYINPUT125), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT125), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1326), .A2(new_n1328), .A3(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(KEYINPUT61), .B1(new_n1330), .B2(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1289), .B1(new_n1322), .B2(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1298), .A2(new_n1274), .A3(new_n1318), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(KEYINPUT62), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT62), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1320), .A2(new_n1337), .A3(new_n1318), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1336), .A2(new_n1289), .A3(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1298), .A2(new_n1274), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1329), .A2(KEYINPUT125), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1340), .A2(new_n1332), .A3(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT61), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1339), .A2(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(KEYINPUT127), .B1(new_n1334), .B2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1289), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT63), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1335), .A2(new_n1348), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1320), .A2(KEYINPUT63), .A3(new_n1318), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1347), .B1(new_n1344), .B2(new_n1351), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT127), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1333), .A2(new_n1289), .A3(new_n1336), .A4(new_n1338), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1352), .A2(new_n1353), .A3(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1346), .A2(new_n1355), .ZN(G405));
  NAND2_X1  g1156(.A1(G375), .A2(new_n1272), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1357), .A2(new_n1290), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1358), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1357), .A2(new_n1318), .A3(new_n1290), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1359), .A2(new_n1360), .ZN(new_n1361));
  XNOR2_X1  g1161(.A(new_n1361), .B(new_n1347), .ZN(G402));
endmodule


