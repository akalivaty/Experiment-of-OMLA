//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n445, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n553, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n607, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1146, new_n1147, new_n1148;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT66), .ZN(new_n455));
  NOR4_X1   g030(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT2), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G325));
  XOR2_X1   g034(.A(new_n458), .B(KEYINPUT67), .Z(G261));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2106), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g040(.A(new_n465), .B(KEYINPUT68), .ZN(G319));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  AND3_X1   g042(.A1(new_n467), .A2(KEYINPUT70), .A3(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(KEYINPUT70), .B1(new_n467), .B2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(G101), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n471), .B1(new_n472), .B2(KEYINPUT3), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n472), .A2(KEYINPUT3), .ZN(new_n476));
  NAND4_X1  g051(.A1(new_n473), .A2(new_n475), .A3(new_n467), .A4(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G137), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n470), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  XNOR2_X1  g054(.A(KEYINPUT3), .B(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G125), .ZN(new_n481));
  NAND2_X1  g056(.A1(G113), .A2(G2104), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n467), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n479), .A2(new_n483), .ZN(G160));
  NAND4_X1  g059(.A1(new_n473), .A2(new_n475), .A3(G2105), .A4(new_n476), .ZN(new_n485));
  INV_X1    g060(.A(G124), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n467), .A2(G112), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n488));
  OAI22_X1  g063(.A1(new_n485), .A2(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n477), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(G136), .B2(new_n490), .ZN(G162));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n473), .A2(new_n475), .A3(new_n493), .A4(new_n476), .ZN(new_n494));
  NOR3_X1   g069(.A1(new_n492), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n494), .A2(KEYINPUT4), .B1(new_n480), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  AND3_X1   g074(.A1(new_n499), .A2(KEYINPUT71), .A3(G2105), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT71), .B1(new_n499), .B2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n498), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AND2_X1   g077(.A1(G126), .A2(G2105), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n473), .A2(new_n475), .A3(new_n476), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT72), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n502), .A2(new_n507), .A3(new_n504), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n496), .B1(new_n506), .B2(new_n508), .ZN(G164));
  NAND2_X1  g084(.A1(KEYINPUT73), .A2(G543), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  XNOR2_X1  g086(.A(new_n510), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g087(.A(KEYINPUT6), .B(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n513), .A2(G543), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n512), .A2(G62), .ZN(new_n520));
  NAND2_X1  g095(.A1(G75), .A2(G543), .ZN(new_n521));
  XOR2_X1   g096(.A(new_n521), .B(KEYINPUT74), .Z(new_n522));
  AOI21_X1  g097(.A(new_n519), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n518), .A2(new_n523), .ZN(G166));
  INV_X1    g099(.A(new_n514), .ZN(new_n525));
  AND2_X1   g100(.A1(new_n525), .A2(G89), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n512), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  OAI211_X1 g105(.A(new_n527), .B(new_n529), .C1(new_n517), .C2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n526), .A2(new_n531), .ZN(G168));
  AOI22_X1  g107(.A1(new_n512), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n519), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT75), .B(G90), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n514), .A2(new_n535), .B1(new_n536), .B2(new_n517), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(G171));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n510), .B(KEYINPUT5), .ZN(new_n540));
  INV_X1    g115(.A(G56), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT76), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n519), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n544), .B1(new_n543), .B2(new_n542), .ZN(new_n545));
  INV_X1    g120(.A(new_n517), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n525), .A2(G81), .B1(G43), .B2(new_n546), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT77), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(new_n546), .A2(G53), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n525), .A2(G91), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT78), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n540), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n556), .A2(new_n557), .A3(new_n562), .ZN(G299));
  NAND2_X1  g138(.A1(G171), .A2(KEYINPUT79), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n565), .B1(new_n534), .B2(new_n537), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G301));
  INV_X1    g143(.A(G168), .ZN(G286));
  INV_X1    g144(.A(G166), .ZN(G303));
  AOI22_X1  g145(.A1(new_n525), .A2(G87), .B1(G49), .B2(new_n546), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(G288));
  AOI22_X1  g148(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n574), .A2(new_n519), .ZN(new_n575));
  INV_X1    g150(.A(G86), .ZN(new_n576));
  INV_X1    g151(.A(G48), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n514), .A2(new_n576), .B1(new_n577), .B2(new_n517), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G305));
  AOI22_X1  g155(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n581), .A2(new_n519), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n525), .A2(G85), .B1(G47), .B2(new_n546), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n583), .A2(new_n584), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n582), .B1(new_n586), .B2(new_n587), .ZN(G290));
  AND3_X1   g163(.A1(new_n512), .A2(G92), .A3(new_n513), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT81), .Z(new_n590));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n589), .B(KEYINPUT81), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(KEYINPUT10), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n540), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(new_n546), .B2(G54), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n592), .A2(new_n594), .A3(new_n598), .ZN(new_n599));
  MUX2_X1   g174(.A(new_n599), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g175(.A(new_n599), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g176(.A1(G286), .A2(G868), .ZN(new_n602));
  INV_X1    g177(.A(G299), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(G868), .ZN(G297));
  OAI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(G868), .ZN(G280));
  AND3_X1   g180(.A1(new_n592), .A2(new_n594), .A3(new_n598), .ZN(new_n606));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g187(.A(new_n480), .B1(new_n468), .B2(new_n469), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2100), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT82), .B(KEYINPUT13), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT83), .ZN(new_n619));
  INV_X1    g194(.A(G111), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n618), .A2(new_n619), .B1(new_n620), .B2(G2105), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n619), .B2(new_n618), .ZN(new_n622));
  INV_X1    g197(.A(G123), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n485), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(G135), .B2(new_n490), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT84), .B(G2096), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n617), .A2(new_n627), .ZN(G156));
  XNOR2_X1  g203(.A(G1341), .B(G1348), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT15), .B(G2435), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2427), .B(G2430), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT85), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n631), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  AND3_X1   g217(.A1(new_n642), .A2(KEYINPUT86), .A3(new_n629), .ZN(new_n643));
  AOI21_X1  g218(.A(KEYINPUT86), .B1(new_n642), .B2(new_n629), .ZN(new_n644));
  OAI221_X1 g219(.A(G14), .B1(new_n629), .B2(new_n642), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(KEYINPUT87), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(G401));
  XNOR2_X1  g223(.A(G2084), .B(G2090), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT88), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AND2_X1   g227(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  AOI21_X1  g229(.A(KEYINPUT18), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2100), .ZN(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  AOI21_X1  g232(.A(new_n657), .B1(new_n652), .B2(KEYINPUT18), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(G2096), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n656), .B(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(G1971), .B(G1976), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  AND2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT20), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n663), .A2(new_n664), .ZN(new_n668));
  NOR3_X1   g243(.A1(new_n662), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n662), .B2(new_n668), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT89), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT90), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G229));
  INV_X1    g254(.A(G29), .ZN(new_n680));
  NOR2_X1   g255(.A1(G164), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(G27), .B2(new_n680), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n682), .A2(new_n443), .ZN(new_n683));
  INV_X1    g258(.A(G139), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n477), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT96), .ZN(new_n686));
  NAND2_X1  g261(.A1(G115), .A2(G2104), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n474), .A2(G2104), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n476), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G127), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n687), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT25), .ZN(new_n692));
  NAND2_X1  g267(.A1(G103), .A2(G2104), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n692), .B1(new_n693), .B2(G2105), .ZN(new_n694));
  NAND4_X1  g269(.A1(new_n467), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n695));
  AOI22_X1  g270(.A1(new_n691), .A2(G2105), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AND2_X1   g271(.A1(new_n686), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G29), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G29), .B2(G33), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G21), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G168), .B2(new_n700), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT99), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT100), .B(G1966), .ZN(new_n704));
  OAI221_X1 g279(.A(new_n683), .B1(new_n699), .B2(new_n442), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n680), .A2(G26), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  INV_X1    g282(.A(G128), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n467), .A2(G116), .ZN(new_n709));
  OAI21_X1  g284(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n710));
  OAI22_X1  g285(.A1(new_n485), .A2(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G140), .B2(new_n490), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n707), .B1(new_n712), .B2(new_n680), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G2067), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT31), .B(G11), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT30), .B(G28), .Z(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(G29), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n625), .B2(G29), .ZN(new_n718));
  NOR2_X1   g293(.A1(G171), .A2(new_n700), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G5), .B2(new_n700), .ZN(new_n720));
  INV_X1    g295(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n718), .B1(new_n721), .B2(G1961), .ZN(new_n722));
  AOI211_X1 g297(.A(new_n714), .B(new_n722), .C1(G1961), .C2(new_n721), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n680), .A2(G35), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G162), .B2(new_n680), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT29), .B(G2090), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n703), .B2(new_n704), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n700), .A2(G20), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT23), .Z(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G299), .B2(G16), .ZN(new_n731));
  INV_X1    g306(.A(G1956), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n443), .B2(new_n682), .ZN(new_n734));
  INV_X1    g309(.A(G34), .ZN(new_n735));
  AOI21_X1  g310(.A(G29), .B1(new_n735), .B2(KEYINPUT24), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OAI22_X1  g312(.A1(new_n737), .A2(KEYINPUT98), .B1(KEYINPUT24), .B2(new_n735), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(KEYINPUT98), .B2(new_n737), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G160), .B2(G29), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(G2084), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(G2084), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT26), .Z(new_n744));
  OAI21_X1  g319(.A(G105), .B1(new_n468), .B2(new_n469), .ZN(new_n745));
  INV_X1    g320(.A(G129), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n744), .B(new_n745), .C1(new_n746), .C2(new_n485), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G141), .B2(new_n490), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(new_n680), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n680), .B2(G32), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G1996), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n742), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AOI211_X1 g327(.A(new_n741), .B(new_n752), .C1(new_n750), .C2(new_n751), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n723), .A2(new_n728), .A3(new_n734), .A4(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G16), .A2(G19), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n548), .B2(G16), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT95), .ZN(new_n757));
  AOI211_X1 g332(.A(new_n705), .B(new_n754), .C1(G1341), .C2(new_n757), .ZN(new_n758));
  MUX2_X1   g333(.A(G24), .B(G290), .S(G16), .Z(new_n759));
  AND2_X1   g334(.A1(new_n759), .A2(G1986), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n759), .A2(G1986), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n680), .A2(G25), .ZN(new_n762));
  INV_X1    g337(.A(G119), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n467), .A2(G107), .ZN(new_n764));
  OAI21_X1  g339(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n765));
  OAI22_X1  g340(.A1(new_n485), .A2(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G131), .B2(new_n490), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n762), .B1(new_n767), .B2(new_n680), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT35), .B(G1991), .Z(new_n769));
  XOR2_X1   g344(.A(new_n768), .B(new_n769), .Z(new_n770));
  NOR3_X1   g345(.A1(new_n760), .A2(new_n761), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n700), .A2(G22), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT93), .Z(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G166), .B2(new_n700), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(G1971), .Z(new_n775));
  NOR2_X1   g350(.A1(G16), .A2(G23), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT92), .Z(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G288), .B2(new_n700), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT33), .B(G1976), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n700), .A2(G6), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n579), .B2(new_n700), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT32), .B(G1981), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT91), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n782), .B(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n775), .A2(new_n780), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(KEYINPUT34), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n786), .A2(KEYINPUT34), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n771), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n789), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n700), .A2(G4), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n606), .B2(new_n700), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1348), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n699), .A2(new_n442), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT97), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n757), .A2(G1341), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n796), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND4_X1  g375(.A1(new_n758), .A2(new_n791), .A3(new_n793), .A4(new_n800), .ZN(G150));
  INV_X1    g376(.A(G150), .ZN(G311));
  NOR2_X1   g377(.A1(new_n599), .A2(new_n607), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n512), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(new_n519), .ZN(new_n807));
  INV_X1    g382(.A(G93), .ZN(new_n808));
  INV_X1    g383(.A(G55), .ZN(new_n809));
  OAI22_X1  g384(.A1(new_n514), .A2(new_n808), .B1(new_n809), .B2(new_n517), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n548), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n545), .A2(new_n547), .ZN(new_n813));
  INV_X1    g388(.A(new_n811), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n805), .B(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT39), .ZN(new_n818));
  AOI21_X1  g393(.A(G860), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n818), .B2(new_n817), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n814), .A2(G860), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT37), .Z(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n822), .ZN(G145));
  INV_X1    g398(.A(G130), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT104), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n467), .B2(G118), .ZN(new_n826));
  OR2_X1    g401(.A1(G106), .A2(G2105), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n826), .A2(G2104), .A3(new_n827), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n825), .A2(new_n467), .A3(G118), .ZN(new_n829));
  OAI22_X1  g404(.A1(new_n485), .A2(new_n824), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(G142), .B2(new_n490), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n614), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(new_n767), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT105), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n833), .A2(KEYINPUT105), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n697), .A2(KEYINPUT103), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n496), .A2(new_n505), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n748), .B(new_n712), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  MUX2_X1   g415(.A(new_n834), .B(new_n835), .S(new_n840), .Z(new_n841));
  XNOR2_X1  g416(.A(G162), .B(G160), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT102), .Z(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n625), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(G37), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n841), .A2(new_n844), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XOR2_X1   g424(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n850));
  XNOR2_X1  g425(.A(new_n849), .B(new_n850), .ZN(G395));
  NAND2_X1  g426(.A1(new_n606), .A2(new_n603), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n599), .A2(G299), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT41), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n852), .A2(KEYINPUT41), .A3(new_n853), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n609), .B(new_n816), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(KEYINPUT107), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT107), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n858), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  OAI211_X1 g438(.A(new_n861), .B(new_n863), .C1(new_n859), .C2(new_n854), .ZN(new_n864));
  NAND2_X1  g439(.A1(G290), .A2(new_n579), .ZN(new_n865));
  OAI211_X1 g440(.A(G305), .B(new_n582), .C1(new_n586), .C2(new_n587), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(G303), .B(G288), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n865), .A2(new_n868), .A3(new_n866), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n872), .A2(KEYINPUT42), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT108), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n870), .A2(KEYINPUT108), .A3(new_n871), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n873), .B1(new_n877), .B2(KEYINPUT42), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n864), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n864), .A2(new_n878), .ZN(new_n880));
  OAI21_X1  g455(.A(G868), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(G868), .B2(new_n811), .ZN(G295));
  OAI21_X1  g457(.A(new_n881), .B1(G868), .B2(new_n811), .ZN(G331));
  NAND2_X1  g458(.A1(new_n812), .A2(new_n815), .ZN(new_n884));
  NOR2_X1   g459(.A1(G301), .A2(G286), .ZN(new_n885));
  NOR2_X1   g460(.A1(G168), .A2(G171), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n884), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n886), .B1(new_n567), .B2(G168), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n816), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n856), .A2(new_n890), .A3(new_n857), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT109), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n599), .B(new_n603), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n816), .A2(KEYINPUT109), .A3(new_n888), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n893), .A2(new_n894), .A3(new_n887), .A4(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n877), .A2(new_n891), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n846), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n877), .B1(new_n896), .B2(new_n891), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT43), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(KEYINPUT110), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n893), .A2(new_n887), .A3(new_n895), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n858), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n894), .A2(new_n887), .A3(new_n889), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n877), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n898), .A2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT110), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n909), .B(KEYINPUT43), .C1(new_n898), .C2(new_n899), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n901), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n898), .A2(new_n899), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n898), .A2(new_n905), .A3(new_n907), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT44), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n913), .A2(new_n917), .ZN(G397));
  INV_X1    g493(.A(G1384), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(new_n496), .B2(new_n505), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT45), .B1(new_n920), .B2(KEYINPUT111), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(KEYINPUT111), .B2(new_n920), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n490), .A2(G137), .ZN(new_n923));
  INV_X1    g498(.A(G125), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n482), .B1(new_n689), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(G2105), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n923), .A2(new_n926), .A3(G40), .A4(new_n470), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n922), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n748), .B(G1996), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n712), .B(G2067), .ZN(new_n930));
  AOI211_X1 g505(.A(new_n927), .B(new_n922), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n931), .B(KEYINPUT112), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n932), .A2(new_n769), .A3(new_n767), .ZN(new_n933));
  INV_X1    g508(.A(G2067), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n712), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n928), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G1996), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n928), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT46), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n930), .A2(new_n748), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n928), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(KEYINPUT47), .ZN(new_n943));
  XNOR2_X1  g518(.A(new_n767), .B(new_n769), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n928), .A2(new_n944), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n932), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(G290), .A2(G1986), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n928), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT48), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n936), .A2(new_n943), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT127), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n951), .B(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n927), .A2(new_n920), .ZN(new_n954));
  INV_X1    g529(.A(G8), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(G305), .A2(G1981), .ZN(new_n957));
  INV_X1    g532(.A(G1981), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n579), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT49), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n957), .A2(KEYINPUT49), .A3(new_n959), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(new_n956), .A3(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(G288), .A2(G1976), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(KEYINPUT116), .ZN(new_n966));
  AND2_X1   g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n959), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n956), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n480), .A2(new_n495), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n502), .A2(new_n504), .ZN(new_n974));
  AOI21_X1  g549(.A(G1384), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n927), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n970), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(G2090), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(G1384), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n981), .B1(new_n496), .B2(new_n505), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT113), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n984), .B(new_n981), .C1(new_n496), .C2(new_n505), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n927), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n980), .B1(G164), .B2(G1384), .ZN(new_n987));
  AOI21_X1  g562(.A(G1971), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n989));
  OR3_X1    g564(.A1(new_n979), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(G166), .B2(new_n955), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT115), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n989), .B1(new_n979), .B2(new_n988), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n990), .A2(new_n995), .A3(G8), .A4(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G1976), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n956), .B1(new_n998), .B2(G288), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT52), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT52), .B1(G288), .B2(new_n998), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n956), .B(new_n1001), .C1(new_n998), .C2(G288), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n964), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n969), .B1(new_n997), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n927), .B1(new_n980), .B2(new_n920), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n502), .A2(new_n507), .A3(new_n504), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n507), .B1(new_n502), .B2(new_n504), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n973), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1008), .A2(KEYINPUT45), .A3(new_n919), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n704), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(G2084), .B2(new_n978), .ZN(new_n1012));
  AND3_X1   g587(.A1(new_n1012), .A2(G8), .A3(G168), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT63), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n991), .A2(new_n993), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n990), .A2(new_n996), .A3(G8), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1003), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1017), .A2(new_n997), .A3(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1008), .A2(new_n976), .A3(new_n919), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT117), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G40), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n479), .A2(new_n483), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1024), .B1(new_n975), .B2(new_n976), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1008), .A2(KEYINPUT117), .A3(new_n976), .A4(new_n919), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1022), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1028), .A2(G2090), .ZN(new_n1029));
  OAI21_X1  g604(.A(G8), .B1(new_n1029), .B2(new_n988), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n1015), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n997), .A2(new_n1018), .A3(new_n1031), .A4(new_n1013), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT63), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1004), .B1(new_n1019), .B2(new_n1034), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1011), .B(G168), .C1(G2084), .C2(new_n978), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1036), .A2(new_n1037), .A3(G8), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1012), .A2(G286), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1039), .A2(G8), .A3(new_n1036), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1038), .B1(new_n1040), .B2(KEYINPUT51), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT62), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n997), .A2(new_n1018), .A3(new_n1031), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT126), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n986), .A2(new_n443), .A3(new_n987), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1961), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n978), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n443), .A2(KEYINPUT53), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1048), .B(new_n1050), .C1(new_n1010), .C2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n567), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .A4(new_n1054), .ZN(new_n1055));
  OR2_X1    g630(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1053), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1045), .B1(new_n1058), .B2(new_n1044), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1035), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1052), .A2(new_n567), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n983), .A2(new_n985), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT124), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n467), .B1(new_n925), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(new_n1064), .B2(new_n925), .ZN(new_n1066));
  OR3_X1    g641(.A1(new_n479), .A2(new_n1023), .A3(new_n1051), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n922), .A2(new_n1063), .A3(new_n1066), .A4(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1048), .A2(new_n1050), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1062), .B1(new_n1070), .B2(G171), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1041), .B1(new_n1061), .B2(new_n1071), .ZN(new_n1072));
  OR2_X1    g647(.A1(new_n1070), .A2(new_n567), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n1053), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT125), .B1(new_n1074), .B2(new_n1062), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1074), .A2(KEYINPUT125), .A3(new_n1062), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1072), .B(new_n1044), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1028), .A2(new_n732), .ZN(new_n1078));
  NAND2_X1  g653(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1079));
  OR2_X1    g654(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT56), .B(G2072), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n986), .A2(new_n987), .A3(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .A4(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(G1348), .B1(new_n970), .B2(new_n977), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n954), .A2(new_n934), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT118), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1348), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n976), .B1(new_n1008), .B2(new_n919), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1024), .B1(KEYINPUT50), .B2(new_n920), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(new_n1092), .A3(new_n1085), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1087), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1094), .A2(new_n599), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1078), .A2(new_n1082), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1083), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n606), .B1(new_n1094), .B2(KEYINPUT60), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1094), .A2(KEYINPUT60), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1094), .A2(KEYINPUT60), .A3(new_n606), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1080), .A2(new_n1079), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1025), .B1(new_n1021), .B2(new_n1020), .ZN(new_n1103));
  AOI21_X1  g678(.A(G1956), .B1(new_n1103), .B2(new_n1027), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1082), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1102), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1106), .A2(new_n1083), .ZN(new_n1107));
  AOI22_X1  g682(.A1(new_n1100), .A2(new_n1101), .B1(new_n1107), .B2(KEYINPUT61), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT61), .B1(new_n1096), .B2(KEYINPUT121), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT121), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1106), .A2(new_n1083), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1109), .A2(new_n1111), .A3(KEYINPUT122), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n1106), .A2(new_n1083), .A3(new_n1110), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT61), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1113), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1108), .A2(new_n1112), .A3(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n987), .A2(new_n1063), .A3(new_n937), .A4(new_n1024), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n986), .A2(new_n1121), .A3(new_n987), .A4(new_n937), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n954), .ZN(new_n1124));
  XOR2_X1   g699(.A(KEYINPUT58), .B(G1341), .Z(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT120), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT120), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1126), .ZN(new_n1129));
  AOI211_X1 g704(.A(new_n1128), .B(new_n1129), .C1(new_n1120), .C2(new_n1122), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n548), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT59), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1133), .B(new_n548), .C1(new_n1127), .C2(new_n1130), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1097), .B1(new_n1118), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1077), .B1(new_n1136), .B2(KEYINPUT123), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT123), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1138), .B(new_n1097), .C1(new_n1118), .C2(new_n1135), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1060), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(G290), .A2(G1986), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n928), .B1(new_n1141), .B2(new_n947), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n946), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n953), .B1(new_n1140), .B2(new_n1143), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g719(.A1(G229), .A2(new_n464), .A3(new_n462), .A4(G227), .ZN(new_n1146));
  AND2_X1   g720(.A1(new_n647), .A2(new_n1146), .ZN(new_n1147));
  OR2_X1    g721(.A1(new_n847), .A2(new_n848), .ZN(new_n1148));
  AND3_X1   g722(.A1(new_n911), .A2(new_n1147), .A3(new_n1148), .ZN(G308));
  NAND3_X1  g723(.A1(new_n911), .A2(new_n1147), .A3(new_n1148), .ZN(G225));
endmodule


