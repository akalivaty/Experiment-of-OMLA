//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:17 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n570, new_n571, new_n572, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n583,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n618, new_n619, new_n622, new_n624, new_n625, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT64), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(new_n460), .A2(G137), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n460), .A2(G2104), .ZN(new_n462));
  AOI22_X1  g037(.A1(new_n459), .A2(new_n461), .B1(new_n462), .B2(G101), .ZN(new_n463));
  AOI22_X1  g038(.A1(new_n459), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n463), .B1(new_n464), .B2(new_n460), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G160));
  AND2_X1   g041(.A1(new_n459), .A2(KEYINPUT65), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n459), .A2(KEYINPUT65), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G136), .ZN(new_n471));
  XNOR2_X1  g046(.A(new_n471), .B(KEYINPUT66), .ZN(new_n472));
  OAI21_X1  g047(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(G112), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n473), .B1(new_n474), .B2(G2105), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n469), .A2(new_n460), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NOR3_X1   g052(.A1(new_n472), .A2(new_n475), .A3(new_n477), .ZN(G162));
  OR2_X1    g053(.A1(new_n460), .A2(G114), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n479), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n460), .A2(G114), .ZN(new_n484));
  OAI21_X1  g059(.A(KEYINPUT67), .B1(new_n484), .B2(new_n480), .ZN(new_n485));
  AND2_X1   g060(.A1(G126), .A2(G2105), .ZN(new_n486));
  AOI22_X1  g061(.A1(new_n483), .A2(new_n485), .B1(new_n459), .B2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT68), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT68), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n492), .A2(new_n459), .A3(new_n493), .A4(new_n495), .ZN(new_n496));
  AND2_X1   g071(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n497));
  NOR2_X1   g072(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(KEYINPUT4), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n460), .A2(G138), .ZN(new_n502));
  INV_X1    g077(.A(new_n498), .ZN(new_n503));
  NAND2_X1  g078(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n493), .B1(new_n505), .B2(new_n492), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n487), .B1(new_n501), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  NAND2_X1  g083(.A1(G75), .A2(G543), .ZN(new_n509));
  NAND3_X1  g084(.A1(KEYINPUT70), .A2(KEYINPUT5), .A3(G543), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g086(.A(G543), .B1(KEYINPUT70), .B2(KEYINPUT5), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G62), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n509), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n515), .A2(G651), .B1(new_n520), .B2(G50), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  OAI21_X1  g097(.A(KEYINPUT71), .B1(new_n513), .B2(new_n518), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT70), .A2(KEYINPUT5), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(new_n519), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(new_n510), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n526), .B(new_n527), .C1(new_n517), .C2(new_n516), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n521), .B1(new_n522), .B2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  NAND2_X1  g106(.A1(new_n520), .A2(G51), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(KEYINPUT72), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT7), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n534), .A2(KEYINPUT72), .ZN(new_n537));
  AND3_X1   g112(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n536), .B1(new_n535), .B2(new_n537), .ZN(new_n539));
  OAI211_X1 g114(.A(new_n532), .B(new_n533), .C1(new_n538), .C2(new_n539), .ZN(new_n540));
  AND3_X1   g115(.A1(new_n523), .A2(G89), .A3(new_n528), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n540), .A2(new_n541), .ZN(G168));
  AOI22_X1  g117(.A1(new_n526), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT73), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n544), .A2(new_n545), .A3(G651), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n523), .A2(new_n528), .A3(G90), .ZN(new_n547));
  INV_X1    g122(.A(G651), .ZN(new_n548));
  OAI21_X1  g123(.A(KEYINPUT73), .B1(new_n543), .B2(new_n548), .ZN(new_n549));
  XOR2_X1   g124(.A(KEYINPUT74), .B(G52), .Z(new_n550));
  NAND2_X1  g125(.A1(new_n520), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n546), .A2(new_n547), .A3(new_n549), .A4(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  NAND3_X1  g128(.A1(new_n523), .A2(new_n528), .A3(G81), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n520), .A2(G43), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT76), .ZN(new_n557));
  NAND2_X1  g132(.A1(G68), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G56), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n513), .B2(new_n559), .ZN(new_n560));
  AND3_X1   g135(.A1(new_n560), .A2(KEYINPUT75), .A3(G651), .ZN(new_n561));
  AOI21_X1  g136(.A(KEYINPUT75), .B1(new_n560), .B2(G651), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n554), .A2(new_n564), .A3(new_n555), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n557), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g144(.A(KEYINPUT77), .B(KEYINPUT8), .Z(new_n570));
  NAND2_X1  g145(.A1(G1), .A2(G3), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n570), .B(new_n571), .ZN(new_n572));
  NAND4_X1  g147(.A1(G319), .A2(G483), .A3(G661), .A4(new_n572), .ZN(G188));
  NAND3_X1  g148(.A1(new_n523), .A2(new_n528), .A3(G91), .ZN(new_n574));
  OAI211_X1 g149(.A(G53), .B(G543), .C1(new_n516), .C2(new_n517), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT9), .ZN(new_n576));
  NAND2_X1  g151(.A1(G78), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n513), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(G651), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n574), .A2(new_n576), .A3(new_n580), .ZN(G299));
  INV_X1    g156(.A(G168), .ZN(G286));
  INV_X1    g157(.A(new_n529), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n583), .A2(G87), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n526), .A2(G74), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n585), .A2(G651), .B1(G49), .B2(new_n520), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n584), .A2(new_n586), .ZN(G288));
  NAND2_X1  g162(.A1(new_n583), .A2(G86), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n589), .B(KEYINPUT78), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n513), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n592), .A2(G651), .B1(new_n520), .B2(G48), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n588), .A2(new_n593), .ZN(G305));
  NAND2_X1  g169(.A1(new_n520), .A2(G47), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n596));
  XNOR2_X1  g171(.A(KEYINPUT79), .B(G85), .ZN(new_n597));
  OAI221_X1 g172(.A(new_n595), .B1(new_n548), .B2(new_n596), .C1(new_n529), .C2(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n523), .A2(new_n528), .A3(G92), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n523), .A2(new_n528), .A3(KEYINPUT10), .A4(G92), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g179(.A(KEYINPUT80), .B(G66), .Z(new_n605));
  AOI22_X1  g180(.A1(new_n605), .A2(new_n526), .B1(G79), .B2(G543), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT81), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n548), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n605), .A2(new_n526), .ZN(new_n609));
  AND2_X1   g184(.A1(G79), .A2(G543), .ZN(new_n610));
  OAI21_X1  g185(.A(KEYINPUT81), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n608), .A2(new_n611), .B1(G54), .B2(new_n520), .ZN(new_n612));
  AND2_X1   g187(.A1(new_n604), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n599), .B1(new_n613), .B2(G868), .ZN(G284));
  XOR2_X1   g189(.A(G284), .B(KEYINPUT82), .Z(G321));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  OR3_X1    g191(.A1(G168), .A2(KEYINPUT83), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(KEYINPUT83), .B1(G168), .B2(new_n616), .ZN(new_n618));
  AND3_X1   g193(.A1(new_n574), .A2(new_n580), .A3(new_n576), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n617), .B(new_n618), .C1(G868), .C2(new_n619), .ZN(G297));
  XNOR2_X1  g195(.A(G297), .B(KEYINPUT84), .ZN(G280));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n613), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n613), .A2(new_n622), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(G868), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(G868), .B2(new_n567), .ZN(G323));
  XOR2_X1   g201(.A(KEYINPUT85), .B(KEYINPUT11), .Z(new_n627));
  XNOR2_X1  g202(.A(G323), .B(new_n627), .ZN(G282));
  NAND2_X1  g203(.A1(new_n470), .A2(G135), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n476), .A2(G123), .ZN(new_n630));
  OR2_X1    g205(.A1(G99), .A2(G2105), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n631), .B(G2104), .C1(G111), .C2(new_n460), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(G2096), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(G2096), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n459), .A2(new_n462), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT13), .B(G2100), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n634), .A2(new_n635), .A3(new_n640), .ZN(G156));
  INV_X1    g216(.A(KEYINPUT14), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT15), .B(G2435), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n646), .B1(new_n645), .B2(new_n644), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2451), .B(G2454), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n647), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(G14), .A3(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  INV_X1    g232(.A(KEYINPUT18), .ZN(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(KEYINPUT17), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n658), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(KEYINPUT87), .B(G2100), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(G2072), .B(G2078), .Z(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n661), .B2(KEYINPUT18), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(G2096), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n666), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  XOR2_X1   g248(.A(G1956), .B(G2474), .Z(new_n674));
  XOR2_X1   g249(.A(G1961), .B(G1966), .Z(new_n675));
  AND2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT20), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n674), .A2(new_n675), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  MUX2_X1   g256(.A(new_n681), .B(new_n680), .S(new_n673), .Z(new_n682));
  NOR2_X1   g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G1981), .ZN(new_n684));
  INV_X1    g259(.A(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT88), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n686), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n686), .A2(new_n688), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n686), .A2(new_n688), .ZN(new_n694));
  NAND3_X1  g269(.A1(new_n693), .A2(new_n690), .A3(new_n694), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n692), .A2(new_n695), .ZN(G229));
  INV_X1    g271(.A(G29), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n697), .A2(G32), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n470), .A2(G141), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n476), .A2(G129), .ZN(new_n700));
  NAND3_X1  g275(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT26), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  AOI22_X1  g279(.A1(new_n703), .A2(new_n704), .B1(G105), .B2(new_n462), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n699), .A2(new_n700), .A3(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT96), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n698), .B1(new_n710), .B2(new_n697), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT97), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT27), .B(G1996), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G5), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(G171), .B2(new_n715), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G1961), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT99), .Z(new_n719));
  OR2_X1    g294(.A1(new_n697), .A2(KEYINPUT89), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n697), .A2(KEYINPUT89), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G26), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT28), .Z(new_n725));
  NAND2_X1  g300(.A1(new_n470), .A2(G140), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n476), .A2(G128), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n460), .A2(G116), .ZN(new_n728));
  OAI21_X1  g303(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n726), .B(new_n727), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  OR2_X1    g305(.A1(new_n730), .A2(KEYINPUT95), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(KEYINPUT95), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n725), .B1(new_n733), .B2(G29), .ZN(new_n734));
  INV_X1    g309(.A(G2067), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(G162), .A2(new_n722), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G35), .B2(new_n722), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT101), .B(KEYINPUT29), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G2090), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n736), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n714), .A2(new_n719), .A3(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n739), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n738), .B(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(G1341), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n567), .A2(new_n715), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n715), .B2(G19), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n745), .A2(G2090), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(G168), .A2(new_n715), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n715), .B2(G21), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G164), .A2(new_n723), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G27), .B2(new_n723), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n752), .A2(G1966), .B1(new_n755), .B2(G2078), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G2078), .B2(new_n755), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT24), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n758), .A2(G34), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(G34), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n723), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n465), .B2(new_n697), .ZN(new_n762));
  INV_X1    g337(.A(G2084), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT25), .Z(new_n766));
  AOI22_X1  g341(.A1(new_n459), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n767), .B2(new_n460), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n470), .B2(G139), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(new_n697), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n697), .B2(G33), .ZN(new_n771));
  INV_X1    g346(.A(G2072), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n764), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n772), .B2(new_n771), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n762), .A2(new_n763), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT100), .Z(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n752), .B2(G1966), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n757), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n715), .A2(G4), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n613), .B2(new_n715), .ZN(new_n780));
  INV_X1    g355(.A(G1348), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n748), .A2(new_n746), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT30), .B(G28), .ZN(new_n784));
  OR2_X1    g359(.A1(KEYINPUT31), .A2(G11), .ZN(new_n785));
  NAND2_X1  g360(.A1(KEYINPUT31), .A2(G11), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n784), .A2(new_n697), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n633), .B2(new_n723), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT98), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n715), .A2(G20), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT23), .Z(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G299), .B2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1956), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n717), .B2(G1961), .ZN(new_n794));
  NOR3_X1   g369(.A1(new_n783), .A2(new_n789), .A3(new_n794), .ZN(new_n795));
  NAND4_X1  g370(.A1(new_n749), .A2(new_n778), .A3(new_n782), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n743), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n723), .A2(G25), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT90), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n476), .A2(G119), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT91), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n802));
  INV_X1    g377(.A(G107), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(G2105), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n470), .B2(G131), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n799), .B1(new_n806), .B2(new_n722), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT35), .B(G1991), .Z(new_n808));
  XOR2_X1   g383(.A(new_n807), .B(new_n808), .Z(new_n809));
  INV_X1    g384(.A(KEYINPUT92), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  OR2_X1    g387(.A1(G16), .A2(G24), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G290), .B2(new_n715), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n814), .A2(new_n685), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(new_n685), .ZN(new_n816));
  OR3_X1    g391(.A1(new_n815), .A2(new_n816), .A3(KEYINPUT94), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n811), .A2(new_n812), .A3(new_n817), .ZN(new_n818));
  MUX2_X1   g393(.A(G6), .B(G305), .S(G16), .Z(new_n819));
  XOR2_X1   g394(.A(KEYINPUT32), .B(G1981), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n821), .A2(KEYINPUT93), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(KEYINPUT93), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n715), .A2(G22), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G166), .B2(new_n715), .ZN(new_n825));
  INV_X1    g400(.A(G1971), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n715), .A2(G23), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n584), .A2(new_n586), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n829), .B2(new_n715), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT33), .B(G1976), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n822), .A2(new_n823), .A3(new_n827), .A4(new_n832), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n833), .A2(KEYINPUT34), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(KEYINPUT34), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n818), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT36), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n818), .A2(new_n834), .A3(KEYINPUT36), .A4(new_n835), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n797), .A2(new_n838), .A3(new_n839), .ZN(G311));
  NAND3_X1  g415(.A1(new_n797), .A2(new_n838), .A3(new_n839), .ZN(G150));
  NAND2_X1  g416(.A1(new_n613), .A2(G559), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT38), .ZN(new_n843));
  AOI22_X1  g418(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n844), .A2(new_n548), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n523), .A2(new_n528), .A3(G93), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n520), .A2(G55), .ZN(new_n847));
  AOI21_X1  g422(.A(KEYINPUT102), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n846), .A2(KEYINPUT102), .A3(new_n847), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n845), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n567), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n850), .ZN(new_n853));
  OAI22_X1  g428(.A1(new_n853), .A2(new_n848), .B1(new_n548), .B2(new_n844), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(new_n566), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n843), .B(new_n856), .Z(new_n857));
  OR2_X1    g432(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n858));
  INV_X1    g433(.A(G860), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(KEYINPUT39), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n851), .A2(new_n859), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(KEYINPUT37), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(G145));
  NAND2_X1  g439(.A1(new_n470), .A2(G142), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n476), .A2(G130), .ZN(new_n866));
  OR3_X1    g441(.A1(new_n460), .A2(KEYINPUT103), .A3(G118), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT103), .B1(new_n460), .B2(G118), .ZN(new_n868));
  OR2_X1    g443(.A1(G106), .A2(G2105), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n867), .A2(G2104), .A3(new_n868), .A4(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n865), .A2(new_n866), .A3(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT104), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n872), .A2(new_n638), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n638), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n731), .A2(new_n769), .A3(new_n732), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n769), .B1(new_n731), .B2(new_n732), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n873), .B(new_n874), .C1(new_n876), .C2(new_n877), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n710), .A2(G164), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n708), .A2(new_n709), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n507), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n806), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n882), .A2(new_n806), .A3(new_n884), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n881), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n633), .B(G160), .ZN(new_n891));
  XNOR2_X1  g466(.A(G162), .B(new_n891), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n879), .A2(new_n887), .A3(new_n880), .A4(new_n888), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n890), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n892), .B1(new_n890), .B2(new_n893), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n898), .A2(KEYINPUT40), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT40), .ZN(new_n900));
  NOR3_X1   g475(.A1(new_n896), .A2(new_n900), .A3(new_n897), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n899), .A2(new_n901), .ZN(G395));
  NAND2_X1  g477(.A1(new_n854), .A2(new_n616), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n856), .B(new_n624), .ZN(new_n904));
  AOI21_X1  g479(.A(G299), .B1(new_n604), .B2(new_n612), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n604), .A2(new_n612), .A3(G299), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT41), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT105), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n912), .A2(new_n905), .ZN(new_n913));
  NOR3_X1   g488(.A1(new_n613), .A2(new_n911), .A3(G299), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n910), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n908), .A2(KEYINPUT41), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n909), .B1(new_n904), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(G288), .B(G303), .ZN(new_n919));
  XNOR2_X1  g494(.A(G305), .B(G290), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n919), .B(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT42), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n918), .B(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n903), .B1(new_n923), .B2(new_n616), .ZN(G295));
  OAI21_X1  g499(.A(new_n903), .B1(new_n923), .B2(new_n616), .ZN(G331));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n926));
  XNOR2_X1  g501(.A(G301), .B(G168), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n852), .A2(new_n855), .A3(new_n927), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n928), .A2(new_n908), .ZN(new_n929));
  XOR2_X1   g504(.A(G301), .B(G168), .Z(new_n930));
  NOR2_X1   g505(.A1(new_n567), .A2(new_n851), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n854), .A2(new_n566), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT106), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n856), .A2(new_n935), .A3(new_n930), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n929), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n933), .A2(new_n928), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(new_n916), .A3(new_n915), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n940), .A2(new_n921), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n937), .A2(new_n939), .A3(new_n921), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n895), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT43), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n934), .A2(new_n936), .A3(new_n928), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT41), .B1(new_n913), .B2(new_n914), .ZN(new_n946));
  OR2_X1    g521(.A1(new_n946), .A2(KEYINPUT107), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n908), .A2(new_n910), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n946), .A2(KEYINPUT107), .A3(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n945), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n929), .A2(new_n933), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n921), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n952), .A2(new_n943), .A3(KEYINPUT43), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT108), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n944), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NOR4_X1   g530(.A1(new_n952), .A2(new_n943), .A3(KEYINPUT108), .A4(KEYINPUT43), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n926), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n941), .A2(new_n943), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n952), .A2(new_n943), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT44), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n957), .A2(new_n962), .ZN(G397));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n507), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(G40), .B(new_n463), .C1(new_n464), .C2(new_n460), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n965), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n733), .B(new_n735), .ZN(new_n971));
  INV_X1    g546(.A(G1996), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n883), .B(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n886), .A2(new_n808), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n886), .A2(new_n808), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n971), .A2(new_n973), .A3(new_n974), .A4(new_n975), .ZN(new_n976));
  XNOR2_X1  g551(.A(G290), .B(G1986), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n970), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT118), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT117), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n965), .A2(KEYINPUT50), .ZN(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT68), .B(KEYINPUT4), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT69), .B1(new_n499), .B2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n983), .A2(new_n500), .A3(new_n496), .ZN(new_n984));
  AOI21_X1  g559(.A(G1384), .B1(new_n984), .B2(new_n487), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT50), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g562(.A(KEYINPUT113), .B(G2084), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n981), .A2(new_n967), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n965), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n968), .A2(G1384), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n966), .B1(new_n507), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(G1966), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n989), .B1(new_n994), .B2(KEYINPUT112), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT112), .ZN(new_n996));
  AOI211_X1 g571(.A(new_n996), .B(G1966), .C1(new_n991), .C2(new_n993), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n980), .B(G8), .C1(new_n995), .C2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G8), .ZN(new_n999));
  NOR2_X1   g574(.A1(G168), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n1000), .A2(KEYINPUT51), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1966), .ZN(new_n1003));
  INV_X1    g578(.A(new_n993), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n985), .A2(KEYINPUT45), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n996), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n994), .A2(KEYINPUT112), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(new_n1008), .A3(new_n989), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n980), .B1(new_n1009), .B2(G8), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n979), .B1(new_n1002), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(G8), .B1(new_n995), .B2(new_n997), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT117), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n1013), .A2(KEYINPUT118), .A3(new_n998), .A4(new_n1001), .ZN(new_n1014));
  OAI211_X1 g589(.A(KEYINPUT51), .B(G8), .C1(new_n1009), .C2(G286), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n967), .B1(new_n985), .B2(new_n986), .ZN(new_n1018));
  AOI211_X1 g593(.A(KEYINPUT50), .B(G1384), .C1(new_n984), .C2(new_n487), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI22_X1  g595(.A1(new_n1006), .A2(new_n996), .B1(new_n1020), .B2(new_n988), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n999), .B1(new_n1021), .B2(new_n1008), .ZN(new_n1022));
  OAI211_X1 g597(.A(KEYINPUT116), .B(KEYINPUT51), .C1(new_n1022), .C2(new_n1000), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1011), .A2(new_n1014), .A3(new_n1017), .A4(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT62), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1009), .A2(new_n1000), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1025), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1028));
  OAI21_X1  g603(.A(G8), .B1(new_n965), .B2(new_n966), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1976), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT52), .B1(G288), .B2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1030), .B(new_n1032), .C1(new_n1031), .C2(G288), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1029), .B1(G1976), .B2(new_n829), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(G305), .A2(G1981), .ZN(new_n1037));
  INV_X1    g612(.A(G1981), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n588), .A2(new_n1038), .A3(new_n593), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1037), .A2(KEYINPUT49), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT111), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1040), .B(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(KEYINPUT49), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(new_n1029), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1036), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1020), .A2(new_n741), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n965), .A2(new_n968), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n985), .A2(KEYINPUT45), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(new_n967), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n826), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n999), .B1(new_n1046), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(G303), .A2(G8), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1052), .B(new_n1053), .ZN(new_n1054));
  OR2_X1    g629(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1045), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n1049), .B2(G2078), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1058), .B(KEYINPUT120), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1020), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT119), .B(G1961), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1057), .A2(G2078), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1061), .A2(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(G301), .B1(new_n1060), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1051), .A2(new_n1054), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1056), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1027), .A2(new_n1028), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1070));
  XNOR2_X1  g645(.A(G299), .B(KEYINPUT57), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n966), .B1(new_n965), .B2(KEYINPUT50), .ZN(new_n1072));
  AOI21_X1  g647(.A(G1956), .B1(new_n1072), .B2(new_n987), .ZN(new_n1073));
  INV_X1    g648(.A(new_n968), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n967), .B1(new_n985), .B2(new_n1074), .ZN(new_n1075));
  AOI211_X1 g650(.A(new_n990), .B(G1384), .C1(new_n984), .C2(new_n487), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT56), .B(G2072), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1077), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1075), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1071), .B1(new_n1073), .B2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n619), .B(KEYINPUT57), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1047), .A2(new_n967), .A3(new_n1048), .A4(new_n1077), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1081), .B(new_n1082), .C1(new_n1020), .C2(G1956), .ZN(new_n1083));
  AOI21_X1  g658(.A(KEYINPUT61), .B1(new_n1080), .B2(new_n1083), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1075), .A2(new_n1076), .A3(G1996), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n965), .A2(new_n966), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT58), .B(G1341), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n567), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n1090));
  AND2_X1   g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1084), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1080), .A2(new_n1083), .A3(KEYINPUT61), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT115), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1080), .A2(new_n1083), .A3(new_n1096), .A4(KEYINPUT61), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n781), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT114), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1086), .A2(new_n735), .ZN(new_n1101));
  AND3_X1   g676(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1100), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT60), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  OR2_X1    g679(.A1(new_n1104), .A2(new_n613), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1103), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT60), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1109), .A2(new_n1104), .A3(new_n613), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1093), .A2(new_n1098), .A3(new_n1105), .A4(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1080), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1083), .A2(new_n613), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1111), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1045), .A2(new_n1067), .A3(new_n1055), .ZN(new_n1117));
  XOR2_X1   g692(.A(G301), .B(KEYINPUT54), .Z(new_n1118));
  NOR3_X1   g693(.A1(new_n1076), .A2(new_n1057), .A3(G2078), .ZN(new_n1119));
  XOR2_X1   g694(.A(new_n966), .B(KEYINPUT122), .Z(new_n1120));
  AND3_X1   g695(.A1(new_n1120), .A2(KEYINPUT123), .A3(new_n1047), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT123), .B1(new_n1120), .B2(new_n1047), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1119), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  OAI211_X1 g700(.A(KEYINPUT124), .B(new_n1119), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT121), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1061), .A2(KEYINPUT121), .A3(new_n1062), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1125), .B(new_n1126), .C1(new_n1127), .C2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1118), .B1(new_n1130), .B2(new_n1059), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1118), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1060), .A2(new_n1065), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1117), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1070), .A2(new_n1116), .A3(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1045), .A2(new_n1051), .A3(new_n1054), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1039), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1138));
  NOR2_X1   g713(.A1(G288), .A2(G1976), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1137), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1136), .B1(new_n1140), .B2(new_n1029), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1022), .A2(G168), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1056), .A2(KEYINPUT63), .A3(new_n1067), .A4(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT63), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1145), .B1(new_n1117), .B2(new_n1142), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1141), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1135), .A2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n978), .B1(new_n1069), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n883), .B1(KEYINPUT46), .B2(new_n972), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n971), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(new_n970), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT46), .B1(new_n970), .B2(new_n972), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT125), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1152), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1155), .A2(KEYINPUT126), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1152), .A2(new_n1157), .A3(new_n1154), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1156), .A2(KEYINPUT47), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT47), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n969), .A2(G1986), .A3(G290), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT48), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1162), .B1(new_n976), .B2(new_n970), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n971), .A2(new_n973), .A3(new_n808), .A4(new_n886), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n731), .A2(new_n735), .A3(new_n732), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n969), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  OR2_X1    g741(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1159), .A2(new_n1160), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1149), .A2(new_n1168), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g744(.A1(new_n955), .A2(new_n956), .ZN(new_n1171));
  NAND2_X1  g745(.A1(new_n670), .A2(G319), .ZN(new_n1172));
  XNOR2_X1  g746(.A(new_n1172), .B(KEYINPUT127), .ZN(new_n1173));
  NAND2_X1  g747(.A1(new_n1173), .A2(new_n656), .ZN(new_n1174));
  AOI21_X1  g748(.A(new_n1174), .B1(new_n692), .B2(new_n695), .ZN(new_n1175));
  OAI21_X1  g749(.A(new_n1175), .B1(new_n897), .B2(new_n896), .ZN(new_n1176));
  NOR2_X1   g750(.A1(new_n1171), .A2(new_n1176), .ZN(G308));
  OAI221_X1 g751(.A(new_n1175), .B1(new_n897), .B2(new_n896), .C1(new_n955), .C2(new_n956), .ZN(G225));
endmodule


