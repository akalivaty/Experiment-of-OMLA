//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n439, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n542, new_n543, new_n545, new_n546,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188, new_n1189, new_n1190,
    new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G69), .ZN(new_n439));
  INV_X1    g014(.A(new_n439), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(G452), .ZN(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n439), .A2(G57), .A3(G108), .A4(G120), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT66), .Z(new_n453));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT67), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n470));
  XNOR2_X1  g045(.A(new_n470), .B(KEYINPUT68), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n464), .A2(new_n466), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  NOR3_X1   g048(.A1(new_n472), .A2(new_n473), .A3(G2105), .ZN(new_n474));
  NOR3_X1   g049(.A1(new_n469), .A2(new_n471), .A3(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n472), .A2(KEYINPUT69), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n462), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT70), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n482), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  NAND3_X1  g064(.A1(new_n464), .A2(new_n466), .A3(G126), .ZN(new_n490));
  NAND2_X1  g065(.A1(G114), .A2(G2104), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n463), .A2(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G102), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n462), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n477), .A2(KEYINPUT4), .A3(G138), .A4(new_n462), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n493), .A2(new_n495), .A3(new_n498), .A4(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n503), .B(new_n505), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI21_X1  g088(.A(G543), .B1(new_n510), .B2(new_n511), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n509), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  OAI21_X1  g093(.A(G89), .B1(new_n510), .B2(new_n511), .ZN(new_n519));
  INV_X1    g094(.A(G63), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n520), .B2(new_n508), .ZN(new_n521));
  INV_X1    g096(.A(new_n514), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n521), .A2(new_n506), .B1(new_n522), .B2(G51), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(G286));
  INV_X1    g101(.A(G286), .ZN(G168));
  AOI22_X1  g102(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n508), .ZN(new_n529));
  INV_X1    g104(.A(G90), .ZN(new_n530));
  INV_X1    g105(.A(G52), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n512), .A2(new_n530), .B1(new_n514), .B2(new_n531), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n529), .A2(new_n532), .ZN(G301));
  INV_X1    g108(.A(G301), .ZN(G171));
  AOI22_X1  g109(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n508), .ZN(new_n536));
  INV_X1    g111(.A(G81), .ZN(new_n537));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n512), .A2(new_n537), .B1(new_n514), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  AND3_X1   g116(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G36), .ZN(new_n543));
  XOR2_X1   g118(.A(new_n543), .B(KEYINPUT71), .Z(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n542), .A2(new_n546), .ZN(G188));
  NAND2_X1  g122(.A1(G78), .A2(G543), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n503), .A2(new_n505), .ZN(new_n549));
  INV_X1    g124(.A(G65), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G651), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(KEYINPUT74), .ZN(new_n553));
  INV_X1    g128(.A(new_n512), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G91), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT72), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  OAI211_X1 g132(.A(G53), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n558));
  OAI211_X1 g133(.A(new_n556), .B(new_n557), .C1(new_n558), .C2(KEYINPUT73), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n551), .A2(new_n560), .A3(G651), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n553), .A2(new_n555), .A3(new_n559), .A4(new_n561), .ZN(new_n562));
  OR2_X1    g137(.A1(new_n558), .A2(new_n556), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n556), .B1(new_n558), .B2(KEYINPUT73), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n563), .A2(KEYINPUT9), .A3(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n562), .A2(new_n566), .ZN(G299));
  NAND2_X1  g142(.A1(new_n554), .A2(G87), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n522), .A2(G49), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  NAND3_X1  g146(.A1(new_n503), .A2(new_n505), .A3(G61), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n508), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n554), .A2(G86), .ZN(new_n576));
  OAI211_X1 g151(.A(G48), .B(G543), .C1(new_n510), .C2(new_n511), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G305));
  AOI22_X1  g153(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n508), .ZN(new_n580));
  XOR2_X1   g155(.A(new_n580), .B(KEYINPUT75), .Z(new_n581));
  XOR2_X1   g156(.A(KEYINPUT76), .B(G85), .Z(new_n582));
  NAND2_X1  g157(.A1(new_n554), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n522), .A2(G47), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  INV_X1    g161(.A(G92), .ZN(new_n587));
  OR3_X1    g162(.A1(new_n512), .A2(KEYINPUT10), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(G79), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G66), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n549), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(G651), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n522), .A2(G54), .ZN(new_n593));
  OAI21_X1  g168(.A(KEYINPUT10), .B1(new_n512), .B2(new_n587), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n588), .A2(new_n592), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n595), .A2(KEYINPUT77), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(KEYINPUT77), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n586), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n586), .B1(new_n598), .B2(G868), .ZN(G321));
  NAND2_X1  g175(.A1(G286), .A2(G868), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n562), .A2(new_n566), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G297));
  OAI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n598), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND2_X1  g181(.A1(new_n598), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G868), .B2(new_n540), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g185(.A1(new_n481), .A2(G123), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n483), .A2(G135), .ZN(new_n612));
  NOR2_X1   g187(.A1(G99), .A2(G2105), .ZN(new_n613));
  OAI21_X1  g188(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n611), .B(new_n612), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT79), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(G2096), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n477), .A2(new_n494), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT12), .Z(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT78), .B(KEYINPUT13), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2100), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n619), .B(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n617), .A2(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2430), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2435), .ZN(new_n625));
  XOR2_X1   g200(.A(G2427), .B(G2438), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(KEYINPUT14), .ZN(new_n628));
  XOR2_X1   g203(.A(G2451), .B(G2454), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT16), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n628), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G1341), .B(G1348), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n633), .B(new_n634), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(G14), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(G401));
  XNOR2_X1  g212(.A(G2067), .B(G2678), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT80), .Z(new_n639));
  XOR2_X1   g214(.A(G2072), .B(G2078), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT17), .ZN(new_n641));
  XOR2_X1   g216(.A(G2084), .B(G2090), .Z(new_n642));
  NAND3_X1  g217(.A1(new_n639), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT81), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n639), .A2(new_n640), .ZN(new_n645));
  INV_X1    g220(.A(new_n642), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n645), .B(new_n646), .C1(new_n641), .C2(new_n639), .ZN(new_n647));
  INV_X1    g222(.A(new_n640), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n648), .A2(new_n642), .A3(new_n638), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT18), .Z(new_n650));
  NAND3_X1  g225(.A1(new_n644), .A2(new_n647), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2096), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2100), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G227));
  XNOR2_X1  g229(.A(G1971), .B(G1976), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT19), .ZN(new_n656));
  XOR2_X1   g231(.A(G1956), .B(G2474), .Z(new_n657));
  XOR2_X1   g232(.A(G1961), .B(G1966), .Z(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT20), .Z(new_n661));
  NOR2_X1   g236(.A1(new_n657), .A2(new_n658), .ZN(new_n662));
  INV_X1    g237(.A(new_n659), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n662), .B1(new_n656), .B2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT82), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n656), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n664), .B(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n661), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1991), .B(G1996), .ZN(new_n669));
  INV_X1    g244(.A(G1981), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n668), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT83), .B(G1986), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n674), .B(new_n675), .Z(G229));
  INV_X1    g251(.A(G29), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n615), .A2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G4), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(new_n598), .B2(new_n679), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT85), .ZN(new_n682));
  INV_X1    g257(.A(G1348), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n677), .A2(G27), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G164), .B2(new_n677), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G2078), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(KEYINPUT91), .ZN(new_n688));
  NOR2_X1   g263(.A1(G160), .A2(new_n677), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT24), .B(G34), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n690), .A2(G29), .ZN(new_n691));
  OAI21_X1  g266(.A(G2084), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n679), .A2(G5), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G171), .B2(new_n679), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT90), .Z(new_n695));
  OAI211_X1 g270(.A(new_n688), .B(new_n692), .C1(new_n695), .C2(G1961), .ZN(new_n696));
  NOR2_X1   g271(.A1(G168), .A2(new_n679), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n679), .B2(G21), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT88), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(G1966), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n483), .A2(G141), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n481), .A2(G129), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n494), .A2(G105), .ZN(new_n704));
  NAND3_X1  g279(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT26), .Z(new_n706));
  NAND4_X1  g281(.A1(new_n702), .A2(new_n703), .A3(new_n704), .A4(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G29), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G29), .B2(G32), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT27), .B(G1996), .ZN(new_n711));
  OAI22_X1  g286(.A1(new_n700), .A2(new_n701), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT31), .B(G11), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n698), .B(KEYINPUT88), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(G1966), .ZN(new_n715));
  NOR3_X1   g290(.A1(new_n696), .A2(new_n712), .A3(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(G29), .A2(G35), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G162), .B2(G29), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT29), .B(G2090), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n679), .A2(G19), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n540), .B2(new_n679), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(G1341), .Z(new_n723));
  AND4_X1   g298(.A1(new_n684), .A2(new_n716), .A3(new_n720), .A4(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n679), .A2(G22), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G166), .B2(new_n679), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n726), .A2(G1971), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n726), .A2(G1971), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(KEYINPUT34), .ZN(new_n730));
  NOR2_X1   g305(.A1(G16), .A2(G23), .ZN(new_n731));
  INV_X1    g306(.A(G288), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(G16), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT33), .B(G1976), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n679), .A2(G6), .ZN(new_n736));
  INV_X1    g311(.A(G305), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n736), .B1(new_n737), .B2(new_n679), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT32), .B(G1981), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n729), .A2(new_n730), .A3(new_n735), .A4(new_n740), .ZN(new_n741));
  OR2_X1    g316(.A1(G16), .A2(G24), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G290), .B2(new_n679), .ZN(new_n743));
  INV_X1    g318(.A(G1986), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n727), .A2(new_n728), .A3(new_n735), .ZN(new_n746));
  INV_X1    g321(.A(new_n740), .ZN(new_n747));
  OAI21_X1  g322(.A(KEYINPUT34), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  AND3_X1   g323(.A1(new_n741), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT36), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n743), .A2(new_n744), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n677), .A2(G25), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n481), .A2(G119), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n483), .A2(G131), .ZN(new_n754));
  OR2_X1    g329(.A1(G95), .A2(G2105), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n755), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n756));
  AND3_X1   g331(.A1(new_n753), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n752), .B1(new_n757), .B2(new_n677), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT35), .B(G1991), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT84), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n758), .B(new_n760), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n749), .A2(new_n750), .A3(new_n751), .A4(new_n761), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n741), .A2(new_n751), .A3(new_n748), .A4(new_n745), .ZN(new_n763));
  INV_X1    g338(.A(new_n761), .ZN(new_n764));
  OAI21_X1  g339(.A(KEYINPUT36), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n762), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n679), .A2(KEYINPUT23), .A3(G20), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT23), .ZN(new_n768));
  INV_X1    g343(.A(G20), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(G16), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n767), .B(new_n770), .C1(new_n602), .C2(new_n679), .ZN(new_n771));
  INV_X1    g346(.A(G1956), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n710), .A2(new_n711), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n773), .B(new_n774), .C1(KEYINPUT91), .C2(new_n687), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n695), .A2(G1961), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n481), .A2(G128), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n483), .A2(G140), .ZN(new_n778));
  OR2_X1    g353(.A1(G104), .A2(G2105), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n779), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n777), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G29), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n677), .A2(G26), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(G2067), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT30), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n677), .B1(new_n789), .B2(G28), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT89), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n789), .A2(G28), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n790), .A2(new_n791), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n788), .A2(new_n795), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n775), .A2(new_n776), .A3(new_n796), .ZN(new_n797));
  AND4_X1   g372(.A1(new_n678), .A2(new_n724), .A3(new_n766), .A4(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(G29), .A2(G33), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n483), .A2(G139), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT87), .B(KEYINPUT25), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n494), .A2(G103), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n800), .B(new_n803), .C1(new_n462), .C2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n799), .B1(new_n805), .B2(new_n677), .ZN(new_n806));
  XOR2_X1   g381(.A(new_n806), .B(G2072), .Z(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  OR3_X1    g383(.A1(new_n689), .A2(G2084), .A3(new_n691), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n798), .A2(KEYINPUT92), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT92), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n716), .A2(new_n684), .A3(new_n720), .A4(new_n723), .ZN(new_n812));
  INV_X1    g387(.A(new_n797), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n814), .A2(new_n809), .A3(new_n678), .A4(new_n766), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n811), .B1(new_n815), .B2(new_n807), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n810), .A2(new_n816), .ZN(G311));
  NAND4_X1  g392(.A1(new_n798), .A2(KEYINPUT93), .A3(new_n808), .A4(new_n809), .ZN(new_n818));
  INV_X1    g393(.A(KEYINPUT93), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n815), .B2(new_n807), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n818), .A2(new_n820), .ZN(G150));
  AOI22_X1  g396(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n822), .A2(new_n508), .ZN(new_n823));
  INV_X1    g398(.A(G93), .ZN(new_n824));
  INV_X1    g399(.A(G55), .ZN(new_n825));
  OAI22_X1  g400(.A1(new_n512), .A2(new_n824), .B1(new_n514), .B2(new_n825), .ZN(new_n826));
  OR3_X1    g401(.A1(new_n823), .A2(KEYINPUT94), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(KEYINPUT94), .B1(new_n823), .B2(new_n826), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n829), .A2(G860), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT37), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n598), .A2(G559), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n540), .B1(new_n827), .B2(new_n828), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n823), .A2(new_n826), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n836), .A2(new_n536), .A3(new_n539), .ZN(new_n837));
  OR3_X1    g412(.A1(new_n835), .A2(KEYINPUT95), .A3(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(KEYINPUT95), .B1(new_n835), .B2(new_n837), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n834), .B(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n831), .B1(new_n841), .B2(G860), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT96), .Z(G145));
  XNOR2_X1  g418(.A(new_n488), .B(G160), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(new_n615), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n781), .B(G164), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(new_n707), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(new_n805), .Z(new_n848));
  INV_X1    g423(.A(new_n619), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n483), .A2(G142), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(KEYINPUT97), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n481), .A2(G130), .ZN(new_n852));
  OR2_X1    g427(.A1(G106), .A2(G2105), .ZN(new_n853));
  OAI211_X1 g428(.A(new_n853), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT97), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n483), .A2(new_n855), .A3(G142), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n851), .A2(new_n852), .A3(new_n854), .A4(new_n856), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n857), .A2(new_n757), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(new_n757), .ZN(new_n859));
  OAI21_X1  g434(.A(KEYINPUT98), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NOR3_X1   g436(.A1(new_n858), .A2(new_n859), .A3(KEYINPUT98), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n849), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n858), .A2(new_n859), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT98), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n866), .A2(new_n619), .A3(new_n860), .ZN(new_n867));
  AOI21_X1  g442(.A(KEYINPUT99), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n863), .A2(KEYINPUT99), .A3(new_n867), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n848), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n870), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n847), .B(new_n805), .ZN(new_n873));
  NOR3_X1   g448(.A1(new_n872), .A2(new_n868), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n845), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n873), .B1(new_n872), .B2(new_n868), .ZN(new_n876));
  INV_X1    g451(.A(new_n845), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n863), .A2(new_n867), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n876), .B(new_n877), .C1(new_n878), .C2(new_n873), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n875), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT40), .ZN(G395));
  AOI21_X1  g457(.A(new_n840), .B1(new_n605), .B2(new_n598), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n607), .B1(new_n838), .B2(new_n839), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n886));
  INV_X1    g461(.A(new_n595), .ZN(new_n887));
  NAND3_X1  g462(.A1(G299), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(G299), .A2(new_n887), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n602), .A2(new_n595), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n888), .B1(new_n891), .B2(new_n886), .ZN(new_n892));
  XOR2_X1   g467(.A(KEYINPUT101), .B(KEYINPUT41), .Z(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  AOI22_X1  g469(.A1(new_n892), .A2(new_n893), .B1(new_n894), .B2(new_n891), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n885), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n892), .B1(new_n883), .B2(new_n884), .ZN(new_n897));
  AND2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g473(.A(G303), .B(new_n732), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n737), .ZN(new_n900));
  XNOR2_X1  g475(.A(G303), .B(G288), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(G305), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n903), .A2(G290), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(G290), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(KEYINPUT42), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n898), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n898), .A2(new_n907), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n898), .A2(KEYINPUT102), .A3(new_n907), .ZN(new_n912));
  AND4_X1   g487(.A1(G868), .A2(new_n910), .A3(new_n911), .A4(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n829), .A2(G868), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(G295));
  NOR2_X1   g490(.A1(new_n913), .A2(new_n914), .ZN(G331));
  NAND3_X1  g491(.A1(new_n889), .A2(KEYINPUT41), .A3(new_n890), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT103), .ZN(new_n918));
  XNOR2_X1  g493(.A(G301), .B(G286), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n838), .A2(new_n839), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n919), .ZN(new_n921));
  INV_X1    g496(.A(new_n839), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n835), .A2(KEYINPUT95), .A3(new_n837), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n918), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n920), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n892), .B1(new_n926), .B2(new_n893), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n906), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n895), .A2(new_n926), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n924), .A2(new_n892), .A3(new_n920), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(new_n906), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n928), .A2(new_n933), .A3(new_n880), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n928), .A2(new_n933), .A3(KEYINPUT105), .A4(new_n880), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(KEYINPUT43), .A3(new_n937), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n929), .A2(new_n906), .A3(new_n930), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n906), .B1(new_n929), .B2(new_n930), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n939), .A2(new_n940), .A3(G37), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n938), .A2(KEYINPUT44), .A3(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n928), .A2(new_n933), .A3(new_n942), .A4(new_n880), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(new_n941), .B2(new_n942), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n946), .A2(KEYINPUT104), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT104), .B1(new_n946), .B2(new_n947), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n944), .B1(new_n948), .B2(new_n949), .ZN(G397));
  OR2_X1    g525(.A1(G290), .A2(G1986), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n952));
  NAND2_X1  g527(.A1(G290), .A2(G1986), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G1384), .ZN(new_n955));
  INV_X1    g530(.A(new_n491), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n956), .B1(new_n477), .B2(G126), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n495), .B1(new_n957), .B2(new_n462), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n498), .A2(new_n499), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  XOR2_X1   g535(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n467), .A2(new_n468), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n464), .A2(new_n466), .A3(new_n462), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n964), .A2(G2105), .B1(new_n965), .B2(G137), .ZN(new_n966));
  INV_X1    g541(.A(new_n471), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(G40), .A3(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n963), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(G290), .A2(KEYINPUT107), .A3(G1986), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n954), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G1996), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n707), .B(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n781), .B(new_n787), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n757), .B(new_n760), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n969), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n971), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n575), .A2(new_n576), .A3(new_n670), .A4(new_n577), .ZN(new_n979));
  INV_X1    g554(.A(G86), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n577), .B1(new_n512), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(G1981), .B1(new_n981), .B2(new_n574), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT49), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT49), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n979), .A2(new_n982), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n988));
  XOR2_X1   g563(.A(KEYINPUT110), .B(G8), .Z(new_n989));
  OAI211_X1 g564(.A(new_n988), .B(new_n989), .C1(new_n960), .C2(new_n968), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NAND4_X1  g566(.A1(G160), .A2(new_n500), .A3(G40), .A4(new_n955), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n988), .B1(new_n992), .B2(new_n989), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n987), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1976), .ZN(new_n995));
  NOR2_X1   g570(.A1(G288), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n989), .B1(new_n960), .B2(new_n968), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT111), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n996), .B1(new_n998), .B2(new_n990), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n994), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1000), .B1(new_n732), .B2(G1976), .ZN(new_n1002));
  AOI211_X1 g577(.A(new_n996), .B(new_n1002), .C1(new_n998), .C2(new_n990), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1971), .ZN(new_n1006));
  INV_X1    g581(.A(G40), .ZN(new_n1007));
  NOR4_X1   g582(.A1(new_n469), .A2(new_n471), .A3(new_n474), .A4(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT45), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1008), .B1(new_n960), .B2(new_n1009), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n498), .A2(new_n499), .ZN(new_n1011));
  AOI22_X1  g586(.A1(new_n492), .A2(G2105), .B1(G102), .B2(new_n494), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1384), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1013), .A2(new_n961), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1006), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT108), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n968), .B1(new_n1013), .B2(KEYINPUT45), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n963), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT108), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1018), .A2(new_n1019), .A3(new_n1006), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT50), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n960), .A2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n500), .A2(KEYINPUT50), .A3(new_n955), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n968), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G2090), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1016), .A2(new_n1020), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(G303), .A2(G8), .ZN(new_n1028));
  XNOR2_X1  g603(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1028), .B(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1027), .A2(G8), .A3(new_n1031), .ZN(new_n1032));
  XOR2_X1   g607(.A(new_n979), .B(KEYINPUT112), .Z(new_n1033));
  AND2_X1   g608(.A1(new_n994), .A2(new_n995), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1033), .B1(new_n1034), .B2(new_n732), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n991), .A2(new_n993), .ZN(new_n1036));
  OAI22_X1  g611(.A1(new_n1005), .A2(new_n1032), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1971), .B1(new_n1017), .B2(new_n963), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT113), .ZN(new_n1039));
  AOI21_X1  g614(.A(G2090), .B1(new_n1024), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1023), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT50), .B1(new_n500), .B2(new_n955), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1008), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT113), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1038), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n989), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1030), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n955), .B(new_n961), .C1(new_n958), .C2(new_n959), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n500), .A2(KEYINPUT115), .A3(new_n955), .A4(new_n961), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1053), .B(new_n1008), .C1(new_n1013), .C2(KEYINPUT45), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n966), .A2(KEYINPUT45), .A3(G40), .A4(new_n967), .ZN(new_n1055));
  OAI211_X1 g630(.A(KEYINPUT114), .B(new_n1055), .C1(new_n960), .C2(new_n968), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1052), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G2084), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1057), .A2(new_n701), .B1(new_n1058), .B2(new_n1024), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n1059), .A2(G286), .A3(new_n1046), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1047), .A2(new_n1004), .A3(new_n1060), .A4(new_n1032), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT63), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1061), .A2(KEYINPUT116), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT116), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1004), .A2(new_n1032), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1027), .A2(G8), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1062), .B1(new_n1067), .B2(new_n1030), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1066), .A2(new_n1060), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1037), .B1(new_n1065), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n1071));
  INV_X1    g646(.A(G2078), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1017), .A2(new_n1072), .A3(new_n963), .ZN(new_n1073));
  INV_X1    g648(.A(G1961), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1071), .A2(new_n1073), .B1(new_n1043), .B2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1052), .A2(new_n1072), .A3(new_n1054), .A4(new_n1056), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1076), .A2(KEYINPUT122), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT53), .B1(new_n1076), .B2(KEYINPUT122), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1075), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT123), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1079), .A2(new_n1080), .A3(G171), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1080), .B1(new_n1079), .B2(G171), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1075), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(G171), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1081), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT124), .B1(new_n1085), .B2(KEYINPUT54), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT124), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT54), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1079), .A2(G171), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(KEYINPUT123), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1079), .A2(new_n1080), .A3(G171), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1087), .B(new_n1088), .C1(new_n1092), .C2(new_n1084), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1086), .A2(new_n1093), .ZN(new_n1094));
  XOR2_X1   g669(.A(KEYINPUT56), .B(G2072), .Z(new_n1095));
  OAI22_X1  g670(.A1(new_n1018), .A2(new_n1095), .B1(new_n1024), .B2(G1956), .ZN(new_n1096));
  OR2_X1    g671(.A1(new_n1096), .A2(KEYINPUT119), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n602), .A2(KEYINPUT117), .A3(new_n1098), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1098), .A2(KEYINPUT117), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(KEYINPUT117), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1100), .B(new_n1101), .C1(new_n562), .C2(new_n566), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1096), .A2(KEYINPUT119), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1097), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n598), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n992), .B(KEYINPUT118), .ZN(new_n1107));
  OAI22_X1  g682(.A1(new_n1107), .A2(G2067), .B1(G1348), .B2(new_n1024), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1105), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1096), .A2(new_n1103), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(new_n1096), .B2(new_n1103), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1112), .B1(new_n1115), .B2(KEYINPUT61), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT61), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n1096), .A2(new_n1114), .A3(new_n1103), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1117), .B1(new_n1118), .B2(new_n1111), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT60), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1108), .A2(new_n1120), .ZN(new_n1121));
  OAI221_X1 g696(.A(KEYINPUT60), .B1(G1348), .B2(new_n1024), .C1(new_n1107), .C2(G2067), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(new_n598), .A3(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1109), .A2(KEYINPUT60), .A3(new_n1106), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1116), .A2(new_n1119), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT58), .B(G1341), .Z(new_n1126));
  AND2_X1   g701(.A1(new_n1107), .A2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1018), .A2(G1996), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n540), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n1129), .B(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1113), .B1(new_n1125), .B2(new_n1131), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1066), .A2(new_n1047), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1083), .A2(G171), .ZN(new_n1134));
  OAI211_X1 g709(.A(new_n1134), .B(KEYINPUT54), .C1(new_n1079), .C2(G171), .ZN(new_n1135));
  NOR2_X1   g710(.A1(G168), .A2(new_n1046), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1059), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1057), .A2(new_n701), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1024), .A2(new_n1058), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1046), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT121), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT51), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(new_n1059), .B2(new_n1046), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1142), .A2(new_n1143), .A3(new_n1145), .A4(new_n1137), .ZN(new_n1146));
  INV_X1    g721(.A(G8), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1137), .B1(new_n1059), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT51), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1138), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1132), .A2(new_n1133), .A3(new_n1135), .A4(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1070), .B1(new_n1094), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1138), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n1092), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1133), .B1(new_n1150), .B2(new_n1156), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1154), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AOI22_X1  g736(.A1(new_n1150), .A2(new_n1156), .B1(new_n1091), .B2(new_n1090), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n989), .ZN(new_n1164));
  AOI21_X1  g739(.A(KEYINPUT51), .B1(new_n1164), .B2(new_n1144), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1136), .B1(new_n1141), .B2(KEYINPUT121), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n1165), .A2(new_n1166), .B1(KEYINPUT51), .B2(new_n1148), .ZN(new_n1167));
  OAI21_X1  g742(.A(KEYINPUT62), .B1(new_n1167), .B2(new_n1138), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1162), .A2(KEYINPUT125), .A3(new_n1133), .A4(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1161), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n978), .B1(new_n1153), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n969), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n973), .A2(new_n974), .A3(new_n760), .A4(new_n757), .ZN(new_n1173));
  OR2_X1    g748(.A1(new_n781), .A2(G2067), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1172), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1172), .B1(new_n974), .B2(new_n708), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT127), .ZN(new_n1177));
  XNOR2_X1  g752(.A(KEYINPUT126), .B(KEYINPUT46), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1178), .B1(new_n1172), .B2(G1996), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n969), .B(new_n972), .C1(KEYINPUT126), .C2(KEYINPUT46), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1177), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1181), .B(KEYINPUT47), .Z(new_n1182));
  NOR2_X1   g757(.A1(new_n951), .A2(new_n1172), .ZN(new_n1183));
  XOR2_X1   g758(.A(new_n1183), .B(KEYINPUT48), .Z(new_n1184));
  AOI211_X1 g759(.A(new_n1175), .B(new_n1182), .C1(new_n977), .C2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1171), .A2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g761(.A1(new_n881), .A2(G319), .ZN(new_n1188));
  INV_X1    g762(.A(G229), .ZN(new_n1189));
  NAND4_X1  g763(.A1(new_n946), .A2(new_n636), .A3(new_n653), .A4(new_n1189), .ZN(new_n1190));
  NOR2_X1   g764(.A1(new_n1188), .A2(new_n1190), .ZN(G308));
  AND3_X1   g765(.A1(new_n946), .A2(new_n636), .A3(new_n1189), .ZN(new_n1192));
  NAND4_X1  g766(.A1(new_n1192), .A2(G319), .A3(new_n653), .A4(new_n881), .ZN(G225));
endmodule


