//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n536, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n549, new_n551, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n567, new_n568,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1164, new_n1165;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT65), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n453), .A2(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT69), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  AND2_X1   g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(G2105), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n470), .A2(G137), .B1(G101), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n475), .B1(new_n468), .B2(new_n469), .ZN(new_n476));
  MUX2_X1   g051(.A(G100), .B(G112), .S(G2105), .Z(new_n477));
  AOI22_X1  g052(.A1(G124), .A2(new_n476), .B1(new_n477), .B2(G2104), .ZN(new_n478));
  INV_X1    g053(.A(G136), .ZN(new_n479));
  INV_X1    g054(.A(new_n470), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT70), .Z(G162));
  AND2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  OAI211_X1 g059(.A(G138), .B(new_n475), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n485), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(G114), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G102), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(G2105), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n476), .A2(G126), .B1(G2104), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT4), .B1(new_n485), .B2(new_n486), .ZN(new_n493));
  AOI21_X1  g068(.A(KEYINPUT71), .B1(new_n470), .B2(G138), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n488), .B(new_n492), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  INV_X1    g071(.A(G88), .ZN(new_n497));
  AOI21_X1  g072(.A(KEYINPUT72), .B1(KEYINPUT73), .B2(G651), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT6), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n500), .B1(new_n503), .B2(new_n498), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT74), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n505), .A2(KEYINPUT75), .A3(KEYINPUT5), .A4(G543), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n507), .B1(KEYINPUT74), .B2(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT75), .A2(G543), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n504), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n504), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n497), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n511), .A2(G62), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT76), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n517), .B(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(KEYINPUT77), .A3(G651), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT77), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n519), .B1(new_n511), .B2(G62), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n524), .B2(new_n502), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n515), .B1(new_n522), .B2(new_n525), .ZN(G166));
  INV_X1    g101(.A(new_n512), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G89), .ZN(new_n528));
  INV_X1    g103(.A(new_n513), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G51), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND4_X1  g108(.A1(new_n528), .A2(new_n530), .A3(new_n531), .A4(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  AOI22_X1  g110(.A1(new_n511), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(new_n502), .ZN(new_n537));
  XOR2_X1   g112(.A(KEYINPUT78), .B(G90), .Z(new_n538));
  NAND2_X1  g113(.A1(new_n527), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n529), .A2(G52), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n537), .A2(new_n539), .A3(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  AOI22_X1  g117(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n502), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT79), .ZN(new_n545));
  AOI22_X1  g120(.A1(G81), .A2(new_n527), .B1(new_n529), .B2(G43), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  XOR2_X1   g125(.A(KEYINPUT80), .B(KEYINPUT8), .Z(new_n551));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n549), .A2(new_n553), .ZN(G188));
  INV_X1    g129(.A(G53), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT81), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n555), .B1(new_n556), .B2(KEYINPUT9), .ZN(new_n557));
  OAI211_X1 g132(.A(new_n529), .B(new_n557), .C1(new_n556), .C2(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n527), .A2(G91), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n511), .A2(G65), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT82), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  OAI211_X1 g139(.A(KEYINPUT81), .B(new_n564), .C1(new_n513), .C2(new_n555), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n558), .A2(new_n559), .A3(new_n563), .A4(new_n565), .ZN(G299));
  NAND2_X1  g141(.A1(new_n522), .A2(new_n525), .ZN(new_n567));
  INV_X1    g142(.A(new_n515), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(G303));
  OAI21_X1  g144(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n570));
  INV_X1    g145(.A(G49), .ZN(new_n571));
  INV_X1    g146(.A(G87), .ZN(new_n572));
  OAI221_X1 g147(.A(new_n570), .B1(new_n513), .B2(new_n571), .C1(new_n572), .C2(new_n512), .ZN(G288));
  AOI22_X1  g148(.A1(new_n511), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n574));
  OR2_X1    g149(.A1(new_n574), .A2(new_n502), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n527), .A2(G86), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n529), .A2(G48), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n575), .A2(new_n576), .A3(KEYINPUT83), .A4(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT83), .ZN(new_n579));
  INV_X1    g154(.A(G86), .ZN(new_n580));
  INV_X1    g155(.A(G48), .ZN(new_n581));
  OAI22_X1  g156(.A1(new_n580), .A2(new_n512), .B1(new_n513), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n574), .A2(new_n502), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n579), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n578), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G305));
  NAND2_X1  g161(.A1(new_n529), .A2(G47), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  XOR2_X1   g163(.A(KEYINPUT84), .B(G85), .Z(new_n589));
  OAI221_X1 g164(.A(new_n587), .B1(new_n502), .B2(new_n588), .C1(new_n512), .C2(new_n589), .ZN(G290));
  INV_X1    g165(.A(G868), .ZN(new_n591));
  NOR2_X1   g166(.A1(G301), .A2(new_n591), .ZN(new_n592));
  AND3_X1   g167(.A1(new_n504), .A2(new_n511), .A3(G92), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n593), .B(KEYINPUT10), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  XOR2_X1   g170(.A(new_n595), .B(KEYINPUT85), .Z(new_n596));
  INV_X1    g171(.A(new_n511), .ZN(new_n597));
  XNOR2_X1  g172(.A(KEYINPUT86), .B(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(new_n529), .B2(G54), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n592), .B1(new_n602), .B2(new_n591), .ZN(G284));
  AOI21_X1  g178(.A(new_n592), .B1(new_n602), .B2(new_n591), .ZN(G321));
  MUX2_X1   g179(.A(G286), .B(G299), .S(new_n591), .Z(G297));
  MUX2_X1   g180(.A(G286), .B(G299), .S(new_n591), .Z(G280));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n602), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n547), .A2(new_n591), .ZN(new_n609));
  NOR2_X1   g184(.A1(new_n601), .A2(G559), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT11), .Z(G282));
  INV_X1    g188(.A(new_n612), .ZN(G323));
  NAND2_X1  g189(.A1(new_n470), .A2(G2104), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XOR2_X1   g191(.A(KEYINPUT87), .B(KEYINPUT13), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT88), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G2100), .ZN(new_n620));
  INV_X1    g195(.A(G2100), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(KEYINPUT88), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n618), .A2(new_n619), .A3(G2100), .ZN(new_n623));
  MUX2_X1   g198(.A(G99), .B(G111), .S(G2105), .Z(new_n624));
  AOI22_X1  g199(.A1(G123), .A2(new_n476), .B1(new_n624), .B2(G2104), .ZN(new_n625));
  INV_X1    g200(.A(G135), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(new_n480), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  NAND3_X1  g203(.A1(new_n622), .A2(new_n623), .A3(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT16), .ZN(new_n631));
  XOR2_X1   g206(.A(G2443), .B(G2446), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G1341), .B(G1348), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT89), .B(KEYINPUT14), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT15), .B(G2435), .Z(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT90), .B(G2438), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2430), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n636), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n639), .B2(new_n640), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n635), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n635), .A2(new_n642), .ZN(new_n644));
  AND3_X1   g219(.A1(new_n643), .A2(G14), .A3(new_n644), .ZN(G401));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  XNOR2_X1  g221(.A(G2072), .B(G2078), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT18), .Z(new_n650));
  INV_X1    g225(.A(new_n646), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n647), .A2(KEYINPUT17), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(new_n648), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n651), .B2(new_n652), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n646), .A2(new_n648), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n647), .B1(new_n656), .B2(KEYINPUT17), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n650), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT91), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2096), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2100), .ZN(G227));
  XOR2_X1   g236(.A(G1956), .B(G2474), .Z(new_n662));
  XOR2_X1   g237(.A(G1961), .B(G1966), .Z(new_n663));
  AND2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT92), .Z(new_n665));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT20), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n662), .A2(new_n663), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n667), .A2(new_n664), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n667), .B2(new_n670), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n675), .B(new_n678), .ZN(G229));
  NAND2_X1  g254(.A1(G166), .A2(G16), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(G16), .B2(G22), .ZN(new_n681));
  INV_X1    g256(.A(G1971), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(G16), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G23), .ZN(new_n685));
  INV_X1    g260(.A(G288), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n685), .B1(new_n686), .B2(new_n684), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT33), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n681), .A2(new_n682), .ZN(new_n690));
  AND3_X1   g265(.A1(new_n683), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(G6), .A2(G16), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n693), .B1(G305), .B2(new_n684), .ZN(new_n694));
  XOR2_X1   g269(.A(KEYINPUT32), .B(G1981), .Z(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n694), .B(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n691), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(KEYINPUT34), .ZN(new_n699));
  INV_X1    g274(.A(KEYINPUT34), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n691), .A2(new_n697), .A3(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(G95), .B(G107), .S(G2105), .Z(new_n702));
  AOI22_X1  g277(.A1(G119), .A2(new_n476), .B1(new_n702), .B2(G2104), .ZN(new_n703));
  INV_X1    g278(.A(G131), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(new_n480), .ZN(new_n705));
  MUX2_X1   g280(.A(G25), .B(new_n705), .S(G29), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT93), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT35), .B(G1991), .Z(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n707), .B(new_n709), .ZN(new_n710));
  OR2_X1    g285(.A1(G16), .A2(G24), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G290), .B2(new_n684), .ZN(new_n712));
  INV_X1    g287(.A(G1986), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n712), .A2(new_n713), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT94), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT36), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR4_X1   g293(.A1(new_n710), .A2(new_n714), .A3(new_n715), .A4(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n699), .A2(new_n701), .A3(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(G16), .A2(G19), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n547), .B2(G16), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(KEYINPUT95), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(KEYINPUT95), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1341), .ZN(new_n728));
  INV_X1    g303(.A(G29), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G26), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT28), .Z(new_n731));
  MUX2_X1   g306(.A(G104), .B(G116), .S(G2105), .Z(new_n732));
  AOI22_X1  g307(.A1(G128), .A2(new_n476), .B1(new_n732), .B2(G2104), .ZN(new_n733));
  INV_X1    g308(.A(G140), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(new_n480), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT96), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n731), .B1(new_n737), .B2(G29), .ZN(new_n738));
  INV_X1    g313(.A(G2067), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(G1348), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n602), .A2(G16), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G4), .B2(G16), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n740), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(new_n741), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OR2_X1    g321(.A1(G162), .A2(new_n729), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n729), .A2(G35), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT29), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n749), .A2(new_n750), .ZN(new_n753));
  OAI21_X1  g328(.A(G2090), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n753), .ZN(new_n755));
  INV_X1    g330(.A(G2090), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n755), .A2(new_n756), .A3(new_n751), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n746), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n729), .A2(G32), .ZN(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT26), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G105), .B2(new_n471), .ZN(new_n762));
  INV_X1    g337(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n476), .A2(G129), .ZN(new_n764));
  INV_X1    g339(.A(G141), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n765), .B2(new_n480), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n759), .B1(new_n767), .B2(G29), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT27), .B(G1996), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  AND2_X1   g345(.A1(KEYINPUT24), .A2(G34), .ZN(new_n771));
  NOR2_X1   g346(.A1(KEYINPUT24), .A2(G34), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n729), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n473), .B2(new_n729), .ZN(new_n774));
  INV_X1    g349(.A(G2084), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n770), .A2(new_n776), .ZN(new_n777));
  XOR2_X1   g352(.A(KEYINPUT97), .B(KEYINPUT25), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n471), .A2(G103), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  AND2_X1   g355(.A1(new_n462), .A2(G127), .ZN(new_n781));
  AND2_X1   g356(.A1(G115), .A2(G2104), .ZN(new_n782));
  OAI21_X1  g357(.A(G2105), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n470), .A2(G139), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n780), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  MUX2_X1   g360(.A(G33), .B(new_n785), .S(G29), .Z(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(G2072), .Z(new_n787));
  XOR2_X1   g362(.A(KEYINPUT31), .B(G11), .Z(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT30), .B(G28), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n788), .B1(new_n729), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n627), .B2(new_n729), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(new_n774), .B2(new_n775), .ZN(new_n792));
  NOR2_X1   g367(.A1(G27), .A2(G29), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G164), .B2(G29), .ZN(new_n794));
  INV_X1    g369(.A(G2078), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n777), .A2(new_n787), .A3(new_n792), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n684), .A2(G20), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(KEYINPUT23), .Z(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(G299), .B2(G16), .ZN(new_n800));
  INV_X1    g375(.A(G1956), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n684), .A2(G21), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G168), .B2(new_n684), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1966), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n684), .A2(G5), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G171), .B2(new_n684), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1961), .ZN(new_n808));
  NOR4_X1   g383(.A1(new_n797), .A2(new_n802), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  AND3_X1   g384(.A1(new_n728), .A2(new_n758), .A3(new_n809), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n722), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n720), .A2(new_n721), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(G311));
  INV_X1    g388(.A(KEYINPUT98), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n811), .B2(new_n812), .ZN(new_n815));
  AND4_X1   g390(.A1(new_n814), .A2(new_n722), .A3(new_n810), .A4(new_n812), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(G150));
  NAND2_X1  g392(.A1(G80), .A2(G543), .ZN(new_n818));
  INV_X1    g393(.A(G67), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n818), .B1(new_n597), .B2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT99), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n502), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n821), .B2(new_n820), .ZN(new_n823));
  AOI22_X1  g398(.A1(G93), .A2(new_n527), .B1(new_n529), .B2(G55), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G860), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT37), .Z(new_n827));
  NAND4_X1  g402(.A1(new_n545), .A2(new_n823), .A3(new_n546), .A4(new_n824), .ZN(new_n828));
  INV_X1    g403(.A(new_n828), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n545), .A2(new_n546), .B1(new_n823), .B2(new_n824), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT38), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n602), .A2(G559), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT100), .Z(new_n836));
  INV_X1    g411(.A(G860), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n834), .B2(KEYINPUT39), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n827), .B1(new_n836), .B2(new_n838), .ZN(G145));
  XNOR2_X1  g414(.A(new_n737), .B(G164), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n767), .B(new_n785), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n616), .B(new_n705), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n476), .A2(G130), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT101), .ZN(new_n845));
  MUX2_X1   g420(.A(G106), .B(G118), .S(G2105), .Z(new_n846));
  AOI22_X1  g421(.A1(G142), .A2(new_n470), .B1(new_n846), .B2(G2104), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n843), .B(new_n848), .Z(new_n849));
  NAND2_X1  g424(.A1(new_n842), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(G162), .B(new_n473), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n627), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n842), .A2(new_n849), .ZN(new_n854));
  AOI21_X1  g429(.A(G37), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n850), .A2(KEYINPUT102), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n850), .A2(KEYINPUT102), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n856), .A2(new_n857), .A3(new_n854), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n855), .B1(new_n858), .B2(new_n852), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g435(.A1(new_n825), .A2(G868), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT105), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n578), .A2(new_n862), .A3(new_n584), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n862), .B1(new_n578), .B2(new_n584), .ZN(new_n865));
  OAI21_X1  g440(.A(G166), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n585), .A2(KEYINPUT105), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n867), .A2(G303), .A3(new_n863), .ZN(new_n868));
  XNOR2_X1  g443(.A(G290), .B(new_n686), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n866), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT106), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n866), .A2(new_n868), .A3(new_n869), .A4(KEYINPUT106), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n866), .A2(new_n868), .ZN(new_n875));
  INV_X1    g450(.A(new_n869), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT42), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n831), .B(new_n610), .Z(new_n880));
  INV_X1    g455(.A(G299), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n601), .ZN(new_n882));
  NAND3_X1  g457(.A1(G299), .A2(new_n594), .A3(new_n600), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT104), .B1(new_n885), .B2(KEYINPUT41), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n602), .A2(KEYINPUT103), .A3(G299), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT103), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n887), .A2(new_n889), .A3(KEYINPUT41), .A4(new_n882), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n884), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n886), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n880), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n887), .A2(new_n889), .A3(new_n882), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n895), .B1(new_n897), .B2(new_n880), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n879), .B(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n861), .B1(new_n899), .B2(G868), .ZN(G295));
  AOI21_X1  g475(.A(new_n861), .B1(new_n899), .B2(G868), .ZN(G331));
  XNOR2_X1  g476(.A(G301), .B(G286), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n902), .B1(new_n829), .B2(new_n830), .ZN(new_n903));
  XOR2_X1   g478(.A(G301), .B(G286), .Z(new_n904));
  NAND2_X1  g479(.A1(new_n545), .A2(new_n546), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n825), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n904), .A2(new_n906), .A3(new_n828), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n903), .A2(new_n907), .A3(new_n896), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n903), .A2(new_n907), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n908), .B1(new_n894), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(G37), .B1(new_n910), .B2(new_n878), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n892), .B1(new_n903), .B2(new_n907), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n912), .A2(new_n896), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n884), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n913), .A2(new_n874), .A3(new_n877), .A4(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g493(.A1(new_n910), .A2(new_n878), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n919), .A2(new_n911), .A3(KEYINPUT43), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT44), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n911), .A2(KEYINPUT107), .A3(new_n915), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT107), .B1(new_n911), .B2(new_n915), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT43), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n919), .A2(new_n917), .A3(new_n911), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n921), .B1(new_n926), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g502(.A(G1981), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n575), .A2(new_n576), .A3(new_n928), .A4(new_n577), .ZN(new_n929));
  OAI21_X1  g504(.A(G1981), .B1(new_n582), .B2(new_n583), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT49), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n491), .A2(G2104), .ZN(new_n934));
  OAI211_X1 g509(.A(G126), .B(G2105), .C1(new_n483), .C2(new_n484), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(new_n494), .B2(new_n487), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n485), .A2(new_n486), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n462), .A2(KEYINPUT71), .A3(G138), .A4(new_n475), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n938), .A2(new_n939), .A3(KEYINPUT4), .ZN(new_n940));
  AOI21_X1  g515(.A(G1384), .B1(new_n937), .B2(new_n940), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n465), .A2(G40), .A3(new_n472), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G8), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n929), .A2(KEYINPUT49), .A3(new_n930), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n933), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n527), .A2(G87), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n529), .A2(G49), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n949), .A2(new_n950), .A3(G1976), .A4(new_n570), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n943), .A2(new_n951), .A3(G8), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT52), .ZN(new_n953));
  INV_X1    g528(.A(G1976), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT52), .B1(G288), .B2(new_n954), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n955), .A2(G8), .A3(new_n943), .A4(new_n951), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n948), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT55), .ZN(new_n960));
  NOR4_X1   g535(.A1(G166), .A2(new_n959), .A3(new_n960), .A4(new_n945), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(G303), .A2(G8), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n959), .B1(new_n963), .B2(new_n960), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n960), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n967));
  INV_X1    g542(.A(G1384), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n938), .A2(new_n939), .A3(KEYINPUT4), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n492), .A2(new_n488), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n967), .B(new_n968), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT111), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT50), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n465), .A2(G40), .A3(new_n472), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n967), .B1(new_n495), .B2(new_n968), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n976), .B1(new_n977), .B2(KEYINPUT111), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n975), .A2(new_n978), .A3(new_n756), .ZN(new_n979));
  XNOR2_X1  g554(.A(KEYINPUT108), .B(G1384), .ZN(new_n980));
  OAI211_X1 g555(.A(KEYINPUT45), .B(new_n980), .C1(new_n969), .C2(new_n970), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n981), .B(new_n942), .C1(new_n941), .C2(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n682), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n945), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n958), .B1(new_n966), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT118), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n979), .A2(new_n983), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(G8), .ZN(new_n988));
  NOR2_X1   g563(.A1(G166), .A2(new_n945), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT112), .B1(new_n989), .B2(KEYINPUT55), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(KEYINPUT55), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n961), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT113), .B1(new_n988), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n966), .A2(new_n994), .A3(new_n984), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n975), .A2(new_n978), .A3(new_n775), .ZN(new_n997));
  INV_X1    g572(.A(G1966), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n942), .B1(new_n941), .B2(KEYINPUT45), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT45), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n973), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n998), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n945), .B1(new_n997), .B2(new_n1002), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n1003), .A2(G168), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n986), .A2(KEYINPUT63), .A3(new_n996), .A4(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n1006), .B1(new_n977), .B2(new_n976), .ZN(new_n1007));
  OAI211_X1 g582(.A(KEYINPUT114), .B(new_n942), .C1(new_n941), .C2(new_n967), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(new_n971), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT115), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT115), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1007), .A2(new_n1008), .A3(new_n1011), .A4(new_n971), .ZN(new_n1012));
  AOI21_X1  g587(.A(G2090), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(new_n983), .ZN(new_n1014));
  OAI21_X1  g589(.A(G8), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(new_n992), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT116), .B1(new_n948), .B2(new_n957), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n933), .A2(new_n946), .A3(new_n947), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1018), .A2(new_n1019), .A3(new_n956), .A4(new_n953), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1016), .A2(new_n996), .A3(new_n1004), .A4(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT63), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1022), .A2(KEYINPUT117), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT117), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1005), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n993), .A2(new_n995), .A3(new_n958), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n686), .A2(new_n954), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n929), .B1(new_n948), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n946), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n993), .A2(new_n995), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n977), .B1(KEYINPUT111), .B2(new_n971), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n973), .A2(KEYINPUT111), .A3(KEYINPUT50), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n942), .ZN(new_n1035));
  OAI21_X1  g610(.A(KEYINPUT120), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1961), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n975), .A2(new_n978), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1036), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n976), .B1(new_n973), .B2(new_n1000), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n941), .A2(KEYINPUT45), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(new_n795), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT124), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1041), .A2(KEYINPUT124), .A3(new_n795), .A4(new_n1042), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1045), .A2(KEYINPUT53), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n982), .B2(G2078), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1040), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1050), .A2(KEYINPUT125), .A3(G171), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT125), .B1(new_n1050), .B2(G171), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1032), .B(new_n1016), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n997), .A2(new_n1002), .ZN(new_n1055));
  OAI211_X1 g630(.A(KEYINPUT123), .B(G8), .C1(new_n1055), .C2(G286), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(G168), .A2(new_n945), .ZN(new_n1059));
  OAI211_X1 g634(.A(KEYINPUT123), .B(KEYINPUT51), .C1(new_n1003), .C2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT62), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT122), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1003), .A2(new_n1063), .A3(G286), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1063), .B1(new_n1003), .B2(G286), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  AND3_X1   g641(.A1(new_n1061), .A2(new_n1062), .A3(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1054), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1055), .A2(G8), .A3(G286), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT122), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1003), .A2(new_n1063), .A3(G286), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1072), .B1(new_n1060), .B2(new_n1058), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n1073), .A2(new_n1062), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1031), .B1(new_n1068), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1032), .A2(new_n1016), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1050), .A2(G301), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT45), .B1(new_n495), .B2(new_n980), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1048), .B1(KEYINPUT126), .B2(new_n795), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(KEYINPUT126), .B2(new_n795), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1079), .A2(new_n976), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n981), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1040), .A2(G171), .A3(new_n1049), .A4(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1077), .B1(new_n1078), .B2(new_n1084), .ZN(new_n1085));
  NOR3_X1   g660(.A1(new_n1076), .A2(new_n1073), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1009), .A2(new_n801), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1009), .A2(KEYINPUT119), .A3(new_n801), .ZN(new_n1090));
  XNOR2_X1  g665(.A(KEYINPUT56), .B(G2072), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1041), .A2(new_n981), .A3(new_n1091), .ZN(new_n1092));
  XOR2_X1   g667(.A(G299), .B(KEYINPUT57), .Z(new_n1093));
  NAND4_X1  g668(.A1(new_n1089), .A2(new_n1090), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1036), .A2(new_n741), .A3(new_n1039), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n944), .A2(new_n739), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n601), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1094), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1093), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT119), .B1(new_n1009), .B2(new_n801), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1098), .A2(new_n1102), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n601), .A2(KEYINPUT60), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT58), .B(G1341), .Z(new_n1106));
  NAND2_X1  g681(.A1(new_n943), .A2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n982), .B2(G1996), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1108), .A2(new_n547), .A3(KEYINPUT121), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(KEYINPUT59), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1108), .A2(new_n547), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1111), .A2(new_n1112), .A3(KEYINPUT59), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1104), .A2(new_n1105), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1095), .A2(new_n601), .A3(new_n1096), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT60), .B1(new_n1117), .B2(new_n1097), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1102), .A2(KEYINPUT61), .A3(new_n1094), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1116), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(KEYINPUT61), .B1(new_n1102), .B2(new_n1094), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1103), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1053), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1040), .A2(new_n1049), .A3(new_n1083), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1123), .B(new_n1051), .C1(G171), .C2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n1077), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1086), .A2(new_n1122), .A3(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1026), .A2(new_n1075), .A3(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1079), .A2(new_n942), .ZN(new_n1129));
  INV_X1    g704(.A(G1996), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(new_n767), .ZN(new_n1132));
  XOR2_X1   g707(.A(new_n1132), .B(KEYINPUT110), .Z(new_n1133));
  XNOR2_X1  g708(.A(new_n737), .B(new_n739), .ZN(new_n1134));
  INV_X1    g709(.A(new_n767), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1134), .B1(new_n1130), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1133), .B1(new_n1129), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n705), .A2(new_n709), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n705), .A2(new_n709), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1129), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1137), .A2(new_n1140), .ZN(new_n1141));
  AND2_X1   g716(.A1(G290), .A2(G1986), .ZN(new_n1142));
  NOR2_X1   g717(.A1(G290), .A2(G1986), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1129), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1144), .B(KEYINPUT109), .ZN(new_n1145));
  AND2_X1   g720(.A1(new_n1141), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1128), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT127), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT46), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1148), .A2(KEYINPUT46), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1149), .B1(new_n1131), .B2(new_n1150), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1129), .ZN(new_n1153));
  OAI221_X1 g728(.A(new_n1151), .B1(new_n1131), .B2(new_n1149), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g729(.A(new_n1154), .B(KEYINPUT47), .Z(new_n1155));
  NAND2_X1  g730(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n737), .A2(G2067), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1153), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1143), .A2(new_n1129), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT48), .ZN(new_n1160));
  AOI211_X1 g735(.A(new_n1155), .B(new_n1158), .C1(new_n1141), .C2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1147), .A2(new_n1161), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g737(.A1(G229), .A2(G227), .A3(new_n460), .A4(G401), .ZN(new_n1164));
  AND2_X1   g738(.A1(new_n859), .A2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g739(.A1(new_n1165), .A2(new_n918), .A3(new_n920), .ZN(G225));
  INV_X1    g740(.A(G225), .ZN(G308));
endmodule


