//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n818, new_n819, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(KEYINPUT85), .B(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(G29gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g009(.A1(G29gat), .A2(G36gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n211), .B(KEYINPUT14), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT15), .ZN(new_n213));
  OR3_X1    g012(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G43gat), .B(G50gat), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n213), .B1(new_n210), .B2(new_n212), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n214), .A2(new_n217), .A3(new_n215), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G8gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(G15gat), .B(G22gat), .ZN(new_n221));
  OR2_X1    g020(.A1(new_n221), .A2(G1gat), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n220), .B1(new_n222), .B2(KEYINPUT86), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n221), .B1(new_n224), .B2(G1gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  OR2_X1    g025(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n223), .A2(new_n226), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n219), .B(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n231), .B(KEYINPUT13), .Z(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n229), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT17), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n216), .A2(new_n235), .A3(new_n218), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n235), .B1(new_n216), .B2(new_n218), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n234), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT87), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n219), .A2(KEYINPUT17), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n236), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT87), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(new_n243), .A3(new_n234), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n219), .A2(new_n229), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n240), .A2(new_n244), .A3(new_n245), .A4(new_n231), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT18), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n233), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n207), .B1(new_n249), .B2(KEYINPUT89), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT88), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT18), .B1(new_n246), .B2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n229), .B1(new_n241), .B2(new_n236), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n253), .A2(new_n243), .B1(new_n229), .B2(new_n219), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n254), .A2(KEYINPUT88), .A3(new_n231), .A4(new_n240), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n256), .A2(new_n249), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n250), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n248), .B1(new_n255), .B2(new_n252), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT89), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n206), .B1(new_n248), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G78gat), .B(G106gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(KEYINPUT31), .B(G50gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G141gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(G148gat), .ZN(new_n268));
  INV_X1    g067(.A(G148gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G141gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G155gat), .ZN(new_n272));
  INV_X1    g071(.A(G162gat), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT2), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G155gat), .B(G162gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT3), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n271), .A2(new_n276), .A3(new_n274), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT29), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G197gat), .B(G204gat), .ZN(new_n284));
  AND2_X1   g083(.A1(G211gat), .A2(G218gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n284), .B1(KEYINPUT22), .B2(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(G211gat), .A2(G218gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  OR2_X1    g088(.A1(new_n285), .A2(KEYINPUT22), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n290), .B(new_n284), .C1(new_n285), .C2(new_n287), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n283), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n286), .A2(new_n288), .ZN(new_n295));
  AOI21_X1  g094(.A(KEYINPUT29), .B1(new_n295), .B2(KEYINPUT79), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT79), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n289), .A2(new_n291), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT3), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n280), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n276), .B1(new_n274), .B2(new_n271), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n294), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(G228gat), .A2(G233gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT3), .B1(new_n292), .B2(new_n282), .ZN(new_n307));
  OR2_X1    g106(.A1(new_n307), .A2(new_n302), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n305), .B1(new_n283), .B2(new_n293), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G22gat), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n303), .A2(new_n305), .B1(new_n308), .B2(new_n309), .ZN(new_n313));
  INV_X1    g112(.A(G22gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n266), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n266), .B1(new_n315), .B2(KEYINPUT81), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT81), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n318), .B1(new_n313), .B2(new_n314), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT80), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n314), .B1(new_n311), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(new_n321), .B2(new_n311), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n316), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT70), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT64), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT24), .ZN(new_n327));
  INV_X1    g126(.A(G183gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G190gat), .ZN(new_n329));
  INV_X1    g128(.A(G190gat), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(G183gat), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n327), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n327), .A2(G183gat), .A3(G190gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n326), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G183gat), .B(G190gat), .ZN(new_n336));
  OAI211_X1 g135(.A(KEYINPUT64), .B(new_n333), .C1(new_n336), .C2(new_n327), .ZN(new_n337));
  NOR2_X1   g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT23), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n340), .B1(G169gat), .B2(G176gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n335), .A2(new_n337), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT25), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n333), .B1(new_n336), .B2(new_n327), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n341), .A2(KEYINPUT25), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n339), .A2(KEYINPUT65), .A3(new_n342), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT65), .B1(new_n339), .B2(new_n342), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n345), .A2(new_n346), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n328), .A2(KEYINPUT27), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT27), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n355), .A2(G183gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n354), .A2(new_n356), .A3(new_n330), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT66), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n357), .A2(new_n358), .A3(KEYINPUT28), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT28), .B1(new_n357), .B2(new_n358), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n338), .A2(KEYINPUT26), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT26), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n362), .B1(G169gat), .B2(G176gat), .ZN(new_n363));
  INV_X1    g162(.A(new_n342), .ZN(new_n364));
  OAI221_X1 g163(.A(new_n361), .B1(new_n328), .B2(new_n330), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  NOR3_X1   g164(.A1(new_n359), .A2(new_n360), .A3(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n282), .B1(new_n353), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(G226gat), .A2(G233gat), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n325), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n345), .A2(new_n346), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n349), .A2(new_n352), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n366), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n368), .B1(new_n372), .B2(KEYINPUT29), .ZN(new_n373));
  OR3_X1    g172(.A1(new_n359), .A2(new_n360), .A3(new_n365), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n343), .B1(new_n347), .B2(new_n326), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT25), .B1(new_n375), .B2(new_n337), .ZN(new_n376));
  NOR4_X1   g175(.A1(new_n347), .A2(new_n350), .A3(new_n351), .A4(new_n348), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n374), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n368), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n373), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n369), .B1(new_n381), .B2(new_n325), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT71), .B1(new_n382), .B2(new_n292), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT71), .ZN(new_n384));
  AOI21_X1  g183(.A(KEYINPUT70), .B1(new_n373), .B2(new_n380), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n384), .B(new_n293), .C1(new_n385), .C2(new_n369), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n381), .A2(new_n293), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G8gat), .B(G36gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(G64gat), .B(G92gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n391), .B(new_n392), .Z(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n390), .A2(new_n394), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n393), .A2(KEYINPUT30), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n379), .B1(new_n378), .B2(new_n282), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n372), .A2(new_n368), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n325), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n369), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n384), .B1(new_n401), .B2(new_n293), .ZN(new_n402));
  AOI211_X1 g201(.A(KEYINPUT71), .B(new_n292), .C1(new_n399), .C2(new_n400), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n389), .B(new_n396), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  AOI211_X1 g203(.A(new_n394), .B(new_n388), .C1(new_n383), .C2(new_n386), .ZN(new_n405));
  XOR2_X1   g204(.A(KEYINPUT72), .B(KEYINPUT30), .Z(new_n406));
  OAI211_X1 g205(.A(new_n395), .B(new_n404), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT78), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT3), .B1(new_n300), .B2(new_n301), .ZN(new_n409));
  XOR2_X1   g208(.A(G127gat), .B(G134gat), .Z(new_n410));
  XNOR2_X1  g209(.A(G113gat), .B(G120gat), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n410), .B1(KEYINPUT1), .B2(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(G113gat), .B(G120gat), .Z(new_n413));
  INV_X1    g212(.A(KEYINPUT1), .ZN(new_n414));
  XNOR2_X1  g213(.A(G127gat), .B(G134gat), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n412), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n409), .A2(new_n281), .A3(new_n417), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n412), .A2(new_n416), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n419), .A2(new_n302), .A3(KEYINPUT4), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n278), .A2(new_n412), .A3(new_n416), .A4(new_n280), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT4), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n418), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT5), .ZN(new_n425));
  NAND2_X1  g224(.A1(G225gat), .A2(G233gat), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n424), .A2(KEYINPUT76), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT76), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n418), .A2(new_n420), .A3(new_n426), .A4(new_n423), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n428), .B1(new_n429), .B2(KEYINPUT5), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n421), .B(KEYINPUT4), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT73), .ZN(new_n433));
  NAND4_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n426), .A4(new_n418), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n429), .A2(KEYINPUT73), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT74), .ZN(new_n436));
  INV_X1    g235(.A(new_n426), .ZN(new_n437));
  INV_X1    g236(.A(new_n421), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n278), .A2(new_n280), .B1(new_n412), .B2(new_n416), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n436), .B(new_n437), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n425), .B1(new_n441), .B2(KEYINPUT74), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n434), .A2(new_n435), .A3(new_n440), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n431), .A2(new_n443), .ZN(new_n444));
  XOR2_X1   g243(.A(G1gat), .B(G29gat), .Z(new_n445));
  XNOR2_X1  g244(.A(KEYINPUT75), .B(KEYINPUT0), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G57gat), .B(G85gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(new_n447), .B(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n444), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n408), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n449), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n453), .B1(new_n431), .B2(new_n443), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n454), .A2(KEYINPUT78), .A3(KEYINPUT6), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n431), .A2(new_n443), .A3(new_n453), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n450), .A2(new_n451), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT77), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n450), .A2(KEYINPUT77), .A3(new_n451), .A4(new_n457), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n456), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n324), .B1(new_n407), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT36), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT67), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n465), .B1(new_n353), .B2(new_n366), .ZN(new_n466));
  OAI211_X1 g265(.A(KEYINPUT67), .B(new_n374), .C1(new_n376), .C2(new_n377), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n417), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n378), .A2(new_n465), .A3(new_n419), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT34), .ZN(new_n471));
  NAND2_X1  g270(.A1(G227gat), .A2(G233gat), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n471), .B1(new_n470), .B2(new_n472), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(G15gat), .B(G43gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(KEYINPUT69), .ZN(new_n478));
  XNOR2_X1  g277(.A(G71gat), .B(G99gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n468), .A2(G227gat), .A3(G233gat), .A4(new_n469), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT33), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n484), .A2(KEYINPUT68), .B1(KEYINPUT32), .B2(new_n482), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n481), .A2(new_n483), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n482), .A2(KEYINPUT32), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT68), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n487), .B1(new_n484), .B2(new_n488), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n476), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n484), .A2(KEYINPUT68), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n482), .A2(KEYINPUT32), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n482), .A2(new_n483), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n494), .A2(new_n488), .A3(new_n480), .ZN(new_n495));
  INV_X1    g294(.A(new_n487), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n475), .B1(new_n493), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n464), .B1(new_n490), .B2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n476), .B1(new_n485), .B2(new_n489), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n493), .A2(new_n497), .A3(new_n475), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT36), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n388), .A2(KEYINPUT37), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(new_n402), .B2(new_n403), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n394), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT37), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n507), .B1(new_n387), .B2(new_n389), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT38), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n399), .A2(new_n292), .A3(new_n400), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT82), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n381), .A2(new_n511), .A3(new_n293), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n293), .B1(new_n397), .B2(new_n398), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT82), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n510), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(KEYINPUT38), .B1(new_n515), .B2(KEYINPUT37), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n505), .A2(new_n516), .A3(new_n394), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT83), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n452), .A2(new_n458), .A3(new_n455), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(new_n405), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT83), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n505), .A2(new_n516), .A3(new_n521), .A4(new_n394), .ZN(new_n522));
  AND4_X1   g321(.A1(new_n509), .A2(new_n518), .A3(new_n520), .A4(new_n522), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n424), .A2(new_n426), .ZN(new_n524));
  OR3_X1    g323(.A1(new_n438), .A2(new_n439), .A3(new_n437), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n524), .A2(KEYINPUT39), .A3(new_n525), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n526), .B(new_n453), .C1(KEYINPUT39), .C2(new_n524), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT40), .ZN(new_n528));
  AND2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n529), .A2(new_n530), .A3(new_n454), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n388), .B1(new_n383), .B2(new_n386), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n404), .B1(new_n393), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n406), .B1(new_n532), .B2(new_n393), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n531), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n324), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n463), .B(new_n503), .C1(new_n523), .C2(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n533), .A2(new_n534), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n324), .B1(new_n500), .B2(new_n501), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n460), .A2(new_n461), .ZN(new_n541));
  INV_X1    g340(.A(new_n456), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n539), .A2(new_n540), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT35), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT35), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n539), .A2(new_n540), .A3(new_n546), .A4(new_n519), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n538), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT84), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n538), .A2(KEYINPUT84), .A3(new_n548), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n263), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(G232gat), .A2(G233gat), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n554), .A2(KEYINPUT41), .ZN(new_n555));
  XNOR2_X1  g354(.A(G134gat), .B(G162gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n554), .A2(KEYINPUT41), .ZN(new_n559));
  INV_X1    g358(.A(new_n219), .ZN(new_n560));
  NAND2_X1  g359(.A1(G85gat), .A2(G92gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n561), .B(KEYINPUT7), .ZN(new_n562));
  NAND2_X1  g361(.A1(G99gat), .A2(G106gat), .ZN(new_n563));
  INV_X1    g362(.A(G85gat), .ZN(new_n564));
  INV_X1    g363(.A(G92gat), .ZN(new_n565));
  AOI22_X1  g364(.A1(KEYINPUT8), .A2(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G99gat), .B(G106gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n569), .A2(KEYINPUT92), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(KEYINPUT92), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n559), .B1(new_n560), .B2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  XOR2_X1   g373(.A(G190gat), .B(G218gat), .Z(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n242), .A2(new_n572), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n576), .B1(new_n574), .B2(new_n577), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n558), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n580), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(new_n557), .A3(new_n578), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT90), .ZN(new_n585));
  XNOR2_X1  g384(.A(G57gat), .B(G64gat), .ZN(new_n586));
  AOI21_X1  g385(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G71gat), .B(G78gat), .Z(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n590), .A2(KEYINPUT21), .ZN(new_n591));
  AND2_X1   g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G127gat), .B(G155gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT20), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n593), .B(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(G183gat), .B(G211gat), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n229), .B1(KEYINPUT21), .B2(new_n590), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n598), .A2(new_n602), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n584), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(G230gat), .ZN(new_n606));
  INV_X1    g405(.A(G233gat), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n570), .A2(KEYINPUT10), .A3(new_n590), .A4(new_n571), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n590), .B1(KEYINPUT93), .B2(new_n568), .ZN(new_n610));
  INV_X1    g409(.A(new_n569), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n569), .B(new_n590), .C1(KEYINPUT93), .C2(new_n568), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT94), .B(KEYINPUT10), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n608), .B1(new_n609), .B2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n608), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n612), .A2(new_n613), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  XOR2_X1   g419(.A(G120gat), .B(G148gat), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT95), .ZN(new_n622));
  XNOR2_X1  g421(.A(G176gat), .B(G204gat), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n622), .B(new_n623), .Z(new_n624));
  NAND2_X1  g423(.A1(new_n620), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT96), .ZN(new_n626));
  INV_X1    g425(.A(new_n624), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n617), .B(new_n627), .C1(new_n618), .C2(new_n619), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n620), .A2(KEYINPUT96), .A3(new_n624), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n605), .A2(KEYINPUT97), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(KEYINPUT97), .B1(new_n605), .B2(new_n631), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n553), .B(new_n462), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(KEYINPUT98), .B(G1gat), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(G1324gat));
  NOR2_X1   g435(.A1(new_n632), .A2(new_n633), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n637), .A2(new_n539), .ZN(new_n638));
  XOR2_X1   g437(.A(KEYINPUT16), .B(G8gat), .Z(new_n639));
  AND3_X1   g438(.A1(new_n553), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n220), .B1(new_n553), .B2(new_n638), .ZN(new_n641));
  OAI21_X1  g440(.A(KEYINPUT42), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n642), .B1(KEYINPUT42), .B2(new_n640), .ZN(G1325gat));
  OAI21_X1  g442(.A(new_n553), .B1(new_n632), .B2(new_n633), .ZN(new_n644));
  OAI21_X1  g443(.A(G15gat), .B1(new_n644), .B2(new_n503), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n490), .A2(new_n498), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n646), .A2(G15gat), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n645), .B1(new_n644), .B2(new_n647), .ZN(G1326gat));
  NOR2_X1   g447(.A1(new_n644), .A2(new_n536), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT43), .B(G22gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n649), .B(new_n650), .Z(G1327gat));
  INV_X1    g450(.A(new_n263), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n603), .A2(new_n604), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n654), .A2(new_n584), .A3(new_n631), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT99), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n538), .A2(KEYINPUT84), .A3(new_n548), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT84), .B1(new_n538), .B2(new_n548), .ZN(new_n658));
  OAI211_X1 g457(.A(new_n652), .B(new_n656), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n659), .A2(G29gat), .A3(new_n543), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n660), .A2(KEYINPUT45), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n581), .A2(new_n583), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n664), .B1(new_n657), .B2(new_n658), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n549), .A2(new_n584), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n663), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n631), .B(KEYINPUT100), .Z(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n669), .A2(new_n263), .A3(new_n653), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n665), .A2(new_n667), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(G29gat), .B1(new_n671), .B2(new_n543), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n660), .A2(KEYINPUT45), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n661), .A2(new_n672), .A3(new_n673), .ZN(G1328gat));
  INV_X1    g473(.A(KEYINPUT101), .ZN(new_n675));
  INV_X1    g474(.A(new_n208), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n539), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n675), .B1(new_n659), .B2(new_n678), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n553), .A2(KEYINPUT101), .A3(new_n656), .A4(new_n677), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n681), .A2(KEYINPUT46), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n676), .B1(new_n671), .B2(new_n539), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n681), .A2(KEYINPUT102), .A3(KEYINPUT46), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT102), .B1(new_n681), .B2(KEYINPUT46), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n682), .B(new_n683), .C1(new_n684), .C2(new_n685), .ZN(G1329gat));
  NOR3_X1   g485(.A1(new_n659), .A2(G43gat), .A3(new_n646), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT47), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n688), .A2(KEYINPUT103), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  OR2_X1    g489(.A1(new_n688), .A2(KEYINPUT103), .ZN(new_n691));
  OAI21_X1  g490(.A(G43gat), .B1(new_n671), .B2(new_n503), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n691), .B1(new_n690), .B2(new_n692), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(G1330gat));
  OAI21_X1  g494(.A(G50gat), .B1(new_n671), .B2(new_n536), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT104), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT48), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OR3_X1    g497(.A1(new_n659), .A2(G50gat), .A3(new_n536), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n696), .B(new_n699), .C1(new_n697), .C2(KEYINPUT48), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(G1331gat));
  NAND2_X1  g502(.A1(new_n263), .A2(new_n605), .ZN(new_n704));
  AOI211_X1 g503(.A(new_n668), .B(new_n704), .C1(new_n538), .C2(new_n548), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n462), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g506(.A(new_n539), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n709), .B(new_n710), .Z(G1333gat));
  INV_X1    g510(.A(new_n503), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n705), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n646), .A2(G71gat), .ZN(new_n714));
  AOI22_X1  g513(.A1(new_n713), .A2(G71gat), .B1(new_n705), .B2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(KEYINPUT105), .B(KEYINPUT50), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1334gat));
  NAND2_X1  g516(.A1(new_n705), .A2(new_n324), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT106), .B(G78gat), .Z(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1335gat));
  NOR2_X1   g519(.A1(new_n652), .A2(new_n653), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n549), .A2(KEYINPUT51), .A3(new_n584), .A4(new_n721), .ZN(new_n722));
  OR2_X1    g521(.A1(new_n722), .A2(KEYINPUT107), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(KEYINPUT107), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n549), .A2(new_n584), .A3(new_n721), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT51), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n723), .A2(new_n724), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT108), .ZN(new_n729));
  INV_X1    g528(.A(new_n631), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n462), .A2(new_n730), .A3(new_n564), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n665), .A2(new_n667), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n652), .A2(new_n653), .A3(new_n631), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n732), .A2(new_n543), .A3(new_n734), .ZN(new_n735));
  OAI22_X1  g534(.A1(new_n729), .A2(new_n731), .B1(new_n564), .B2(new_n735), .ZN(G1336gat));
  NOR3_X1   g535(.A1(new_n668), .A2(G92gat), .A3(new_n539), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n728), .A2(new_n737), .ZN(new_n738));
  NAND4_X1  g537(.A1(new_n665), .A2(new_n407), .A3(new_n667), .A4(new_n733), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT52), .B1(new_n739), .B2(G92gat), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT52), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n737), .B(KEYINPUT109), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n743), .B1(new_n727), .B2(new_n722), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n744), .B1(G92gat), .B2(new_n739), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n741), .B1(new_n742), .B2(new_n745), .ZN(G1337gat));
  NOR3_X1   g545(.A1(new_n646), .A2(G99gat), .A3(new_n631), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT110), .ZN(new_n748));
  INV_X1    g547(.A(G99gat), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n732), .A2(new_n503), .A3(new_n734), .ZN(new_n750));
  OAI22_X1  g549(.A1(new_n729), .A2(new_n748), .B1(new_n749), .B2(new_n750), .ZN(G1338gat));
  NOR3_X1   g550(.A1(new_n668), .A2(G106gat), .A3(new_n536), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n728), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n665), .A2(new_n324), .A3(new_n667), .A4(new_n733), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G106gat), .ZN(new_n755));
  XOR2_X1   g554(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n756));
  NAND3_X1  g555(.A1(new_n753), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n758));
  AND3_X1   g557(.A1(new_n754), .A2(new_n758), .A3(G106gat), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n758), .B1(new_n754), .B2(G106gat), .ZN(new_n760));
  INV_X1    g559(.A(new_n752), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n761), .B1(new_n727), .B2(new_n722), .ZN(new_n762));
  NOR3_X1   g561(.A1(new_n759), .A2(new_n760), .A3(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n757), .B1(new_n763), .B2(new_n764), .ZN(G1339gat));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n609), .A2(new_n615), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n767), .A2(new_n618), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT54), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n768), .A2(new_n769), .A3(new_n616), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n627), .B1(new_n616), .B2(new_n769), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n766), .B1(new_n770), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n617), .A2(KEYINPUT54), .ZN(new_n774));
  OAI211_X1 g573(.A(KEYINPUT55), .B(new_n771), .C1(new_n774), .C2(new_n768), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n773), .A2(new_n775), .A3(new_n628), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n250), .A2(new_n257), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n259), .A2(new_n261), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n231), .B1(new_n254), .B2(new_n240), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n780), .A2(KEYINPUT113), .B1(new_n230), .B2(new_n232), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n254), .A2(new_n240), .ZN(new_n782));
  INV_X1    g581(.A(new_n231), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(KEYINPUT113), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n205), .B1(new_n781), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n256), .A2(new_n249), .A3(new_n207), .ZN(new_n787));
  AND3_X1   g586(.A1(new_n730), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n662), .B1(new_n779), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n786), .A2(new_n787), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n776), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n786), .A2(new_n787), .A3(KEYINPUT114), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n792), .A2(new_n584), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n653), .B1(new_n789), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n704), .A2(new_n730), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n540), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n799), .A2(new_n407), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n798), .A2(new_n462), .A3(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n801), .B(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(G113gat), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n803), .A2(new_n804), .A3(new_n652), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n407), .A2(new_n543), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n798), .A2(new_n540), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G113gat), .B1(new_n807), .B2(new_n263), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(new_n808), .ZN(G1340gat));
  INV_X1    g608(.A(G120gat), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n803), .A2(new_n810), .A3(new_n730), .ZN(new_n811));
  OAI21_X1  g610(.A(G120gat), .B1(new_n807), .B2(new_n668), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n812), .A2(KEYINPUT116), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT116), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n814), .B(G120gat), .C1(new_n807), .C2(new_n668), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n811), .B1(new_n813), .B2(new_n816), .ZN(G1341gat));
  OAI21_X1  g616(.A(G127gat), .B1(new_n807), .B2(new_n654), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n654), .A2(G127gat), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n818), .B1(new_n801), .B2(new_n819), .ZN(G1342gat));
  NOR2_X1   g619(.A1(new_n662), .A2(G134gat), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  OR3_X1    g621(.A1(new_n801), .A2(KEYINPUT56), .A3(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(G134gat), .B1(new_n807), .B2(new_n662), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT56), .B1(new_n801), .B2(new_n822), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT117), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n823), .A2(new_n824), .A3(KEYINPUT117), .A4(new_n825), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(G1343gat));
  NAND2_X1  g629(.A1(new_n503), .A2(new_n806), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n796), .A2(new_n797), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(new_n833), .B2(new_n536), .ZN(new_n834));
  OAI211_X1 g633(.A(KEYINPUT57), .B(new_n324), .C1(new_n796), .C2(new_n797), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n831), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n267), .B1(new_n836), .B2(new_n652), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n833), .A2(new_n543), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n712), .A2(new_n536), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n407), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n263), .A2(G141gat), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT118), .ZN(new_n843));
  AND3_X1   g642(.A1(new_n838), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT58), .B1(new_n837), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n844), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT58), .ZN(new_n847));
  AOI211_X1 g646(.A(new_n263), .B(new_n831), .C1(new_n834), .C2(new_n835), .ZN(new_n848));
  OAI211_X1 g647(.A(new_n846), .B(new_n847), .C1(new_n848), .C2(new_n267), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n845), .A2(new_n849), .ZN(G1344gat));
  INV_X1    g649(.A(KEYINPUT122), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n793), .B1(new_n258), .B2(new_n262), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n730), .A2(new_n786), .A3(new_n787), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n584), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n775), .A2(new_n628), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n584), .A2(new_n855), .A3(new_n773), .A4(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT121), .B1(new_n776), .B2(new_n662), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n786), .A2(new_n787), .A3(KEYINPUT114), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT114), .B1(new_n786), .B2(new_n787), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n654), .B1(new_n854), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n263), .B1(new_n632), .B2(new_n633), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n536), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n835), .B1(new_n865), .B2(KEYINPUT57), .ZN(new_n866));
  INV_X1    g665(.A(new_n831), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n867), .A2(KEYINPUT120), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(KEYINPUT120), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n730), .A3(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n269), .B1(new_n866), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n851), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n792), .A2(new_n794), .A3(new_n858), .A4(new_n857), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n653), .B1(new_n789), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n864), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n324), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n832), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n870), .B1(new_n879), .B2(new_n835), .ZN(new_n880));
  OAI211_X1 g679(.A(KEYINPUT122), .B(KEYINPUT59), .C1(new_n880), .C2(new_n269), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n834), .A2(new_n835), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n730), .A3(new_n867), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n269), .A2(KEYINPUT59), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n874), .A2(new_n881), .A3(new_n885), .ZN(new_n886));
  AND4_X1   g685(.A1(new_n269), .A2(new_n838), .A3(new_n730), .A4(new_n841), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT119), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(G1345gat));
  NAND2_X1  g688(.A1(new_n838), .A2(new_n841), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n272), .A3(new_n653), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n836), .A2(new_n653), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n892), .B1(new_n893), .B2(new_n272), .ZN(G1346gat));
  NOR2_X1   g693(.A1(new_n662), .A2(G162gat), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n891), .A2(KEYINPUT123), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT123), .B1(new_n891), .B2(new_n895), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n836), .A2(new_n584), .ZN(new_n898));
  OAI22_X1  g697(.A1(new_n896), .A2(new_n897), .B1(new_n898), .B2(new_n273), .ZN(G1347gat));
  NOR2_X1   g698(.A1(new_n539), .A2(new_n462), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n540), .B(new_n900), .C1(new_n796), .C2(new_n797), .ZN(new_n901));
  INV_X1    g700(.A(G169gat), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n901), .A2(new_n902), .A3(new_n263), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n799), .A2(new_n539), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n798), .A2(new_n543), .A3(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n652), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n903), .B1(new_n907), .B2(new_n902), .ZN(G1348gat));
  OAI21_X1  g707(.A(G176gat), .B1(new_n901), .B2(new_n668), .ZN(new_n909));
  OR2_X1    g708(.A1(new_n631), .A2(G176gat), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n905), .B2(new_n910), .ZN(G1349gat));
  INV_X1    g710(.A(KEYINPUT60), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n912), .A2(KEYINPUT125), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n653), .A2(new_n354), .A3(new_n356), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n906), .B2(new_n914), .ZN(new_n915));
  OR3_X1    g714(.A1(new_n901), .A2(KEYINPUT124), .A3(new_n654), .ZN(new_n916));
  OAI21_X1  g715(.A(KEYINPUT124), .B1(new_n901), .B2(new_n654), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n916), .A2(G183gat), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n912), .A2(KEYINPUT125), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n915), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n915), .B2(new_n918), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n920), .A2(new_n921), .ZN(G1350gat));
  OAI21_X1  g721(.A(G190gat), .B1(new_n901), .B2(new_n662), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT61), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n906), .A2(new_n330), .A3(new_n584), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1351gat));
  NOR2_X1   g725(.A1(new_n840), .A2(new_n539), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n798), .A2(new_n543), .A3(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(G197gat), .B1(new_n929), .B2(new_n652), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n503), .A2(new_n900), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n931), .B1(new_n879), .B2(new_n835), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n652), .A2(G197gat), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(G1352gat));
  INV_X1    g733(.A(G204gat), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n730), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(KEYINPUT62), .B1(new_n928), .B2(new_n936), .ZN(new_n937));
  OR3_X1    g736(.A1(new_n928), .A2(KEYINPUT62), .A3(new_n936), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n932), .A2(new_n669), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n937), .B(new_n938), .C1(new_n939), .C2(new_n935), .ZN(G1353gat));
  OR3_X1    g739(.A1(new_n928), .A2(G211gat), .A3(new_n654), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n932), .A2(new_n653), .ZN(new_n942));
  OAI21_X1  g741(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n943));
  INV_X1    g742(.A(new_n943), .ZN(new_n944));
  AOI22_X1  g743(.A1(new_n942), .A2(new_n944), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n945));
  NAND2_X1  g744(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n946));
  AOI211_X1 g745(.A(new_n946), .B(new_n943), .C1(new_n932), .C2(new_n653), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n941), .B1(new_n945), .B2(new_n947), .ZN(G1354gat));
  AND2_X1   g747(.A1(new_n932), .A2(KEYINPUT127), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n584), .B1(new_n932), .B2(KEYINPUT127), .ZN(new_n950));
  OAI21_X1  g749(.A(G218gat), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OR3_X1    g750(.A1(new_n928), .A2(G218gat), .A3(new_n662), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1355gat));
endmodule


