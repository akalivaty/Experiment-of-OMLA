

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590;

  NOR2_X1 U325 ( .A1(n295), .A2(n407), .ZN(n408) );
  INV_X1 U326 ( .A(KEYINPUT74), .ZN(n359) );
  XOR2_X1 U327 ( .A(n399), .B(n398), .Z(n559) );
  XOR2_X1 U328 ( .A(n388), .B(KEYINPUT11), .Z(n293) );
  XOR2_X1 U329 ( .A(n395), .B(n394), .Z(n294) );
  XOR2_X1 U330 ( .A(n402), .B(KEYINPUT47), .Z(n295) );
  XNOR2_X1 U331 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U332 ( .A(n362), .B(n361), .ZN(n577) );
  NOR2_X1 U333 ( .A1(n534), .A2(n457), .ZN(n567) );
  XNOR2_X1 U334 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U335 ( .A(n461), .B(n460), .ZN(G1349GAT) );
  XOR2_X1 U336 ( .A(KEYINPUT88), .B(G176GAT), .Z(n297) );
  XNOR2_X1 U337 ( .A(KEYINPUT20), .B(KEYINPUT87), .ZN(n296) );
  XNOR2_X1 U338 ( .A(n297), .B(n296), .ZN(n313) );
  XOR2_X1 U339 ( .A(KEYINPUT85), .B(G99GAT), .Z(n299) );
  XNOR2_X1 U340 ( .A(G113GAT), .B(G134GAT), .ZN(n298) );
  XNOR2_X1 U341 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U342 ( .A(n300), .B(G190GAT), .Z(n302) );
  XOR2_X1 U343 ( .A(G120GAT), .B(G71GAT), .Z(n354) );
  XNOR2_X1 U344 ( .A(G43GAT), .B(n354), .ZN(n301) );
  XNOR2_X1 U345 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U346 ( .A(KEYINPUT0), .B(G127GAT), .Z(n428) );
  XOR2_X1 U347 ( .A(n428), .B(KEYINPUT86), .Z(n304) );
  NAND2_X1 U348 ( .A1(G227GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U349 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U350 ( .A(n306), .B(n305), .Z(n311) );
  XOR2_X1 U351 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n308) );
  XNOR2_X1 U352 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n307) );
  XNOR2_X1 U353 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U354 ( .A(G169GAT), .B(n309), .Z(n328) );
  XNOR2_X1 U355 ( .A(G15GAT), .B(n328), .ZN(n310) );
  XNOR2_X1 U356 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X2 U357 ( .A(n313), .B(n312), .Z(n534) );
  XOR2_X1 U358 ( .A(KEYINPUT90), .B(G218GAT), .Z(n315) );
  XNOR2_X1 U359 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n314) );
  XNOR2_X1 U360 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U361 ( .A(G197GAT), .B(n316), .Z(n452) );
  XOR2_X1 U362 ( .A(G92GAT), .B(G64GAT), .Z(n318) );
  XNOR2_X1 U363 ( .A(G204GAT), .B(KEYINPUT77), .ZN(n317) );
  XNOR2_X1 U364 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U365 ( .A(G176GAT), .B(n319), .Z(n353) );
  XNOR2_X1 U366 ( .A(n452), .B(n353), .ZN(n326) );
  XOR2_X1 U367 ( .A(G36GAT), .B(G190GAT), .Z(n390) );
  XOR2_X1 U368 ( .A(KEYINPUT102), .B(KEYINPUT100), .Z(n321) );
  XNOR2_X1 U369 ( .A(G8GAT), .B(KEYINPUT101), .ZN(n320) );
  XNOR2_X1 U370 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U371 ( .A(n390), .B(n322), .Z(n324) );
  NAND2_X1 U372 ( .A1(G226GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U373 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U375 ( .A(n328), .B(n327), .ZN(n498) );
  XOR2_X1 U376 ( .A(G57GAT), .B(KEYINPUT13), .Z(n346) );
  XOR2_X1 U377 ( .A(n346), .B(G78GAT), .Z(n330) );
  XOR2_X1 U378 ( .A(G15GAT), .B(G8GAT), .Z(n371) );
  XNOR2_X1 U379 ( .A(n371), .B(G211GAT), .ZN(n329) );
  XNOR2_X1 U380 ( .A(n330), .B(n329), .ZN(n334) );
  XOR2_X1 U381 ( .A(KEYINPUT12), .B(KEYINPUT84), .Z(n332) );
  XNOR2_X1 U382 ( .A(G1GAT), .B(KEYINPUT83), .ZN(n331) );
  XNOR2_X1 U383 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U384 ( .A(n334), .B(n333), .Z(n336) );
  XNOR2_X1 U385 ( .A(G22GAT), .B(G155GAT), .ZN(n335) );
  XNOR2_X1 U386 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U387 ( .A(KEYINPUT14), .B(KEYINPUT82), .Z(n338) );
  NAND2_X1 U388 ( .A1(G231GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U389 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U390 ( .A(n340), .B(n339), .Z(n345) );
  XOR2_X1 U391 ( .A(G64GAT), .B(G71GAT), .Z(n342) );
  XNOR2_X1 U392 ( .A(G183GAT), .B(G127GAT), .ZN(n341) );
  XNOR2_X1 U393 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U394 ( .A(n343), .B(KEYINPUT15), .ZN(n344) );
  XNOR2_X1 U395 ( .A(n345), .B(n344), .ZN(n564) );
  INV_X1 U396 ( .A(KEYINPUT41), .ZN(n363) );
  XOR2_X1 U397 ( .A(G99GAT), .B(G85GAT), .Z(n391) );
  XOR2_X1 U398 ( .A(n346), .B(n391), .Z(n348) );
  NAND2_X1 U399 ( .A1(G230GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U401 ( .A(KEYINPUT33), .B(KEYINPUT78), .Z(n350) );
  XNOR2_X1 U402 ( .A(KEYINPUT76), .B(KEYINPUT32), .ZN(n349) );
  XNOR2_X1 U403 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U404 ( .A(n352), .B(n351), .Z(n356) );
  XNOR2_X1 U405 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U406 ( .A(n356), .B(n355), .ZN(n362) );
  XOR2_X1 U407 ( .A(G78GAT), .B(G148GAT), .Z(n358) );
  XNOR2_X1 U408 ( .A(G106GAT), .B(KEYINPUT75), .ZN(n357) );
  XNOR2_X1 U409 ( .A(n358), .B(n357), .ZN(n444) );
  XNOR2_X1 U410 ( .A(n444), .B(KEYINPUT31), .ZN(n360) );
  XNOR2_X1 U411 ( .A(n363), .B(n577), .ZN(n551) );
  XOR2_X1 U412 ( .A(KEYINPUT73), .B(KEYINPUT68), .Z(n365) );
  XNOR2_X1 U413 ( .A(KEYINPUT69), .B(KEYINPUT29), .ZN(n364) );
  XNOR2_X1 U414 ( .A(n365), .B(n364), .ZN(n382) );
  XOR2_X1 U415 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n367) );
  XNOR2_X1 U416 ( .A(G36GAT), .B(G50GAT), .ZN(n366) );
  XNOR2_X1 U417 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U418 ( .A(n368), .B(G197GAT), .Z(n370) );
  XOR2_X1 U419 ( .A(G113GAT), .B(G1GAT), .Z(n429) );
  XNOR2_X1 U420 ( .A(G169GAT), .B(n429), .ZN(n369) );
  XNOR2_X1 U421 ( .A(n370), .B(n369), .ZN(n375) );
  XOR2_X1 U422 ( .A(n371), .B(KEYINPUT71), .Z(n373) );
  NAND2_X1 U423 ( .A1(G229GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U424 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U425 ( .A(n375), .B(n374), .Z(n380) );
  XOR2_X1 U426 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n377) );
  XNOR2_X1 U427 ( .A(G43GAT), .B(G29GAT), .ZN(n376) );
  XNOR2_X1 U428 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U429 ( .A(KEYINPUT72), .B(n378), .Z(n396) );
  XOR2_X1 U430 ( .A(G141GAT), .B(G22GAT), .Z(n448) );
  XNOR2_X1 U431 ( .A(n396), .B(n448), .ZN(n379) );
  XNOR2_X1 U432 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U433 ( .A(n382), .B(n381), .ZN(n561) );
  NAND2_X1 U434 ( .A1(n551), .A2(n561), .ZN(n383) );
  XNOR2_X1 U435 ( .A(KEYINPUT46), .B(n383), .ZN(n400) );
  XOR2_X1 U436 ( .A(KEYINPUT9), .B(KEYINPUT81), .Z(n385) );
  XNOR2_X1 U437 ( .A(G106GAT), .B(G92GAT), .ZN(n384) );
  XNOR2_X1 U438 ( .A(n385), .B(n384), .ZN(n399) );
  XOR2_X1 U439 ( .A(KEYINPUT65), .B(KEYINPUT67), .Z(n387) );
  XNOR2_X1 U440 ( .A(KEYINPUT10), .B(KEYINPUT66), .ZN(n386) );
  XNOR2_X1 U441 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U442 ( .A(G50GAT), .B(G162GAT), .Z(n442) );
  XNOR2_X1 U443 ( .A(G218GAT), .B(n442), .ZN(n389) );
  XNOR2_X1 U444 ( .A(n293), .B(n389), .ZN(n395) );
  XOR2_X1 U445 ( .A(n391), .B(n390), .Z(n393) );
  NAND2_X1 U446 ( .A1(G232GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U447 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U448 ( .A(G134GAT), .B(KEYINPUT80), .Z(n413) );
  XNOR2_X1 U449 ( .A(n396), .B(n413), .ZN(n397) );
  XNOR2_X1 U450 ( .A(n294), .B(n397), .ZN(n398) );
  NAND2_X1 U451 ( .A1(n400), .A2(n559), .ZN(n401) );
  NOR2_X1 U452 ( .A1(n564), .A2(n401), .ZN(n402) );
  INV_X1 U453 ( .A(n564), .ZN(n583) );
  XNOR2_X1 U454 ( .A(n559), .B(KEYINPUT36), .ZN(n588) );
  NOR2_X1 U455 ( .A1(n583), .A2(n588), .ZN(n403) );
  XNOR2_X1 U456 ( .A(n403), .B(KEYINPUT45), .ZN(n404) );
  INV_X1 U457 ( .A(n561), .ZN(n573) );
  NAND2_X1 U458 ( .A1(n404), .A2(n573), .ZN(n405) );
  NOR2_X1 U459 ( .A1(n577), .A2(n405), .ZN(n406) );
  XNOR2_X1 U460 ( .A(KEYINPUT114), .B(n406), .ZN(n407) );
  XNOR2_X1 U461 ( .A(KEYINPUT48), .B(n408), .ZN(n531) );
  NOR2_X1 U462 ( .A1(n498), .A2(n531), .ZN(n409) );
  XNOR2_X1 U463 ( .A(n409), .B(KEYINPUT54), .ZN(n438) );
  XOR2_X1 U464 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n411) );
  NAND2_X1 U465 ( .A1(G225GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U466 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U467 ( .A(n413), .B(n412), .ZN(n437) );
  XOR2_X1 U468 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n415) );
  XNOR2_X1 U469 ( .A(KEYINPUT4), .B(KEYINPUT93), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U471 ( .A(KEYINPUT98), .B(G57GAT), .Z(n417) );
  XNOR2_X1 U472 ( .A(G141GAT), .B(G120GAT), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U474 ( .A(n419), .B(n418), .Z(n427) );
  XOR2_X1 U475 ( .A(KEYINPUT3), .B(KEYINPUT92), .Z(n421) );
  XNOR2_X1 U476 ( .A(KEYINPUT91), .B(G155GAT), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U478 ( .A(KEYINPUT2), .B(n422), .Z(n453) );
  XOR2_X1 U479 ( .A(KEYINPUT1), .B(KEYINPUT96), .Z(n424) );
  XNOR2_X1 U480 ( .A(KEYINPUT99), .B(KEYINPUT97), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U482 ( .A(n453), .B(n425), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n433) );
  XOR2_X1 U484 ( .A(G162GAT), .B(G148GAT), .Z(n431) );
  XNOR2_X1 U485 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U487 ( .A(n433), .B(n432), .Z(n435) );
  XNOR2_X1 U488 ( .A(G29GAT), .B(G85GAT), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U490 ( .A(n437), .B(n436), .ZN(n495) );
  NAND2_X1 U491 ( .A1(n438), .A2(n495), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n439), .B(KEYINPUT64), .ZN(n570) );
  XOR2_X1 U493 ( .A(KEYINPUT22), .B(KEYINPUT89), .Z(n441) );
  XNOR2_X1 U494 ( .A(G204GAT), .B(KEYINPUT23), .ZN(n440) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n443) );
  XOR2_X1 U496 ( .A(n443), .B(n442), .Z(n450) );
  XOR2_X1 U497 ( .A(KEYINPUT24), .B(n444), .Z(n446) );
  NAND2_X1 U498 ( .A1(G228GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U499 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U500 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U501 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U502 ( .A(n452), .B(n451), .ZN(n455) );
  INV_X1 U503 ( .A(n453), .ZN(n454) );
  XNOR2_X1 U504 ( .A(n455), .B(n454), .ZN(n473) );
  NOR2_X1 U505 ( .A1(n570), .A2(n473), .ZN(n456) );
  XNOR2_X1 U506 ( .A(n456), .B(KEYINPUT55), .ZN(n457) );
  NAND2_X1 U507 ( .A1(n567), .A2(n551), .ZN(n461) );
  XOR2_X1 U508 ( .A(KEYINPUT122), .B(KEYINPUT56), .Z(n459) );
  XNOR2_X1 U509 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n458) );
  INV_X1 U510 ( .A(n495), .ZN(n518) );
  NOR2_X1 U511 ( .A1(n577), .A2(n573), .ZN(n462) );
  XNOR2_X1 U512 ( .A(n462), .B(KEYINPUT79), .ZN(n492) );
  INV_X1 U513 ( .A(n559), .ZN(n566) );
  NOR2_X1 U514 ( .A1(n566), .A2(n583), .ZN(n463) );
  XNOR2_X1 U515 ( .A(n463), .B(KEYINPUT16), .ZN(n479) );
  NOR2_X1 U516 ( .A1(n534), .A2(n498), .ZN(n464) );
  XNOR2_X1 U517 ( .A(n464), .B(KEYINPUT104), .ZN(n465) );
  NOR2_X1 U518 ( .A1(n473), .A2(n465), .ZN(n466) );
  XOR2_X1 U519 ( .A(KEYINPUT25), .B(n466), .Z(n470) );
  XNOR2_X1 U520 ( .A(KEYINPUT27), .B(n498), .ZN(n474) );
  XOR2_X1 U521 ( .A(KEYINPUT26), .B(KEYINPUT103), .Z(n468) );
  NAND2_X1 U522 ( .A1(n534), .A2(n473), .ZN(n467) );
  XNOR2_X1 U523 ( .A(n468), .B(n467), .ZN(n571) );
  NOR2_X1 U524 ( .A1(n474), .A2(n571), .ZN(n469) );
  NOR2_X1 U525 ( .A1(n470), .A2(n469), .ZN(n471) );
  NOR2_X1 U526 ( .A1(n518), .A2(n471), .ZN(n472) );
  XOR2_X1 U527 ( .A(KEYINPUT105), .B(n472), .Z(n477) );
  XNOR2_X1 U528 ( .A(KEYINPUT28), .B(n473), .ZN(n525) );
  NOR2_X1 U529 ( .A1(n495), .A2(n474), .ZN(n529) );
  NAND2_X1 U530 ( .A1(n534), .A2(n529), .ZN(n475) );
  NOR2_X1 U531 ( .A1(n525), .A2(n475), .ZN(n476) );
  NOR2_X1 U532 ( .A1(n477), .A2(n476), .ZN(n489) );
  INV_X1 U533 ( .A(n489), .ZN(n478) );
  NAND2_X1 U534 ( .A1(n479), .A2(n478), .ZN(n505) );
  NOR2_X1 U535 ( .A1(n492), .A2(n505), .ZN(n487) );
  NAND2_X1 U536 ( .A1(n518), .A2(n487), .ZN(n483) );
  XOR2_X1 U537 ( .A(KEYINPUT107), .B(KEYINPUT34), .Z(n481) );
  XNOR2_X1 U538 ( .A(G1GAT), .B(KEYINPUT106), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n483), .B(n482), .ZN(G1324GAT) );
  INV_X1 U541 ( .A(n498), .ZN(n520) );
  NAND2_X1 U542 ( .A1(n487), .A2(n520), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n484), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U544 ( .A(G15GAT), .B(KEYINPUT35), .Z(n486) );
  INV_X1 U545 ( .A(n534), .ZN(n523) );
  NAND2_X1 U546 ( .A1(n487), .A2(n523), .ZN(n485) );
  XNOR2_X1 U547 ( .A(n486), .B(n485), .ZN(G1326GAT) );
  NAND2_X1 U548 ( .A1(n487), .A2(n525), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n488), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U550 ( .A1(n489), .A2(n588), .ZN(n490) );
  NAND2_X1 U551 ( .A1(n583), .A2(n490), .ZN(n491) );
  XOR2_X1 U552 ( .A(KEYINPUT37), .B(n491), .Z(n517) );
  NOR2_X1 U553 ( .A1(n492), .A2(n517), .ZN(n494) );
  XOR2_X1 U554 ( .A(KEYINPUT38), .B(KEYINPUT108), .Z(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n502) );
  NOR2_X1 U556 ( .A1(n495), .A2(n502), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n496), .B(KEYINPUT39), .ZN(n497) );
  XNOR2_X1 U558 ( .A(G29GAT), .B(n497), .ZN(G1328GAT) );
  NOR2_X1 U559 ( .A1(n498), .A2(n502), .ZN(n499) );
  XOR2_X1 U560 ( .A(G36GAT), .B(n499), .Z(G1329GAT) );
  NOR2_X1 U561 ( .A1(n534), .A2(n502), .ZN(n500) );
  XOR2_X1 U562 ( .A(KEYINPUT40), .B(n500), .Z(n501) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n501), .ZN(G1330GAT) );
  INV_X1 U564 ( .A(n525), .ZN(n532) );
  NOR2_X1 U565 ( .A1(n532), .A2(n502), .ZN(n504) );
  XNOR2_X1 U566 ( .A(G50GAT), .B(KEYINPUT109), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(G1331GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n507) );
  NAND2_X1 U569 ( .A1(n573), .A2(n551), .ZN(n516) );
  NOR2_X1 U570 ( .A1(n516), .A2(n505), .ZN(n511) );
  NAND2_X1 U571 ( .A1(n511), .A2(n518), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U573 ( .A(G57GAT), .B(n508), .Z(G1332GAT) );
  NAND2_X1 U574 ( .A1(n511), .A2(n520), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n509), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U576 ( .A1(n523), .A2(n511), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n510), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n513) );
  NAND2_X1 U579 ( .A1(n511), .A2(n525), .ZN(n512) );
  XNOR2_X1 U580 ( .A(n513), .B(n512), .ZN(n515) );
  XOR2_X1 U581 ( .A(G78GAT), .B(KEYINPUT112), .Z(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(G1335GAT) );
  NOR2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n526) );
  NAND2_X1 U584 ( .A1(n526), .A2(n518), .ZN(n519) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(n519), .ZN(G1336GAT) );
  XOR2_X1 U586 ( .A(G92GAT), .B(KEYINPUT113), .Z(n522) );
  NAND2_X1 U587 ( .A1(n526), .A2(n520), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n523), .A2(n526), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n524), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n527), .B(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n528), .ZN(G1339GAT) );
  INV_X1 U594 ( .A(n529), .ZN(n530) );
  NOR2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n546) );
  NAND2_X1 U596 ( .A1(n546), .A2(n532), .ZN(n533) );
  NOR2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n541), .A2(n561), .ZN(n535) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U601 ( .A1(n541), .A2(n551), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n539) );
  NAND2_X1 U604 ( .A1(n541), .A2(n564), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U606 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT51), .B(KEYINPUT116), .Z(n543) );
  NAND2_X1 U608 ( .A1(n541), .A2(n566), .ZN(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(n544), .ZN(G1343GAT) );
  INV_X1 U611 ( .A(n571), .ZN(n545) );
  NAND2_X1 U612 ( .A1(n546), .A2(n545), .ZN(n558) );
  NOR2_X1 U613 ( .A1(n573), .A2(n558), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT52), .B(KEYINPUT118), .Z(n550) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n554) );
  INV_X1 U619 ( .A(n551), .ZN(n552) );
  NOR2_X1 U620 ( .A1(n552), .A2(n558), .ZN(n553) );
  XOR2_X1 U621 ( .A(n554), .B(n553), .Z(G1345GAT) );
  NOR2_X1 U622 ( .A1(n583), .A2(n558), .ZN(n556) );
  XNOR2_X1 U623 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(G155GAT), .B(n557), .ZN(G1346GAT) );
  NOR2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U627 ( .A(G162GAT), .B(n560), .Z(G1347GAT) );
  NAND2_X1 U628 ( .A1(n567), .A2(n561), .ZN(n563) );
  XOR2_X1 U629 ( .A(G169GAT), .B(KEYINPUT121), .Z(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1348GAT) );
  NAND2_X1 U631 ( .A1(n567), .A2(n564), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U633 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n569) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1351GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n572), .B(KEYINPUT123), .ZN(n587) );
  NOR2_X1 U638 ( .A1(n573), .A2(n587), .ZN(n575) );
  XNOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(G197GAT), .B(n576), .ZN(G1352GAT) );
  INV_X1 U642 ( .A(n577), .ZN(n578) );
  NOR2_X1 U643 ( .A1(n587), .A2(n578), .ZN(n582) );
  XOR2_X1 U644 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n580) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1353GAT) );
  NOR2_X1 U648 ( .A1(n583), .A2(n587), .ZN(n584) );
  XOR2_X1 U649 ( .A(G211GAT), .B(n584), .Z(G1354GAT) );
  XOR2_X1 U650 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n586) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(n590) );
  NOR2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U654 ( .A(n590), .B(n589), .Z(G1355GAT) );
endmodule

