//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 1 0 0 0 1 1 1 1 0 1 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:02 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1245, new_n1246, new_n1247, new_n1248, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XOR2_X1   g0003(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  OAI21_X1  g0014(.A(G50), .B1(G58), .B2(G68), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n209), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n211), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n214), .B(new_n219), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G226), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G58), .B(G77), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(KEYINPUT21), .ZN(new_n245));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  INV_X1    g0046(.A(G116), .ZN(new_n247));
  AOI22_X1  g0047(.A1(new_n246), .A2(new_n217), .B1(G20), .B2(new_n247), .ZN(new_n248));
  AOI21_X1  g0048(.A(G20), .B1(G33), .B2(G283), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G97), .ZN(new_n251));
  AND3_X1   g0051(.A1(new_n249), .A2(new_n251), .A3(KEYINPUT83), .ZN(new_n252));
  AOI21_X1  g0052(.A(KEYINPUT83), .B1(new_n249), .B2(new_n251), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n248), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OAI211_X1 g0056(.A(KEYINPUT20), .B(new_n248), .C1(new_n252), .C2(new_n253), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G116), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n246), .A2(new_n217), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n208), .A2(G33), .ZN(new_n263));
  AND3_X1   g0063(.A1(new_n262), .A2(new_n259), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n260), .B1(new_n264), .B2(G116), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G169), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT82), .ZN(new_n268));
  AND2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  OAI211_X1 g0070(.A(G264), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  OAI211_X1 g0072(.A(G257), .B(new_n272), .C1(new_n269), .C2(new_n270), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(new_n250), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(G303), .A3(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n271), .A2(new_n273), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G41), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n208), .B(G45), .C1(new_n281), .C2(KEYINPUT5), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT77), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G45), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n285), .A2(G1), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT5), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G41), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(KEYINPUT77), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n281), .A2(KEYINPUT5), .ZN(new_n290));
  INV_X1    g0090(.A(G274), .ZN(new_n291));
  AND2_X1   g0091(.A1(G1), .A2(G13), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G41), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND4_X1  g0094(.A1(new_n284), .A2(new_n289), .A3(new_n290), .A4(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n286), .A2(new_n290), .A3(new_n288), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n292), .A2(new_n293), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(G270), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n268), .B1(new_n280), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n278), .A2(new_n279), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n301), .A2(KEYINPUT82), .A3(new_n295), .A4(new_n298), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n245), .B1(new_n267), .B2(new_n303), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n301), .A2(G179), .A3(new_n295), .A4(new_n298), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n266), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(new_n258), .B2(new_n265), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n309), .A2(KEYINPUT21), .A3(new_n300), .A4(new_n302), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n304), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n300), .A2(G200), .A3(new_n302), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n313), .B1(new_n300), .B2(new_n302), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n312), .A2(new_n314), .A3(new_n266), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n262), .A2(new_n259), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n208), .A2(G20), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G50), .ZN(new_n319));
  OAI22_X1  g0119(.A1(new_n317), .A2(new_n319), .B1(G50), .B2(new_n259), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n320), .B(KEYINPUT68), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n204), .A2(new_n209), .ZN(new_n322));
  XNOR2_X1  g0122(.A(KEYINPUT8), .B(G58), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n209), .A2(G33), .ZN(new_n324));
  INV_X1    g0124(.A(G150), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n209), .A2(new_n250), .ZN(new_n326));
  OAI22_X1  g0126(.A1(new_n323), .A2(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n261), .B1(new_n322), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n321), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g0129(.A(new_n329), .B(KEYINPUT9), .ZN(new_n330));
  AOI21_X1  g0130(.A(G1698), .B1(new_n275), .B2(new_n276), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n269), .A2(new_n270), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n331), .A2(G222), .B1(new_n332), .B2(G77), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n275), .A2(new_n276), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(G1698), .ZN(new_n335));
  XOR2_X1   g0135(.A(KEYINPUT67), .B(G223), .Z(new_n336));
  OAI21_X1  g0136(.A(new_n333), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n279), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n294), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G226), .ZN(new_n342));
  NOR2_X1   g0142(.A1(G41), .A2(G45), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT66), .B1(new_n343), .B2(G1), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT66), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n345), .B(new_n208), .C1(G41), .C2(G45), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n344), .A2(new_n297), .A3(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n338), .B(new_n341), .C1(new_n342), .C2(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n348), .A2(new_n313), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(G200), .B2(new_n348), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n330), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT10), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT10), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n330), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n348), .A2(G179), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n348), .A2(new_n308), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(new_n329), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n356), .B1(new_n359), .B2(KEYINPUT69), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(KEYINPUT69), .B2(new_n359), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n344), .A2(G244), .A3(new_n297), .A4(new_n346), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n341), .ZN(new_n363));
  OAI211_X1 g0163(.A(G232), .B(new_n272), .C1(new_n269), .C2(new_n270), .ZN(new_n364));
  OAI211_X1 g0164(.A(G238), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n275), .A2(G107), .A3(new_n276), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n363), .B1(new_n279), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G190), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n318), .A2(G77), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n317), .A2(new_n370), .B1(G77), .B2(new_n259), .ZN(new_n371));
  INV_X1    g0171(.A(G58), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT8), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT8), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(G58), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n326), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n209), .A2(new_n205), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT70), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT70), .ZN(new_n379));
  OAI221_X1 g0179(.A(new_n379), .B1(new_n209), .B2(new_n205), .C1(new_n323), .C2(new_n326), .ZN(new_n380));
  XNOR2_X1  g0180(.A(KEYINPUT15), .B(G87), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n381), .A2(new_n324), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n378), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n371), .B1(new_n384), .B2(new_n261), .ZN(new_n385));
  AND2_X1   g0185(.A1(new_n362), .A2(new_n341), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n367), .A2(new_n279), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(G200), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n369), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n388), .A2(G179), .ZN(new_n391));
  OAI22_X1  g0191(.A1(new_n323), .A2(new_n326), .B1(new_n209), .B2(new_n205), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n382), .B1(new_n392), .B2(KEYINPUT70), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n262), .B1(new_n393), .B2(new_n380), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n394), .A2(new_n371), .B1(new_n368), .B2(G169), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n391), .B1(new_n395), .B2(KEYINPUT71), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n388), .A2(new_n308), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT71), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n397), .B(new_n398), .C1(new_n394), .C2(new_n371), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n390), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n355), .A2(new_n361), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n259), .ZN(new_n402));
  INV_X1    g0202(.A(G68), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g0204(.A(new_n404), .B(KEYINPUT12), .ZN(new_n405));
  INV_X1    g0205(.A(new_n326), .ZN(new_n406));
  AOI22_X1  g0206(.A1(new_n406), .A2(G50), .B1(G20), .B2(new_n403), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n205), .B2(new_n324), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(KEYINPUT11), .A3(new_n261), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n318), .A2(G68), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n405), .B(new_n409), .C1(new_n317), .C2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT11), .B1(new_n408), .B2(new_n261), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT14), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT13), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n342), .A2(G1698), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n269), .B2(new_n270), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT72), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G33), .A2(G97), .ZN(new_n420));
  OAI211_X1 g0220(.A(G232), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT72), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n417), .B(new_n422), .C1(new_n270), .C2(new_n269), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n419), .A2(new_n420), .A3(new_n421), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n279), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT73), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n347), .A2(new_n426), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n339), .A2(KEYINPUT66), .B1(new_n292), .B2(new_n293), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n428), .A2(KEYINPUT73), .A3(new_n346), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n427), .A2(new_n429), .A3(G238), .ZN(new_n430));
  AND4_X1   g0230(.A1(new_n416), .A2(new_n425), .A3(new_n430), .A4(new_n341), .ZN(new_n431));
  NOR3_X1   g0231(.A1(new_n279), .A2(new_n291), .A3(new_n339), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n424), .B2(new_n279), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n416), .B1(new_n433), .B2(new_n430), .ZN(new_n434));
  OAI211_X1 g0234(.A(new_n415), .B(G169), .C1(new_n431), .C2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n425), .A2(new_n430), .A3(new_n341), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT13), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n433), .A2(new_n416), .A3(new_n430), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n437), .A2(G179), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n437), .A2(new_n438), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n415), .B1(new_n441), .B2(G169), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n414), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(G200), .B1(new_n431), .B2(new_n434), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n437), .A2(G190), .A3(new_n438), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(new_n445), .A3(new_n413), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n443), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n344), .A2(G232), .A3(new_n297), .A4(new_n346), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT75), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT75), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n428), .A2(new_n450), .A3(G232), .A4(new_n346), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n342), .A2(G1698), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(G223), .B2(G1698), .ZN(new_n454));
  INV_X1    g0254(.A(G87), .ZN(new_n455));
  OAI22_X1  g0255(.A1(new_n454), .A2(new_n332), .B1(new_n250), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n432), .B1(new_n456), .B2(new_n279), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n452), .A2(new_n457), .A3(new_n313), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n452), .A2(new_n457), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n458), .B1(new_n459), .B2(G200), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT74), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n275), .A2(new_n209), .A3(new_n276), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT7), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n275), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n276), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n403), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n372), .A2(new_n403), .ZN(new_n467));
  OAI21_X1  g0267(.A(G20), .B1(new_n467), .B2(new_n201), .ZN(new_n468));
  INV_X1    g0268(.A(G159), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(new_n326), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n461), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT16), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT16), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n461), .B(new_n473), .C1(new_n466), .C2(new_n470), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n261), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n323), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n318), .ZN(new_n477));
  OAI22_X1  g0277(.A1(new_n477), .A2(new_n317), .B1(new_n259), .B2(new_n476), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n460), .A2(new_n475), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT17), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n475), .A2(new_n479), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT18), .ZN(new_n484));
  AOI21_X1  g0284(.A(G169), .B1(new_n452), .B2(new_n457), .ZN(new_n485));
  INV_X1    g0285(.A(G179), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n485), .B1(new_n486), .B2(new_n459), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n483), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n262), .B1(new_n471), .B2(KEYINPUT16), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n478), .B1(new_n489), .B2(new_n474), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n452), .A2(new_n457), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n308), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(G179), .B2(new_n491), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT18), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n490), .A2(KEYINPUT17), .A3(new_n460), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n482), .A2(new_n488), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n401), .A2(new_n447), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT79), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT6), .ZN(new_n499));
  AND2_X1   g0299(.A1(G97), .A2(G107), .ZN(new_n500));
  NOR2_X1   g0300(.A1(G97), .A2(G107), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(KEYINPUT6), .A2(G97), .ZN(new_n503));
  OAI21_X1  g0303(.A(KEYINPUT76), .B1(new_n503), .B2(G107), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT76), .ZN(new_n505));
  INV_X1    g0305(.A(G107), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT6), .A4(G97), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n502), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n508), .A2(G20), .B1(G77), .B2(new_n406), .ZN(new_n509));
  AOI21_X1  g0309(.A(KEYINPUT7), .B1(new_n332), .B2(new_n209), .ZN(new_n510));
  INV_X1    g0310(.A(new_n465), .ZN(new_n511));
  OAI21_X1  g0311(.A(G107), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n262), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n259), .A2(G97), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(new_n264), .B2(G97), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n498), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n508), .A2(G20), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n406), .A2(G77), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n506), .B1(new_n464), .B2(new_n465), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n261), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n522), .A2(KEYINPUT79), .A3(new_n515), .ZN(new_n523));
  NAND2_X1  g0323(.A1(G33), .A2(G283), .ZN(new_n524));
  OAI211_X1 g0324(.A(G250), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n525));
  OAI211_X1 g0325(.A(G244), .B(new_n272), .C1(new_n269), .C2(new_n270), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT4), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n524), .B(new_n525), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT4), .B1(new_n331), .B2(G244), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n279), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n296), .A2(G257), .A3(new_n297), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT78), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT78), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n296), .A2(new_n533), .A3(G257), .A4(new_n297), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n530), .A2(new_n535), .A3(new_n295), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G169), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n284), .A2(new_n289), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n294), .A2(new_n290), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n532), .A2(new_n534), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n541), .A2(G179), .A3(new_n530), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n517), .A2(new_n523), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n297), .B1(G250), .B2(new_n286), .ZN(new_n544));
  NOR3_X1   g0344(.A1(new_n285), .A2(G1), .A3(G274), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  OAI211_X1 g0347(.A(G238), .B(new_n272), .C1(new_n269), .C2(new_n270), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n250), .A2(new_n247), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT80), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n334), .A2(new_n552), .A3(G244), .A4(G1698), .ZN(new_n553));
  OAI211_X1 g0353(.A(G244), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT80), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n551), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n547), .B1(new_n556), .B2(new_n297), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G200), .ZN(new_n558));
  OAI211_X1 g0358(.A(G190), .B(new_n547), .C1(new_n556), .C2(new_n297), .ZN(new_n559));
  NAND3_X1  g0359(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT81), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n560), .A2(new_n561), .A3(new_n209), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n561), .B1(new_n560), .B2(new_n209), .ZN(new_n563));
  NOR3_X1   g0363(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n564));
  NOR3_X1   g0364(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n209), .B(G68), .C1(new_n269), .C2(new_n270), .ZN(new_n566));
  INV_X1    g0366(.A(G97), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n324), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n566), .B1(KEYINPUT19), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n261), .B1(new_n565), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n381), .A2(new_n402), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n264), .A2(G87), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n558), .A2(new_n559), .A3(new_n573), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n486), .B(new_n547), .C1(new_n556), .C2(new_n297), .ZN(new_n575));
  INV_X1    g0375(.A(new_n381), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n264), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n570), .A2(new_n577), .A3(new_n571), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n555), .A2(new_n553), .ZN(new_n579));
  INV_X1    g0379(.A(new_n551), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n546), .B1(new_n581), .B2(new_n279), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n575), .B(new_n578), .C1(new_n582), .C2(G169), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n574), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n536), .A2(G200), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n513), .A2(new_n516), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n541), .A2(G190), .A3(new_n530), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n543), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n209), .B(G87), .C1(new_n269), .C2(new_n270), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT22), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT22), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n334), .A2(new_n592), .A3(new_n209), .A4(G87), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT24), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT23), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n209), .B2(G107), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n506), .A2(KEYINPUT23), .A3(G20), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n597), .A2(new_n598), .B1(new_n549), .B2(new_n209), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n594), .A2(new_n595), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n595), .B1(new_n594), .B2(new_n599), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n261), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT84), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT25), .ZN(new_n604));
  AOI211_X1 g0404(.A(G107), .B(new_n259), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  OR2_X1    g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n606), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n607), .A2(new_n608), .B1(G107), .B2(new_n264), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n331), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n610));
  OAI211_X1 g0410(.A(G257), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n297), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n287), .A2(G41), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n297), .B(G264), .C1(new_n282), .C2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n295), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(G169), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT85), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n296), .A2(KEYINPUT85), .A3(G264), .A4(new_n297), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(G250), .B(new_n272), .C1(new_n269), .C2(new_n270), .ZN(new_n621));
  INV_X1    g0421(.A(G294), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n611), .B(new_n621), .C1(new_n250), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n279), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n620), .A2(new_n624), .A3(G179), .A4(new_n295), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n602), .A2(new_n609), .B1(new_n616), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT86), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n602), .A2(new_n609), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n612), .A2(new_n615), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n620), .A2(new_n624), .A3(new_n295), .ZN(new_n630));
  INV_X1    g0430(.A(G200), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n313), .A2(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n627), .B1(new_n628), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n630), .A2(new_n631), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n624), .A2(new_n313), .A3(new_n295), .A4(new_n614), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n636), .A2(KEYINPUT86), .A3(new_n602), .A4(new_n609), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n626), .B1(new_n633), .B2(new_n637), .ZN(new_n638));
  AND4_X1   g0438(.A1(new_n316), .A2(new_n497), .A3(new_n589), .A4(new_n638), .ZN(G372));
  INV_X1    g0439(.A(new_n583), .ZN(new_n640));
  INV_X1    g0440(.A(new_n584), .ZN(new_n641));
  XNOR2_X1  g0441(.A(KEYINPUT87), .B(KEYINPUT26), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n641), .A2(new_n543), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n586), .B1(new_n537), .B2(new_n542), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n645), .B1(new_n647), .B2(new_n584), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n640), .B1(new_n644), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n633), .A2(new_n637), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n543), .A2(new_n588), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n616), .A2(new_n625), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n594), .A2(new_n599), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(KEYINPUT24), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n594), .A2(new_n595), .A3(new_n599), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n262), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n607), .A2(new_n608), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n264), .A2(G107), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n652), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n304), .A2(new_n660), .A3(new_n307), .A4(new_n310), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n650), .A2(new_n651), .A3(new_n661), .A4(new_n641), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n649), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n497), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n482), .A2(new_n495), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n446), .A2(new_n399), .A3(new_n396), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n665), .B1(new_n443), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n488), .A2(new_n494), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n355), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n669), .A2(new_n361), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n664), .A2(new_n670), .ZN(G369));
  NAND3_X1  g0471(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(G343), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n266), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n311), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n316), .A2(new_n678), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT88), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n628), .A2(new_n677), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n638), .A2(new_n687), .B1(new_n626), .B2(new_n677), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n311), .A2(new_n676), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n638), .ZN(new_n693));
  XOR2_X1   g0493(.A(new_n676), .B(KEYINPUT89), .Z(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n693), .B1(new_n660), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n690), .A2(new_n697), .ZN(G399));
  NAND3_X1  g0498(.A1(new_n212), .A2(KEYINPUT90), .A3(new_n281), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(KEYINPUT90), .B1(new_n212), .B2(new_n281), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n564), .A2(new_n247), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n703), .A2(G1), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n215), .B2(new_n703), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n695), .B1(new_n649), .B2(new_n662), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n709), .A2(KEYINPUT29), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT91), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n583), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n523), .A2(new_n517), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n537), .A2(new_n542), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n642), .B1(new_n715), .B2(new_n584), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n646), .A2(KEYINPUT26), .A3(new_n583), .A4(new_n574), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n712), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n662), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n719), .A2(KEYINPUT29), .A3(new_n676), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n710), .A2(new_n720), .ZN(new_n721));
  AND4_X1   g0521(.A1(new_n316), .A2(new_n589), .A3(new_n638), .A4(new_n694), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n306), .A2(new_n582), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n618), .A2(new_n619), .B1(new_n623), .B2(new_n279), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n724), .A2(new_n541), .A3(new_n530), .ZN(new_n725));
  OAI21_X1  g0525(.A(KEYINPUT30), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n725), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n557), .A2(new_n305), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT30), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  AND4_X1   g0531(.A1(new_n486), .A2(new_n536), .A3(new_n557), .A4(new_n630), .ZN(new_n732));
  INV_X1    g0532(.A(new_n303), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n695), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT31), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n726), .A2(new_n730), .B1(new_n732), .B2(new_n733), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n737), .B1(new_n738), .B2(new_n676), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n736), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(G330), .B1(new_n722), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n721), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n708), .B1(new_n743), .B2(G1), .ZN(G364));
  INV_X1    g0544(.A(new_n686), .ZN(new_n745));
  INV_X1    g0545(.A(G13), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G20), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n208), .B1(new_n747), .B2(G45), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n702), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n745), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(G330), .B2(new_n685), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n212), .A2(new_n334), .ZN(new_n753));
  INV_X1    g0553(.A(G355), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n753), .A2(new_n754), .B1(G116), .B2(new_n212), .ZN(new_n755));
  INV_X1    g0555(.A(new_n212), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n334), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n758), .B1(new_n285), .B2(new_n216), .ZN(new_n759));
  OR2_X1    g0559(.A1(new_n240), .A2(new_n285), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n755), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G13), .A2(G33), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n217), .B1(G20), .B2(new_n308), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n750), .B1(new_n761), .B2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n765), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n209), .A2(new_n486), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G190), .A2(G200), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n334), .B1(new_n772), .B2(new_n205), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n209), .A2(G179), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(G190), .A3(G200), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n774), .A2(new_n313), .A3(G200), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n455), .A2(new_n775), .B1(new_n776), .B2(new_n506), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n770), .A2(G190), .A3(new_n631), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n773), .B(new_n777), .C1(G58), .C2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n770), .A2(G190), .A3(G200), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT92), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G50), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n313), .A2(G179), .A3(G200), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n209), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n567), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n770), .A2(new_n313), .A3(G200), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n790), .B1(G68), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n774), .A2(new_n771), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n469), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT32), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n780), .A2(new_n787), .A3(new_n793), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n786), .A2(G326), .ZN(new_n798));
  INV_X1    g0598(.A(G303), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n332), .B1(new_n775), .B2(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT93), .ZN(new_n801));
  INV_X1    g0601(.A(G322), .ZN(new_n802));
  INV_X1    g0602(.A(G311), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n778), .A2(new_n802), .B1(new_n772), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n794), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n804), .B1(G329), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G283), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n789), .A2(new_n622), .B1(new_n776), .B2(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(KEYINPUT33), .B(G317), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n808), .B1(new_n792), .B2(new_n809), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n798), .A2(new_n801), .A3(new_n806), .A4(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n769), .B1(new_n797), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n768), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n764), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n683), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n752), .A2(new_n815), .ZN(G396));
  AOI21_X1  g0616(.A(G169), .B1(new_n386), .B2(new_n387), .ZN(new_n817));
  OAI21_X1  g0617(.A(KEYINPUT71), .B1(new_n385), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n391), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n385), .A2(new_n676), .ZN(new_n820));
  AND4_X1   g0620(.A1(new_n399), .A2(new_n818), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n820), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n821), .B1(new_n400), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n709), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n709), .A2(new_n824), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n742), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT96), .ZN(new_n829));
  INV_X1    g0629(.A(new_n750), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n829), .B(new_n830), .C1(new_n742), .C2(new_n827), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n765), .A2(new_n762), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n750), .B1(G77), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(new_n834), .B(KEYINPUT94), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n786), .A2(G303), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n332), .B1(new_n775), .B2(new_n506), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT95), .Z(new_n838));
  NOR2_X1   g0638(.A1(new_n776), .A2(new_n455), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n839), .B(new_n790), .C1(G283), .C2(new_n792), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n778), .A2(new_n622), .B1(new_n772), .B2(new_n247), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(G311), .B2(new_n805), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n836), .A2(new_n838), .A3(new_n840), .A4(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(G132), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n334), .B1(new_n794), .B2(new_n844), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n202), .A2(new_n775), .B1(new_n776), .B2(new_n403), .ZN(new_n846));
  INV_X1    g0646(.A(new_n789), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n845), .B(new_n846), .C1(G58), .C2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n772), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n779), .A2(G143), .B1(new_n849), .B2(G159), .ZN(new_n850));
  INV_X1    g0650(.A(G137), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n850), .B1(new_n325), .B2(new_n791), .C1(new_n785), .C2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n848), .B1(new_n853), .B2(KEYINPUT34), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT34), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n843), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n835), .B1(new_n857), .B2(new_n765), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n824), .B2(new_n763), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n831), .A2(new_n859), .ZN(G384));
  NOR2_X1   g0660(.A1(new_n747), .A2(new_n208), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT98), .ZN(new_n863));
  INV_X1    g0663(.A(new_n675), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n490), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n496), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n480), .B1(new_n490), .B2(new_n493), .ZN(new_n867));
  OAI21_X1  g0667(.A(KEYINPUT37), .B1(new_n867), .B2(new_n865), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n483), .A2(new_n487), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n483), .A2(new_n675), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n869), .A2(new_n870), .A3(new_n871), .A4(new_n480), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n866), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n863), .B1(new_n496), .B2(new_n865), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n862), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n496), .A2(new_n865), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(KEYINPUT98), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n878), .A2(KEYINPUT38), .A3(new_n873), .A4(new_n866), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n876), .A2(KEYINPUT39), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(G169), .B1(new_n431), .B2(new_n434), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT14), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(new_n439), .A3(new_n435), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(new_n414), .A3(new_n676), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n873), .A2(new_n877), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n862), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT39), .B1(new_n879), .B2(new_n886), .ZN(new_n887));
  OR3_X1    g0687(.A1(new_n880), .A2(new_n884), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n396), .A2(new_n399), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n889), .A2(new_n677), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(new_n709), .B2(new_n824), .ZN(new_n891));
  INV_X1    g0691(.A(new_n446), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n883), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n414), .A2(new_n677), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n443), .A2(new_n446), .A3(new_n894), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT97), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n443), .A2(KEYINPUT97), .A3(new_n446), .A4(new_n894), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n895), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n891), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n876), .A2(new_n879), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n901), .A2(new_n902), .B1(new_n668), .B2(new_n864), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n888), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n497), .A2(new_n710), .A3(new_n720), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n905), .A2(new_n670), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n904), .B(new_n906), .Z(new_n907));
  INV_X1    g0707(.A(G330), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT40), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n876), .A2(new_n879), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n898), .A2(new_n899), .ZN(new_n911));
  INV_X1    g0711(.A(new_n895), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n914), .A2(new_n739), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n316), .A2(new_n589), .A3(new_n638), .A4(new_n694), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n823), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n909), .B1(new_n910), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n879), .A2(new_n886), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(KEYINPUT99), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n914), .A2(new_n739), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n824), .B1(new_n722), .B2(new_n922), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n900), .A2(new_n923), .A3(new_n909), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT99), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n879), .A2(new_n925), .A3(new_n886), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n921), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n919), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n915), .A2(new_n916), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n497), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n908), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n928), .B2(new_n930), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n861), .B1(new_n907), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n907), .B2(new_n932), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n508), .A2(KEYINPUT35), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n508), .A2(KEYINPUT35), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n935), .A2(G116), .A3(new_n218), .A4(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT36), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n467), .A2(new_n215), .A3(new_n205), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n403), .A2(G50), .ZN(new_n940));
  OAI211_X1 g0740(.A(G1), .B(new_n746), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n934), .A2(new_n938), .A3(new_n941), .ZN(G367));
  INV_X1    g0742(.A(new_n776), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n847), .A2(G107), .B1(new_n943), .B2(G97), .ZN(new_n944));
  OAI221_X1 g0744(.A(new_n944), .B1(new_n622), .B2(new_n791), .C1(new_n785), .C2(new_n803), .ZN(new_n945));
  AOI22_X1  g0745(.A1(G283), .A2(new_n849), .B1(new_n805), .B2(G317), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n334), .B1(new_n779), .B2(G303), .ZN(new_n947));
  INV_X1    g0747(.A(new_n775), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(KEYINPUT46), .A3(G116), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT46), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(new_n775), .B2(new_n247), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n946), .A2(new_n947), .A3(new_n949), .A4(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n789), .A2(new_n403), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(G58), .B2(new_n948), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n332), .B1(new_n779), .B2(G150), .ZN(new_n955));
  AOI22_X1  g0755(.A1(G50), .A2(new_n849), .B1(new_n805), .B2(G137), .ZN(new_n956));
  AOI22_X1  g0756(.A1(G159), .A2(new_n792), .B1(new_n943), .B2(G77), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n954), .A2(new_n955), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(G143), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n785), .A2(new_n959), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n945), .A2(new_n952), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT105), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT47), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n765), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n573), .A2(new_n676), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n641), .A2(new_n965), .ZN(new_n966));
  OR2_X1    g0766(.A1(new_n965), .A2(new_n583), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n966), .A2(new_n764), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n757), .A2(new_n236), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n767), .B1(new_n756), .B2(new_n576), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n830), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n964), .A2(new_n968), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n651), .B1(new_n586), .B2(new_n694), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n695), .A2(new_n646), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n715), .B1(new_n975), .B2(new_n660), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n694), .ZN(new_n977));
  OAI21_X1  g0777(.A(KEYINPUT42), .B1(new_n975), .B2(new_n693), .ZN(new_n978));
  OR3_X1    g0778(.A1(new_n975), .A2(new_n693), .A3(KEYINPUT42), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT100), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n966), .A2(new_n967), .ZN(new_n982));
  OR3_X1    g0782(.A1(new_n981), .A2(KEYINPUT43), .A3(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n982), .B(KEYINPUT43), .Z(new_n984));
  NAND2_X1  g0784(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT101), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n981), .A2(KEYINPUT101), .A3(new_n984), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n983), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n975), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n689), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n989), .B(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(KEYINPUT104), .B1(new_n697), .B2(new_n990), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT104), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n696), .A2(new_n994), .A3(new_n975), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT44), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n696), .A2(new_n975), .ZN(new_n999));
  XNOR2_X1  g0799(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n993), .A2(KEYINPUT44), .A3(new_n995), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n998), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(new_n689), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n690), .A2(new_n998), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n688), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n693), .B1(new_n1006), .B2(new_n692), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n745), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1007), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n686), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1004), .A2(new_n1005), .A3(new_n743), .A4(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n743), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n702), .B(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n749), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n972), .B1(new_n992), .B2(new_n1016), .ZN(G387));
  NAND2_X1  g0817(.A1(new_n1011), .A2(new_n743), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1008), .B(new_n1010), .C1(new_n742), .C2(new_n721), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n702), .B(KEYINPUT110), .Z(new_n1020));
  NAND3_X1  g0820(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  AOI211_X1 g0821(.A(G45), .B(new_n704), .C1(G68), .C2(G77), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n1023), .A2(KEYINPUT106), .ZN(new_n1024));
  OAI21_X1  g0824(.A(KEYINPUT50), .B1(new_n323), .B2(G50), .ZN(new_n1025));
  OR3_X1    g0825(.A1(new_n323), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT106), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1025), .B(new_n1026), .C1(new_n1022), .C2(new_n1027), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n757), .B1(new_n1024), .B2(new_n1028), .C1(new_n233), .C2(new_n285), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(G107), .B2(new_n212), .C1(new_n705), .C2(new_n753), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n830), .B1(new_n1030), .B2(new_n766), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(new_n1006), .B2(new_n814), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n334), .B1(new_n794), .B2(new_n325), .C1(new_n403), .C2(new_n772), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n205), .A2(new_n775), .B1(new_n776), .B2(new_n567), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1033), .B(new_n1034), .C1(new_n476), .C2(new_n792), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n789), .A2(new_n381), .B1(new_n778), .B2(new_n202), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT107), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1035), .B(new_n1037), .C1(new_n469), .C2(new_n785), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT108), .Z(new_n1039));
  AOI22_X1  g0839(.A1(new_n786), .A2(G322), .B1(G311), .B2(new_n792), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1040), .A2(KEYINPUT109), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(KEYINPUT109), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n779), .A2(G317), .B1(new_n849), .B2(G303), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1041), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT48), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n789), .A2(new_n807), .B1(new_n775), .B2(new_n622), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1046), .A2(KEYINPUT49), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n334), .B1(new_n805), .B2(G326), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(new_n247), .C2(new_n776), .ZN(new_n1051));
  AOI21_X1  g0851(.A(KEYINPUT49), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1039), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1032), .B1(new_n1053), .B2(new_n765), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(new_n1011), .B2(new_n749), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1021), .A2(new_n1055), .ZN(G393));
  INV_X1    g0856(.A(KEYINPUT111), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1057), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n1005), .A2(new_n1057), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n975), .A2(new_n764), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n766), .B1(new_n567), .B2(new_n212), .C1(new_n758), .C2(new_n243), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n750), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n785), .A2(new_n325), .B1(new_n469), .B2(new_n778), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT113), .ZN(new_n1065));
  XOR2_X1   g0865(.A(KEYINPUT112), .B(KEYINPUT51), .Z(new_n1066));
  XOR2_X1   g0866(.A(new_n1065), .B(new_n1066), .Z(new_n1067));
  OAI221_X1 g0867(.A(new_n334), .B1(new_n794), .B2(new_n959), .C1(new_n323), .C2(new_n772), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n839), .B1(G50), .B2(new_n792), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n847), .A2(G77), .B1(new_n948), .B2(G68), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n786), .A2(G317), .B1(G311), .B2(new_n779), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT52), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n332), .B1(new_n794), .B2(new_n802), .C1(new_n622), .C2(new_n772), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n791), .A2(new_n799), .B1(new_n776), .B2(new_n506), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n789), .A2(new_n247), .B1(new_n775), .B2(new_n807), .ZN(new_n1077));
  OR3_X1    g0877(.A1(new_n1075), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n1067), .A2(new_n1072), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1063), .B1(new_n1079), .B2(new_n765), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1060), .A2(new_n749), .B1(new_n1061), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1018), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1082), .A2(new_n1012), .A3(new_n1020), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1083), .ZN(G390));
  INV_X1    g0884(.A(KEYINPUT114), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n677), .B(new_n823), .C1(new_n718), .C2(new_n662), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1085), .B1(new_n1086), .B2(new_n890), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n719), .A2(new_n676), .A3(new_n824), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n890), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1088), .A2(KEYINPUT114), .A3(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1087), .A2(new_n913), .A3(new_n1090), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1091), .A2(new_n884), .A3(new_n921), .A4(new_n926), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n884), .B1(new_n891), .B2(new_n900), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n880), .B2(new_n887), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n900), .A2(new_n741), .A3(new_n823), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n1092), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT115), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n913), .A2(new_n1098), .A3(G330), .A4(new_n917), .ZN(new_n1099));
  OAI211_X1 g0899(.A(G330), .B(new_n824), .C1(new_n722), .C2(new_n922), .ZN(new_n1100));
  OAI21_X1  g0900(.A(KEYINPUT115), .B1(new_n900), .B2(new_n1100), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n900), .B1(new_n741), .B2(new_n823), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1099), .A2(new_n1101), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n891), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n900), .A2(new_n1100), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1095), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1105), .A2(new_n1106), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n497), .A2(G330), .A3(new_n929), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n905), .A2(new_n1111), .A3(new_n670), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n1097), .A2(new_n1103), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1112), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1102), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1092), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1116), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1113), .A2(new_n1121), .A3(new_n1020), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1097), .A2(new_n1103), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n762), .B1(new_n880), .B2(new_n887), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(G137), .A2(new_n792), .B1(new_n943), .B2(G50), .ZN(new_n1125));
  INV_X1    g0925(.A(G128), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1125), .B1(new_n469), .B2(new_n789), .C1(new_n785), .C2(new_n1126), .ZN(new_n1127));
  XOR2_X1   g0927(.A(KEYINPUT54), .B(G143), .Z(new_n1128));
  AOI22_X1  g0928(.A1(new_n849), .A2(new_n1128), .B1(new_n805), .B2(G125), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n332), .B1(new_n779), .B2(G132), .ZN(new_n1130));
  OR3_X1    g0930(.A1(new_n775), .A2(KEYINPUT53), .A3(new_n325), .ZN(new_n1131));
  OAI21_X1  g0931(.A(KEYINPUT53), .B1(new_n775), .B2(new_n325), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n785), .A2(new_n807), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(G77), .A2(new_n847), .B1(new_n792), .B2(G107), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n948), .A2(G87), .B1(new_n943), .B2(G68), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n334), .B1(new_n779), .B2(G116), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(G97), .A2(new_n849), .B1(new_n805), .B2(G294), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n1127), .A2(new_n1133), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT117), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n769), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n1141), .B2(new_n1140), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n750), .B1(new_n476), .B2(new_n833), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT116), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1123), .A2(new_n749), .B1(new_n1124), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1122), .A2(new_n1147), .ZN(G378));
  OR2_X1    g0948(.A1(new_n904), .A2(KEYINPUT121), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n904), .A2(KEYINPUT121), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n355), .A2(new_n361), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n329), .A2(new_n675), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1151), .B(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n919), .A2(new_n927), .A3(G330), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(KEYINPUT119), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n900), .A2(new_n923), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n902), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n908), .B1(new_n1159), .B2(new_n909), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT119), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n1161), .A3(new_n927), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1155), .B1(new_n1157), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1161), .B1(new_n1160), .B2(new_n927), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1155), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1149), .B(new_n1150), .C1(new_n1163), .C2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT57), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1112), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1168), .B1(new_n1121), .B2(new_n1169), .ZN(new_n1170));
  AND4_X1   g0970(.A1(new_n1161), .A2(new_n919), .A3(G330), .A4(new_n927), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1165), .B1(new_n1171), .B2(new_n1164), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1157), .A2(new_n1155), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1172), .A2(KEYINPUT121), .A3(new_n904), .A4(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1167), .A2(new_n1170), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1110), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1112), .B1(new_n1123), .B2(new_n1176), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n904), .A2(KEYINPUT120), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1178), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n904), .A2(KEYINPUT120), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1172), .A2(new_n1173), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1177), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1020), .B(new_n1175), .C1(new_n1182), .C2(KEYINPUT57), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n776), .A2(new_n372), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT118), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G116), .B2(new_n786), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n332), .A2(new_n281), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n772), .A2(new_n381), .B1(new_n794), .B2(new_n807), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1187), .B(new_n1188), .C1(G107), .C2(new_n779), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n775), .A2(new_n205), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1190), .B(new_n953), .C1(G97), .C2(new_n792), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1186), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT58), .ZN(new_n1193));
  AOI21_X1  g0993(.A(G50), .B1(new_n250), .B2(new_n281), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1192), .A2(new_n1193), .B1(new_n1187), .B2(new_n1194), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n778), .A2(new_n1126), .B1(new_n772), .B2(new_n851), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1196), .B1(G132), .B2(new_n792), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n847), .A2(G150), .B1(new_n948), .B2(new_n1128), .ZN(new_n1198));
  INV_X1    g0998(.A(G125), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1197), .B(new_n1198), .C1(new_n1199), .C2(new_n785), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n943), .A2(G159), .ZN(new_n1203));
  AOI211_X1 g1003(.A(G33), .B(G41), .C1(new_n805), .C2(G124), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1195), .B1(new_n1193), .B2(new_n1192), .C1(new_n1201), .C2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n765), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n830), .B1(new_n202), .B2(new_n832), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1207), .B(new_n1208), .C1(new_n1155), .C2(new_n763), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1210), .B1(new_n1211), .B2(new_n749), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1183), .A2(new_n1212), .ZN(G375));
  INV_X1    g1013(.A(new_n1116), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1214), .A2(new_n1215), .A3(new_n1015), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT122), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n334), .B1(new_n805), .B2(G303), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n506), .B2(new_n772), .C1(new_n807), .C2(new_n778), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(G116), .A2(new_n792), .B1(new_n948), .B2(G97), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1220), .B1(new_n205), .B2(new_n776), .C1(new_n381), .C2(new_n789), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n1219), .B(new_n1221), .C1(G294), .C2(new_n786), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G50), .A2(new_n847), .B1(new_n792), .B2(new_n1128), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n332), .B1(new_n849), .B2(G150), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1223), .B(new_n1224), .C1(new_n851), .C2(new_n778), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1185), .B(new_n1225), .C1(G132), .C2(new_n786), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n775), .A2(new_n469), .B1(new_n794), .B2(new_n1126), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT123), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1222), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1229));
  OAI221_X1 g1029(.A(new_n750), .B1(G68), .B2(new_n833), .C1(new_n1229), .C2(new_n769), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n900), .B2(new_n762), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1176), .B2(new_n749), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1217), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1233), .ZN(G381));
  NAND4_X1  g1034(.A1(new_n1021), .A2(new_n815), .A3(new_n752), .A4(new_n1055), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(G384), .A2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1081), .A2(new_n1083), .A3(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(G387), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n1233), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT124), .ZN(new_n1240));
  INV_X1    g1040(.A(G378), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1183), .A2(new_n1241), .A3(new_n1212), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1240), .A2(new_n1243), .ZN(G407));
  INV_X1    g1044(.A(G343), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(G213), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1242), .A2(new_n1246), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT125), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(G407), .A2(G213), .A3(new_n1248), .ZN(G409));
  NAND2_X1  g1049(.A1(G393), .A2(G396), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n1235), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n1083), .B2(new_n1081), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  XOR2_X1   g1053(.A(new_n989), .B(new_n991), .Z(new_n1254));
  INV_X1    g1054(.A(new_n1016), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1081), .A2(new_n1083), .A3(new_n1251), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1253), .A2(new_n972), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1257), .ZN(new_n1259));
  OAI21_X1  g1059(.A(G387), .B1(new_n1259), .B2(new_n1252), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1258), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT61), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT60), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1215), .A2(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1110), .A2(KEYINPUT60), .A3(new_n1112), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1264), .A2(new_n1020), .A3(new_n1214), .A4(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(G384), .B1(new_n1266), .B2(new_n1232), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1266), .A2(G384), .A3(new_n1232), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1245), .A2(G213), .A3(G2897), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1268), .A2(new_n1269), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1269), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1270), .B1(new_n1273), .B2(new_n1267), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1241), .B1(new_n1183), .B2(new_n1212), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1121), .A2(new_n1169), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(new_n1163), .A2(new_n1178), .A3(new_n1166), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1180), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1015), .B(new_n1277), .C1(new_n1278), .C2(new_n1279), .ZN(new_n1280));
  AND3_X1   g1080(.A1(new_n1122), .A2(new_n1147), .A3(new_n1209), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1167), .A2(new_n749), .A3(new_n1174), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1280), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1246), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1275), .B1(new_n1276), .B2(new_n1284), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1273), .A2(new_n1267), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1276), .A2(new_n1284), .A3(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT62), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1262), .B(new_n1285), .C1(new_n1288), .C2(new_n1289), .ZN(new_n1290));
  NOR4_X1   g1090(.A1(new_n1276), .A2(new_n1284), .A3(new_n1287), .A4(KEYINPUT62), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1261), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT63), .ZN(new_n1293));
  OR2_X1    g1093(.A1(new_n1276), .A2(new_n1284), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1293), .B1(new_n1294), .B2(new_n1287), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1261), .A2(KEYINPUT61), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1288), .A2(KEYINPUT63), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1275), .A2(KEYINPUT126), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT126), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1272), .A2(new_n1274), .A3(new_n1299), .ZN(new_n1300));
  OAI211_X1 g1100(.A(new_n1298), .B(new_n1300), .C1(new_n1276), .C2(new_n1284), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1295), .A2(new_n1296), .A3(new_n1297), .A4(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1292), .A2(new_n1302), .ZN(G405));
  OAI21_X1  g1103(.A(new_n1287), .B1(new_n1243), .B2(new_n1276), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1276), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1305), .A2(new_n1242), .A3(new_n1286), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1258), .A2(KEYINPUT127), .A3(new_n1260), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1304), .A2(new_n1306), .A3(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT127), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1308), .A2(new_n1309), .A3(new_n1261), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1261), .A2(new_n1309), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1311), .A2(new_n1304), .A3(new_n1307), .A4(new_n1306), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1310), .A2(new_n1312), .ZN(G402));
endmodule


