//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n813, new_n814,
    new_n815, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n864, new_n865, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915;
  INV_X1    g000(.A(KEYINPUT86), .ZN(new_n202));
  INV_X1    g001(.A(G141gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n203), .A2(KEYINPUT77), .A3(G148gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT77), .ZN(new_n205));
  INV_X1    g004(.A(G148gat), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n205), .B1(G141gat), .B2(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(G141gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n204), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT78), .ZN(new_n210));
  XNOR2_X1  g009(.A(G155gat), .B(G162gat), .ZN(new_n211));
  INV_X1    g010(.A(G155gat), .ZN(new_n212));
  INV_X1    g011(.A(G162gat), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT2), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT78), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n215), .B(new_n204), .C1(new_n207), .C2(new_n208), .ZN(new_n216));
  NAND4_X1  g015(.A1(new_n210), .A2(new_n211), .A3(new_n214), .A4(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n218));
  XNOR2_X1  g017(.A(G141gat), .B(G148gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(KEYINPUT2), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n220), .A2(new_n211), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n217), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT79), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT79), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n217), .A2(new_n224), .A3(new_n218), .A4(new_n221), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT29), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G211gat), .ZN(new_n229));
  INV_X1    g028(.A(G218gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G211gat), .A2(G218gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT74), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n231), .A2(KEYINPUT74), .A3(new_n232), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  XOR2_X1   g036(.A(G197gat), .B(G204gat), .Z(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n229), .A2(KEYINPUT72), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT72), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G211gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(new_n242), .A3(G218gat), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT22), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n243), .A2(KEYINPUT73), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT73), .B1(new_n243), .B2(new_n244), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n237), .B(new_n239), .C1(new_n245), .C2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT75), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n243), .A2(new_n244), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT73), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n243), .A2(KEYINPUT73), .A3(new_n244), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT75), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n253), .A2(new_n254), .A3(new_n237), .A4(new_n239), .ZN(new_n255));
  INV_X1    g054(.A(new_n237), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n239), .B1(new_n245), .B2(new_n246), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n248), .A2(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n202), .B1(new_n228), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT29), .B1(new_n223), .B2(new_n225), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n238), .B1(new_n251), .B2(new_n252), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n254), .B1(new_n261), .B2(new_n237), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n247), .A2(KEYINPUT75), .ZN(new_n263));
  OAI22_X1  g062(.A1(new_n262), .A2(new_n263), .B1(new_n237), .B2(new_n261), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n260), .A2(new_n264), .A3(KEYINPUT86), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(KEYINPUT85), .A3(new_n227), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT85), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n268), .B1(new_n258), .B2(KEYINPUT29), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n269), .A3(new_n218), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n217), .A2(new_n221), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G228gat), .ZN(new_n273));
  INV_X1    g072(.A(G233gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n266), .A2(new_n272), .A3(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT84), .B1(new_n261), .B2(new_n237), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT84), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n257), .A2(new_n278), .A3(new_n256), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n277), .B(new_n279), .C1(new_n262), .C2(new_n263), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT3), .B1(new_n280), .B2(new_n227), .ZN(new_n281));
  INV_X1    g080(.A(new_n271), .ZN(new_n282));
  OAI22_X1  g081(.A1(new_n281), .A2(new_n282), .B1(new_n264), .B2(new_n260), .ZN(new_n283));
  INV_X1    g082(.A(new_n275), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n276), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT87), .ZN(new_n287));
  INV_X1    g086(.A(G22gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  XOR2_X1   g088(.A(G78gat), .B(G106gat), .Z(new_n290));
  XNOR2_X1  g089(.A(new_n290), .B(G50gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT83), .ZN(new_n292));
  XOR2_X1   g091(.A(new_n292), .B(KEYINPUT31), .Z(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(KEYINPUT87), .A2(G22gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n287), .A2(new_n288), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n276), .A2(new_n285), .A3(new_n295), .A4(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n289), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n288), .A2(KEYINPUT88), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n284), .B1(new_n270), .B2(new_n271), .ZN(new_n300));
  AOI221_X4 g099(.A(new_n299), .B1(new_n283), .B2(new_n284), .C1(new_n300), .C2(new_n266), .ZN(new_n301));
  INV_X1    g100(.A(new_n299), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n302), .B1(new_n276), .B2(new_n285), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT89), .B1(new_n304), .B2(new_n293), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT89), .ZN(new_n306));
  NOR4_X1   g105(.A1(new_n301), .A2(new_n303), .A3(new_n306), .A4(new_n294), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n298), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G120gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G113gat), .ZN(new_n310));
  INV_X1    g109(.A(G113gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G120gat), .ZN(new_n312));
  AND2_X1   g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(G127gat), .B1(new_n313), .B2(KEYINPUT1), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT1), .B1(new_n310), .B2(new_n312), .ZN(new_n315));
  INV_X1    g114(.A(G127gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n314), .A2(G134gat), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G134gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n315), .A2(new_n316), .ZN(new_n320));
  AOI211_X1 g119(.A(KEYINPUT1), .B(G127gat), .C1(new_n310), .C2(new_n312), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n319), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n217), .A2(new_n221), .A3(new_n318), .A4(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT4), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n323), .B(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n271), .A2(KEYINPUT3), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n318), .A2(new_n322), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n327), .B1(new_n223), .B2(new_n225), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n325), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT5), .ZN(new_n330));
  NAND2_X1  g129(.A1(G225gat), .A2(G233gat), .ZN(new_n331));
  NAND4_X1  g130(.A1(new_n329), .A2(KEYINPUT81), .A3(new_n330), .A4(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n328), .A2(new_n326), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n323), .B(KEYINPUT4), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n333), .A2(new_n330), .A3(new_n331), .A4(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT81), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(G57gat), .B(G85gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(G1gat), .B(G29gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n341), .B(new_n342), .Z(new_n343));
  XNOR2_X1  g142(.A(new_n327), .B(new_n271), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n344), .A2(new_n331), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n333), .A2(new_n334), .ZN(new_n346));
  INV_X1    g145(.A(new_n331), .ZN(new_n347));
  OAI211_X1 g146(.A(KEYINPUT5), .B(new_n345), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n338), .A2(new_n343), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT82), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n338), .A2(new_n348), .ZN(new_n352));
  INV_X1    g151(.A(new_n343), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT6), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n338), .A2(KEYINPUT82), .A3(new_n348), .A4(new_n343), .ZN(new_n356));
  NAND4_X1  g155(.A1(new_n351), .A2(new_n354), .A3(new_n355), .A4(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n352), .A2(KEYINPUT6), .A3(new_n353), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT23), .ZN(new_n360));
  INV_X1    g159(.A(G169gat), .ZN(new_n361));
  INV_X1    g160(.A(G176gat), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n364));
  AOI22_X1  g163(.A1(new_n363), .A2(new_n364), .B1(G169gat), .B2(G176gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(G183gat), .A2(G190gat), .ZN(new_n366));
  XOR2_X1   g165(.A(new_n366), .B(KEYINPUT24), .Z(new_n367));
  NOR2_X1   g166(.A1(G183gat), .A2(G190gat), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n365), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT25), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT27), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(G183gat), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT28), .B1(new_n372), .B2(KEYINPUT66), .ZN(new_n373));
  INV_X1    g172(.A(G190gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(KEYINPUT27), .B(G183gat), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n373), .B(new_n374), .C1(KEYINPUT66), .C2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n374), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT28), .ZN(new_n378));
  OR3_X1    g177(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n379), .B(new_n380), .C1(new_n361), .C2(new_n362), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n376), .A2(new_n378), .A3(new_n366), .A4(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n365), .B1(KEYINPUT65), .B2(KEYINPUT25), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n366), .B(KEYINPUT24), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT64), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n368), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n383), .B(new_n388), .C1(KEYINPUT65), .C2(new_n365), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n327), .A2(new_n370), .A3(new_n382), .A4(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n370), .A3(new_n382), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n318), .A2(new_n322), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G227gat), .A2(G233gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G71gat), .B(G99gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(G15gat), .B(G43gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n400), .B(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n395), .B1(new_n390), .B2(new_n393), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT32), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n402), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n394), .A2(new_n396), .ZN(new_n406));
  XOR2_X1   g205(.A(KEYINPUT67), .B(KEYINPUT33), .Z(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n406), .A2(KEYINPUT68), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT68), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n410), .B1(new_n403), .B2(new_n407), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n405), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n402), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n406), .B(KEYINPUT32), .C1(new_n408), .C2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n397), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n413), .B1(new_n406), .B2(KEYINPUT32), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT68), .B1(new_n406), .B2(new_n408), .ZN(new_n418));
  NOR3_X1   g217(.A1(new_n403), .A2(new_n410), .A3(new_n407), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n397), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n421), .A3(new_n414), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT34), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n423), .B1(new_n395), .B2(KEYINPUT71), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n416), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n424), .B1(new_n416), .B2(new_n422), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n391), .A2(new_n227), .ZN(new_n429));
  NAND2_X1  g228(.A1(G226gat), .A2(G233gat), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n430), .B(KEYINPUT76), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n391), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n264), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n429), .A2(new_n432), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n391), .A2(G226gat), .A3(G233gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n436), .B1(new_n264), .B2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G8gat), .B(G36gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(G64gat), .ZN(new_n442));
  INV_X1    g241(.A(G92gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(new_n442), .B(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT30), .B1(new_n440), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n440), .A2(new_n444), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n308), .A2(new_n359), .A3(new_n428), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT35), .ZN(new_n450));
  INV_X1    g249(.A(new_n428), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n286), .A2(new_n299), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n276), .A2(new_n285), .A3(new_n302), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(new_n293), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(new_n306), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n452), .A2(KEYINPUT89), .A3(new_n453), .A4(new_n293), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n451), .B1(new_n457), .B2(new_n298), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT35), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n458), .A2(new_n459), .A3(new_n359), .A4(new_n448), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n450), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT37), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n444), .B1(new_n440), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT38), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n439), .A2(new_n264), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n465), .B(KEYINPUT37), .C1(new_n264), .C2(new_n435), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n463), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n446), .ZN(new_n468));
  OR2_X1    g267(.A1(new_n440), .A2(new_n462), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n464), .B1(new_n469), .B2(new_n463), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n357), .A2(new_n471), .A3(new_n358), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n344), .A2(new_n331), .ZN(new_n473));
  OAI211_X1 g272(.A(KEYINPUT39), .B(new_n473), .C1(new_n329), .C2(new_n331), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n346), .A2(new_n347), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n474), .B(new_n343), .C1(KEYINPUT39), .C2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT90), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT40), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n477), .B1(new_n476), .B2(new_n478), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n476), .A2(new_n478), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n481), .A2(new_n354), .A3(new_n447), .A4(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n308), .A2(new_n472), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n359), .A2(new_n448), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n485), .A2(new_n298), .A3(new_n457), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT36), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n426), .A2(new_n427), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n416), .A2(new_n422), .ZN(new_n489));
  INV_X1    g288(.A(new_n424), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT36), .B1(new_n491), .B2(new_n425), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n484), .B(new_n486), .C1(new_n488), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n461), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(G43gat), .B(G50gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(KEYINPUT15), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  OR3_X1    g296(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT93), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT94), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(G29gat), .ZN(new_n504));
  INV_X1    g303(.A(G36gat), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n497), .B(new_n498), .C1(new_n503), .C2(new_n506), .ZN(new_n507));
  XOR2_X1   g306(.A(new_n496), .B(KEYINPUT95), .Z(new_n508));
  OAI21_X1  g307(.A(new_n498), .B1(new_n501), .B2(new_n506), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n495), .A2(KEYINPUT15), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT96), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT17), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n507), .A2(KEYINPUT17), .A3(new_n512), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(G15gat), .B(G22gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT16), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n519), .B1(new_n520), .B2(G1gat), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(G1gat), .B2(new_n519), .ZN(new_n522));
  INV_X1    g321(.A(G8gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n522), .B(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n524), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n513), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G229gat), .A2(G233gat), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n525), .A2(KEYINPUT18), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n513), .B(new_n526), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n528), .B(KEYINPUT13), .Z(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n527), .B(new_n528), .C1(new_n517), .C2(new_n526), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT18), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n529), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n537));
  XNOR2_X1  g336(.A(G113gat), .B(G141gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G169gat), .B(G197gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(KEYINPUT12), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n542), .B(KEYINPUT92), .Z(new_n543));
  NAND2_X1  g342(.A1(new_n536), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT97), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n529), .A2(new_n532), .A3(new_n535), .A4(new_n542), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT97), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n536), .A2(new_n547), .A3(new_n543), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G120gat), .B(G148gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(new_n362), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(G204gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(G230gat), .A2(G233gat), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n554), .B(KEYINPUT103), .Z(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G57gat), .B(G64gat), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n558));
  OR2_X1    g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G71gat), .B(G78gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562));
  INV_X1    g361(.A(G85gat), .ZN(new_n563));
  AOI22_X1  g362(.A1(KEYINPUT8), .A2(new_n562), .B1(new_n563), .B2(new_n443), .ZN(new_n564));
  NAND2_X1  g363(.A1(G85gat), .A2(G92gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(KEYINPUT99), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT99), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n567), .A2(G85gat), .A3(G92gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT7), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n569), .B1(new_n566), .B2(new_n568), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n564), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G99gat), .B(G106gat), .Z(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n573), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n575), .B(new_n564), .C1(new_n570), .C2(new_n571), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n561), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n574), .A2(KEYINPUT100), .A3(new_n576), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n559), .B(new_n560), .Z(new_n579));
  INV_X1    g378(.A(KEYINPUT100), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n572), .A2(new_n580), .A3(new_n573), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT102), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT102), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n578), .A2(new_n579), .A3(new_n584), .A4(new_n581), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n577), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT10), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI211_X1 g387(.A(new_n587), .B(new_n579), .C1(new_n578), .C2(new_n581), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT104), .B1(new_n591), .B2(new_n556), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n589), .B1(new_n586), .B2(new_n587), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT104), .ZN(new_n594));
  NOR3_X1   g393(.A1(new_n593), .A2(new_n594), .A3(new_n555), .ZN(new_n595));
  OAI221_X1 g394(.A(new_n553), .B1(new_n556), .B2(new_n586), .C1(new_n592), .C2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n553), .B(KEYINPUT105), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n593), .A2(new_n555), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n586), .A2(new_n556), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n550), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n561), .A2(KEYINPUT21), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n526), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT21), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n604), .B1(new_n605), .B2(new_n579), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n526), .A2(new_n603), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G127gat), .B(G155gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n610), .B(new_n611), .Z(new_n612));
  XNOR2_X1  g411(.A(G183gat), .B(G211gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT20), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n612), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G190gat), .B(G218gat), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n578), .A2(new_n581), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n513), .A2(new_n620), .ZN(new_n621));
  AND2_X1   g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT41), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n621), .A2(KEYINPUT101), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT101), .B1(new_n621), .B2(new_n623), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n517), .A2(new_n620), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n622), .A2(KEYINPUT41), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n626), .B(new_n627), .C1(KEYINPUT41), .C2(new_n622), .ZN(new_n631));
  XNOR2_X1  g430(.A(G134gat), .B(G162gat), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n633), .B1(new_n630), .B2(new_n631), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n619), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n630), .A2(new_n631), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n632), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n638), .A2(new_n639), .A3(new_n618), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n636), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n617), .A2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n494), .A2(new_n602), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n359), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g446(.A1(new_n643), .A2(new_n448), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n648), .A2(new_n523), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT106), .ZN(new_n650));
  NOR2_X1   g449(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n648), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n654), .A2(KEYINPUT42), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n654), .A2(KEYINPUT42), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n650), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT107), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n650), .B(new_n659), .C1(new_n655), .C2(new_n656), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(G1325gat));
  INV_X1    g460(.A(KEYINPUT108), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n488), .B2(new_n492), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n487), .B1(new_n426), .B2(new_n427), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n491), .A2(KEYINPUT36), .A3(new_n425), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n664), .A2(new_n665), .A3(KEYINPUT108), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n644), .A2(G15gat), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(G15gat), .B1(new_n644), .B2(new_n428), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(G1326gat));
  OR3_X1    g470(.A1(new_n643), .A2(KEYINPUT109), .A3(new_n308), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT109), .B1(new_n643), .B2(new_n308), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT43), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(G22gat), .ZN(G1327gat));
  NAND2_X1  g475(.A1(new_n461), .A2(KEYINPUT112), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n484), .A2(new_n667), .A3(new_n486), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(KEYINPUT111), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT111), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n484), .A2(new_n667), .A3(new_n486), .A4(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT112), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n450), .A2(new_n460), .A3(new_n682), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n677), .A2(new_n679), .A3(new_n681), .A4(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(new_n685), .A3(new_n641), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n494), .A2(new_n641), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT44), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n602), .A2(new_n617), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT110), .Z(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(G29gat), .B1(new_n692), .B2(new_n359), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n687), .A2(new_n690), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n694), .A2(new_n504), .A3(new_n645), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT45), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n696), .ZN(G1328gat));
  NAND3_X1  g496(.A1(new_n694), .A2(new_n505), .A3(new_n447), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n698), .B(KEYINPUT46), .Z(new_n699));
  OAI21_X1  g498(.A(G36gat), .B1(new_n692), .B2(new_n448), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(G1329gat));
  NAND2_X1  g500(.A1(new_n668), .A2(G43gat), .ZN(new_n702));
  INV_X1    g501(.A(new_n694), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n703), .A2(new_n451), .ZN(new_n704));
  OAI22_X1  g503(.A1(new_n692), .A2(new_n702), .B1(new_n704), .B2(G43gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g505(.A1(new_n703), .A2(G50gat), .A3(new_n308), .ZN(new_n707));
  INV_X1    g506(.A(new_n308), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n689), .A2(new_n708), .A3(new_n691), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n707), .B1(new_n709), .B2(G50gat), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g510(.A1(new_n617), .A2(new_n641), .A3(new_n549), .ZN(new_n712));
  AND3_X1   g511(.A1(new_n684), .A2(new_n601), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n645), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT113), .B(G57gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1332gat));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n447), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT49), .B(G64gat), .Z(new_n719));
  OAI21_X1  g518(.A(new_n718), .B1(new_n717), .B2(new_n719), .ZN(G1333gat));
  AND2_X1   g519(.A1(new_n713), .A2(new_n428), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n721), .A2(G71gat), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n713), .A2(G71gat), .A3(new_n668), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT50), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT50), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n722), .A2(new_n726), .A3(new_n723), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(G1334gat));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n708), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(G78gat), .ZN(G1335gat));
  INV_X1    g529(.A(new_n617), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(new_n549), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n689), .A2(new_n601), .A3(new_n732), .ZN(new_n733));
  OR3_X1    g532(.A1(new_n733), .A2(KEYINPUT114), .A3(new_n359), .ZN(new_n734));
  OAI21_X1  g533(.A(KEYINPUT114), .B1(new_n733), .B2(new_n359), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n734), .A2(G85gat), .A3(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n601), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n359), .A2(new_n737), .A3(G85gat), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT115), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n684), .A2(new_n739), .A3(new_n641), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n739), .B1(new_n684), .B2(new_n641), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT51), .B1(new_n742), .B2(new_n732), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n679), .A2(new_n681), .ZN(new_n744));
  AND3_X1   g543(.A1(new_n450), .A2(new_n682), .A3(new_n460), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n682), .B1(new_n450), .B2(new_n460), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n744), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n636), .A2(new_n640), .ZN(new_n748));
  OAI21_X1  g547(.A(KEYINPUT115), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n684), .A2(new_n739), .A3(new_n641), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n749), .A2(KEYINPUT51), .A3(new_n732), .A4(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n738), .B1(new_n743), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n736), .A2(new_n753), .ZN(G1336gat));
  NAND2_X1  g553(.A1(new_n601), .A2(new_n447), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(G92gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n743), .B2(new_n752), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758));
  OAI21_X1  g557(.A(G92gat), .B1(new_n733), .B2(new_n448), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n756), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n749), .A2(new_n732), .A3(new_n750), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n761), .B1(new_n764), .B2(new_n751), .ZN(new_n765));
  INV_X1    g564(.A(new_n732), .ZN(new_n766));
  AOI211_X1 g565(.A(new_n737), .B(new_n766), .C1(new_n686), .C2(new_n688), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n443), .B1(new_n767), .B2(new_n447), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT52), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n760), .A2(new_n769), .ZN(G1337gat));
  NOR3_X1   g569(.A1(new_n451), .A2(G99gat), .A3(new_n737), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(new_n743), .B2(new_n752), .ZN(new_n772));
  OAI21_X1  g571(.A(G99gat), .B1(new_n733), .B2(new_n667), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(G1338gat));
  NOR3_X1   g573(.A1(new_n308), .A2(G106gat), .A3(new_n737), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(new_n743), .B2(new_n752), .ZN(new_n776));
  INV_X1    g575(.A(G106gat), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n767), .B2(new_n708), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n776), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n780), .ZN(new_n782));
  INV_X1    g581(.A(new_n775), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n783), .B1(new_n764), .B2(new_n751), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n782), .B1(new_n784), .B2(new_n778), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n781), .A2(new_n785), .ZN(G1339gat));
  NAND2_X1  g585(.A1(new_n593), .A2(new_n555), .ZN(new_n787));
  OAI211_X1 g586(.A(KEYINPUT54), .B(new_n787), .C1(new_n592), .C2(new_n595), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789));
  XNOR2_X1  g588(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n553), .B1(new_n598), .B2(new_n790), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n789), .B1(new_n788), .B2(new_n791), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n596), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n528), .B1(new_n525), .B2(new_n527), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n530), .A2(new_n531), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n541), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n546), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n748), .A2(new_n794), .A3(new_n798), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n549), .B(new_n596), .C1(new_n793), .C2(new_n792), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n601), .A2(new_n546), .A3(new_n797), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n641), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n617), .B1(new_n799), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n712), .A2(new_n737), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n359), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AND3_X1   g604(.A1(new_n805), .A2(new_n448), .A3(new_n458), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n549), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n807), .A2(KEYINPUT118), .A3(new_n311), .ZN(new_n808));
  XNOR2_X1  g607(.A(KEYINPUT118), .B(G113gat), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n808), .B1(new_n807), .B2(new_n809), .ZN(G1340gat));
  NAND2_X1  g609(.A1(new_n806), .A2(new_n601), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g611(.A1(new_n806), .A2(new_n731), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(new_n316), .ZN(new_n814));
  XOR2_X1   g613(.A(new_n814), .B(KEYINPUT119), .Z(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n316), .B2(new_n813), .ZN(G1342gat));
  INV_X1    g615(.A(KEYINPUT56), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n806), .B(new_n641), .C1(new_n817), .C2(new_n319), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n319), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n818), .B(new_n819), .ZN(G1343gat));
  NAND2_X1  g619(.A1(new_n803), .A2(new_n804), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n667), .A2(new_n708), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n822), .A2(KEYINPUT121), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(KEYINPUT121), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n821), .A2(new_n645), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT122), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n805), .A2(KEYINPUT122), .A3(new_n823), .A4(new_n824), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n447), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n550), .A2(G141gat), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT58), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT57), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n821), .A2(new_n832), .A3(new_n708), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n668), .A2(new_n359), .A3(new_n447), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n794), .A2(KEYINPUT120), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT120), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n836), .B(new_n596), .C1(new_n792), .C2(new_n793), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n835), .A2(new_n549), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n641), .B1(new_n838), .B2(new_n801), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n617), .B1(new_n839), .B2(new_n799), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n308), .B1(new_n840), .B2(new_n804), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n833), .B(new_n834), .C1(new_n841), .C2(new_n832), .ZN(new_n842));
  OAI21_X1  g641(.A(G141gat), .B1(new_n842), .B2(new_n550), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n831), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n825), .A2(new_n447), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(new_n830), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n845), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT123), .B1(new_n844), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT123), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n831), .A2(new_n843), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n843), .A2(new_n847), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n850), .B(new_n851), .C1(new_n852), .C2(new_n845), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n849), .A2(new_n853), .ZN(G1344gat));
  NAND2_X1  g653(.A1(new_n840), .A2(new_n804), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT57), .B1(new_n855), .B2(new_n708), .ZN(new_n856));
  AOI211_X1 g655(.A(new_n832), .B(new_n308), .C1(new_n803), .C2(new_n804), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n858), .A2(new_n601), .A3(new_n834), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n206), .B1(new_n859), .B2(KEYINPUT59), .ZN(new_n860));
  OR3_X1    g659(.A1(new_n842), .A2(KEYINPUT59), .A3(new_n737), .ZN(new_n861));
  AOI21_X1  g660(.A(G148gat), .B1(new_n829), .B2(new_n601), .ZN(new_n862));
  AOI22_X1  g661(.A1(new_n860), .A2(new_n861), .B1(KEYINPUT59), .B2(new_n862), .ZN(G1345gat));
  AOI21_X1  g662(.A(G155gat), .B1(new_n829), .B2(new_n731), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n842), .A2(new_n212), .A3(new_n617), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(G1346gat));
  NAND3_X1  g665(.A1(new_n829), .A2(new_n213), .A3(new_n641), .ZN(new_n867));
  OAI21_X1  g666(.A(G162gat), .B1(new_n842), .B2(new_n748), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1347gat));
  AND2_X1   g668(.A1(new_n821), .A2(new_n458), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n645), .A2(new_n448), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n550), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(new_n361), .ZN(G1348gat));
  NOR2_X1   g673(.A1(new_n872), .A2(new_n737), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(new_n362), .ZN(G1349gat));
  OAI21_X1  g675(.A(G183gat), .B1(new_n872), .B2(new_n617), .ZN(new_n877));
  NAND2_X1  g676(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n870), .A2(new_n375), .A3(new_n731), .A4(new_n871), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n880), .B(new_n881), .Z(G1350gat));
  XNOR2_X1  g681(.A(KEYINPUT61), .B(G190gat), .ZN(new_n883));
  NAND2_X1  g682(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n872), .A2(new_n748), .ZN(new_n885));
  MUX2_X1   g684(.A(new_n883), .B(new_n884), .S(new_n885), .Z(G1351gat));
  AND2_X1   g685(.A1(new_n667), .A2(new_n871), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n821), .A2(new_n708), .A3(new_n887), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT125), .Z(new_n889));
  INV_X1    g688(.A(G197gat), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n889), .A2(new_n890), .A3(new_n549), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n858), .A2(new_n887), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n892), .A2(new_n549), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n891), .B1(new_n893), .B2(new_n890), .ZN(G1352gat));
  NAND3_X1  g693(.A1(new_n858), .A2(new_n601), .A3(new_n887), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n895), .A2(KEYINPUT126), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(KEYINPUT126), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(G204gat), .A3(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(new_n822), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n755), .A2(G204gat), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n821), .A2(new_n359), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  XOR2_X1   g700(.A(new_n901), .B(KEYINPUT62), .Z(new_n902));
  NAND2_X1  g701(.A1(new_n898), .A2(new_n902), .ZN(G1353gat));
  AOI21_X1  g702(.A(new_n617), .B1(new_n240), .B2(new_n242), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n731), .B(new_n887), .C1(new_n856), .C2(new_n857), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n906), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT63), .B1(new_n906), .B2(G211gat), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(KEYINPUT127), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT127), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n911), .B(new_n905), .C1(new_n907), .C2(new_n908), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(G1354gat));
  AOI21_X1  g712(.A(G218gat), .B1(new_n889), .B2(new_n641), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n748), .A2(new_n230), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n914), .B1(new_n892), .B2(new_n915), .ZN(G1355gat));
endmodule


