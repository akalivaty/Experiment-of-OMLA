

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804;

  NAND2_X1 U376 ( .A1(n384), .A2(n382), .ZN(n683) );
  NOR2_X2 U377 ( .A1(n585), .A2(n560), .ZN(n563) );
  XNOR2_X2 U378 ( .A(n557), .B(n556), .ZN(n585) );
  XNOR2_X2 U379 ( .A(n648), .B(KEYINPUT1), .ZN(n730) );
  NAND2_X1 U380 ( .A1(n494), .A2(n591), .ZN(n411) );
  XNOR2_X1 U381 ( .A(n407), .B(n363), .ZN(n777) );
  AND2_X1 U382 ( .A1(n386), .A2(n356), .ZN(n384) );
  XNOR2_X1 U383 ( .A(n705), .B(n706), .ZN(n707) );
  XOR2_X1 U384 ( .A(KEYINPUT59), .B(n692), .Z(n693) );
  XNOR2_X1 U385 ( .A(n566), .B(n565), .ZN(n794) );
  XNOR2_X1 U386 ( .A(n443), .B(KEYINPUT69), .ZN(n542) );
  NAND2_X1 U387 ( .A1(n401), .A2(n435), .ZN(n355) );
  NAND2_X1 U388 ( .A1(n401), .A2(n435), .ZN(n714) );
  BUF_X2 U389 ( .A(n703), .Z(n697) );
  OR2_X1 U390 ( .A1(n621), .A2(n455), .ZN(n426) );
  XNOR2_X2 U391 ( .A(n602), .B(n588), .ZN(n718) );
  XNOR2_X1 U392 ( .A(n505), .B(n551), .ZN(n566) );
  INV_X1 U393 ( .A(KEYINPUT47), .ZN(n461) );
  INV_X1 U394 ( .A(KEYINPUT87), .ZN(n463) );
  INV_X1 U395 ( .A(n766), .ZN(n436) );
  XNOR2_X1 U396 ( .A(KEYINPUT15), .B(G902), .ZN(n612) );
  NOR2_X1 U397 ( .A1(G237), .A2(G902), .ZN(n554) );
  XNOR2_X1 U398 ( .A(n542), .B(n442), .ZN(n441) );
  XNOR2_X1 U399 ( .A(KEYINPUT5), .B(G137), .ZN(n442) );
  XNOR2_X1 U400 ( .A(n419), .B(KEYINPUT70), .ZN(n729) );
  BUF_X1 U401 ( .A(n729), .Z(n414) );
  OR2_X1 U402 ( .A1(n620), .A2(n622), .ZN(n455) );
  INV_X1 U403 ( .A(G472), .ZN(n440) );
  INV_X1 U404 ( .A(n637), .ZN(n383) );
  NAND2_X1 U405 ( .A1(n380), .A2(n587), .ZN(n379) );
  INV_X1 U406 ( .A(n654), .ZN(n394) );
  NOR2_X1 U407 ( .A1(n652), .A2(n653), .ZN(n390) );
  XNOR2_X1 U408 ( .A(n445), .B(n498), .ZN(n444) );
  XNOR2_X1 U409 ( .A(n496), .B(G146), .ZN(n445) );
  XNOR2_X1 U410 ( .A(KEYINPUT79), .B(KEYINPUT104), .ZN(n496) );
  XNOR2_X1 U411 ( .A(G113), .B(KEYINPUT98), .ZN(n499) );
  INV_X1 U412 ( .A(KEYINPUT23), .ZN(n520) );
  XNOR2_X1 U413 ( .A(G146), .B(G125), .ZN(n546) );
  INV_X1 U414 ( .A(G101), .ZN(n443) );
  XNOR2_X1 U415 ( .A(KEYINPUT71), .B(KEYINPUT4), .ZN(n503) );
  INV_X1 U416 ( .A(G210), .ZN(n555) );
  XNOR2_X1 U417 ( .A(n481), .B(n480), .ZN(n592) );
  XNOR2_X1 U418 ( .A(n479), .B(n478), .ZN(n480) );
  INV_X1 U419 ( .A(G140), .ZN(n529) );
  BUF_X1 U420 ( .A(n585), .Z(n602) );
  NAND2_X1 U421 ( .A1(n413), .A2(n717), .ZN(n412) );
  XNOR2_X1 U422 ( .A(n615), .B(n420), .ZN(n748) );
  XNOR2_X1 U423 ( .A(KEYINPUT111), .B(KEYINPUT33), .ZN(n420) );
  XNOR2_X1 U424 ( .A(n400), .B(n449), .ZN(n448) );
  OR2_X1 U425 ( .A1(n410), .A2(n560), .ZN(n400) );
  OR2_X1 U426 ( .A1(n427), .A2(KEYINPUT67), .ZN(n385) );
  INV_X1 U427 ( .A(KEYINPUT22), .ZN(n458) );
  NAND2_X1 U428 ( .A1(n668), .A2(n389), .ZN(n715) );
  AND2_X1 U429 ( .A1(n667), .A2(KEYINPUT2), .ZN(n668) );
  INV_X1 U430 ( .A(KEYINPUT86), .ZN(n416) );
  NOR2_X1 U431 ( .A1(n375), .A2(n374), .ZN(n373) );
  INV_X1 U432 ( .A(KEYINPUT91), .ZN(n596) );
  NAND2_X1 U433 ( .A1(n423), .A2(n726), .ZN(n727) );
  INV_X1 U434 ( .A(G110), .ZN(n519) );
  NOR2_X1 U435 ( .A1(n397), .A2(n653), .ZN(n391) );
  XNOR2_X1 U436 ( .A(n421), .B(KEYINPUT20), .ZN(n534) );
  XNOR2_X1 U437 ( .A(n368), .B(G122), .ZN(n467) );
  INV_X1 U438 ( .A(KEYINPUT12), .ZN(n368) );
  XNOR2_X1 U439 ( .A(G113), .B(G104), .ZN(n466) );
  XNOR2_X1 U440 ( .A(G143), .B(G140), .ZN(n469) );
  XNOR2_X1 U441 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n545) );
  INV_X1 U442 ( .A(KEYINPUT48), .ZN(n460) );
  NAND2_X1 U443 ( .A1(G234), .A2(G237), .ZN(n510) );
  NAND2_X1 U444 ( .A1(n718), .A2(n717), .ZN(n721) );
  NOR2_X1 U445 ( .A1(n734), .A2(n439), .ZN(n735) );
  INV_X1 U446 ( .A(n599), .ZN(n413) );
  XNOR2_X1 U447 ( .A(n643), .B(KEYINPUT110), .ZN(n410) );
  INV_X1 U448 ( .A(G902), .ZN(n533) );
  INV_X1 U449 ( .A(n456), .ZN(n454) );
  XNOR2_X1 U450 ( .A(n566), .B(n433), .ZN(n672) );
  XNOR2_X1 U451 ( .A(n434), .B(n501), .ZN(n433) );
  XNOR2_X1 U452 ( .A(n444), .B(n441), .ZN(n434) );
  XNOR2_X1 U453 ( .A(KEYINPUT16), .B(G122), .ZN(n539) );
  XNOR2_X1 U454 ( .A(G128), .B(G119), .ZN(n523) );
  XNOR2_X1 U455 ( .A(G116), .B(G122), .ZN(n483) );
  XOR2_X1 U456 ( .A(KEYINPUT107), .B(KEYINPUT7), .Z(n484) );
  XNOR2_X1 U457 ( .A(G134), .B(G107), .ZN(n482) );
  XNOR2_X1 U458 ( .A(n432), .B(n430), .ZN(n528) );
  XNOR2_X1 U459 ( .A(KEYINPUT8), .B(KEYINPUT72), .ZN(n432) );
  NOR2_X1 U460 ( .A1(n431), .A2(G953), .ZN(n430) );
  INV_X1 U461 ( .A(G234), .ZN(n431) );
  INV_X1 U462 ( .A(G131), .ZN(n473) );
  XNOR2_X1 U463 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n474) );
  NOR2_X1 U464 ( .A1(n406), .A2(n405), .ZN(n408) );
  XNOR2_X1 U465 ( .A(n403), .B(n362), .ZN(n747) );
  NOR2_X1 U466 ( .A1(n720), .A2(n560), .ZN(n402) );
  XNOR2_X1 U467 ( .A(n437), .B(KEYINPUT28), .ZN(n575) );
  NOR2_X1 U468 ( .A1(n410), .A2(n599), .ZN(n437) );
  XNOR2_X1 U469 ( .A(n563), .B(n562), .ZN(n621) );
  XOR2_X1 U470 ( .A(n561), .B(KEYINPUT19), .Z(n562) );
  NOR2_X1 U471 ( .A1(n414), .A2(n439), .ZN(n650) );
  INV_X1 U472 ( .A(KEYINPUT6), .ZN(n438) );
  INV_X1 U473 ( .A(G953), .ZN(n795) );
  XNOR2_X1 U474 ( .A(n676), .B(KEYINPUT97), .ZN(n709) );
  INV_X1 U475 ( .A(KEYINPUT36), .ZN(n369) );
  NOR2_X1 U476 ( .A1(n605), .A2(n602), .ZN(n603) );
  AND2_X1 U477 ( .A1(n448), .A2(n425), .ZN(n424) );
  AND2_X1 U478 ( .A1(n586), .A2(n583), .ZN(n425) );
  NAND2_X1 U479 ( .A1(n383), .A2(n388), .ZN(n382) );
  NOR2_X1 U480 ( .A1(n753), .A2(n752), .ZN(n754) );
  AND2_X1 U481 ( .A1(n385), .A2(n423), .ZN(n356) );
  XOR2_X1 U482 ( .A(n536), .B(n535), .Z(n357) );
  AND2_X1 U483 ( .A1(n457), .A2(n453), .ZN(n358) );
  XNOR2_X1 U484 ( .A(n509), .B(n508), .ZN(n726) );
  AND2_X1 U485 ( .A1(n682), .A2(n415), .ZN(n359) );
  AND2_X1 U486 ( .A1(n426), .A2(n456), .ZN(n360) );
  INV_X1 U487 ( .A(n640), .ZN(n423) );
  XNOR2_X1 U488 ( .A(n537), .B(n357), .ZN(n640) );
  AND2_X1 U489 ( .A1(n579), .A2(KEYINPUT87), .ZN(n361) );
  INV_X1 U490 ( .A(KEYINPUT67), .ZN(n388) );
  XOR2_X1 U491 ( .A(KEYINPUT114), .B(KEYINPUT41), .Z(n362) );
  XOR2_X1 U492 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n363) );
  XOR2_X1 U493 ( .A(n596), .B(KEYINPUT46), .Z(n364) );
  INV_X1 U494 ( .A(KEYINPUT2), .ZN(n435) );
  INV_X1 U495 ( .A(KEYINPUT76), .ZN(n587) );
  NAND2_X1 U496 ( .A1(n409), .A2(n408), .ZN(n407) );
  NAND2_X1 U497 ( .A1(n365), .A2(n448), .ZN(n370) );
  AND2_X2 U498 ( .A1(n399), .A2(n584), .ZN(n365) );
  AND2_X1 U499 ( .A1(n730), .A2(n410), .ZN(n427) );
  INV_X1 U500 ( .A(n366), .ZN(n662) );
  NOR2_X1 U501 ( .A1(n660), .A2(n658), .ZN(n366) );
  NAND2_X1 U502 ( .A1(n429), .A2(n637), .ZN(n428) );
  XNOR2_X2 U503 ( .A(n459), .B(n458), .ZN(n637) );
  XNOR2_X2 U504 ( .A(n367), .B(n636), .ZN(n660) );
  NAND2_X1 U505 ( .A1(n680), .A2(n683), .ZN(n367) );
  XNOR2_X1 U506 ( .A(n603), .B(n369), .ZN(n604) );
  NOR2_X1 U507 ( .A1(n648), .A2(n729), .ZN(n582) );
  XNOR2_X2 U508 ( .A(n572), .B(n571), .ZN(n648) );
  NAND2_X1 U509 ( .A1(n662), .A2(n661), .ZN(n404) );
  NAND2_X1 U510 ( .A1(n631), .A2(n423), .ZN(n632) );
  NOR2_X1 U511 ( .A1(n598), .A2(n412), .ZN(n601) );
  XNOR2_X2 U512 ( .A(n370), .B(n589), .ZN(n610) );
  NAND2_X1 U513 ( .A1(n372), .A2(n371), .ZN(n447) );
  NAND2_X1 U514 ( .A1(n373), .A2(n359), .ZN(n371) );
  NAND2_X1 U515 ( .A1(n376), .A2(n682), .ZN(n372) );
  NAND2_X1 U516 ( .A1(n580), .A2(KEYINPUT76), .ZN(n374) );
  INV_X1 U517 ( .A(n381), .ZN(n375) );
  NAND2_X1 U518 ( .A1(n379), .A2(n377), .ZN(n376) );
  NAND2_X1 U519 ( .A1(n378), .A2(n587), .ZN(n377) );
  NAND2_X1 U520 ( .A1(n381), .A2(n580), .ZN(n378) );
  INV_X1 U521 ( .A(n415), .ZN(n380) );
  NAND2_X1 U522 ( .A1(n462), .A2(n461), .ZN(n381) );
  NAND2_X1 U523 ( .A1(n637), .A2(n387), .ZN(n386) );
  AND2_X1 U524 ( .A1(n427), .A2(KEYINPUT67), .ZN(n387) );
  INV_X1 U525 ( .A(n777), .ZN(n389) );
  AND2_X2 U526 ( .A1(n777), .A2(n435), .ZN(n712) );
  NOR2_X1 U527 ( .A1(n390), .A2(n394), .ZN(n393) );
  AND2_X1 U528 ( .A1(n652), .A2(n653), .ZN(n396) );
  NOR2_X1 U529 ( .A1(n392), .A2(n391), .ZN(n655) );
  NAND2_X1 U530 ( .A1(n395), .A2(n393), .ZN(n392) );
  NAND2_X1 U531 ( .A1(n396), .A2(n397), .ZN(n395) );
  INV_X1 U532 ( .A(n774), .ZN(n397) );
  NAND2_X1 U533 ( .A1(n398), .A2(n803), .ZN(n597) );
  XNOR2_X1 U534 ( .A(n398), .B(G131), .ZN(G33) );
  XNOR2_X2 U535 ( .A(n590), .B(KEYINPUT40), .ZN(n398) );
  AND2_X2 U536 ( .A1(n718), .A2(n583), .ZN(n399) );
  XNOR2_X1 U537 ( .A(n582), .B(n581), .ZN(n584) );
  XNOR2_X1 U538 ( .A(n401), .B(n797), .ZN(n796) );
  XNOR2_X2 U539 ( .A(n665), .B(KEYINPUT90), .ZN(n401) );
  NAND2_X1 U540 ( .A1(n718), .A2(n402), .ZN(n403) );
  INV_X1 U541 ( .A(n747), .ZN(n594) );
  NAND2_X1 U542 ( .A1(n404), .A2(n663), .ZN(n409) );
  INV_X1 U543 ( .A(n656), .ZN(n405) );
  NAND2_X1 U544 ( .A1(n451), .A2(n452), .ZN(n406) );
  NOR2_X1 U545 ( .A1(n629), .A2(n454), .ZN(n453) );
  NAND2_X2 U546 ( .A1(n358), .A2(n426), .ZN(n459) );
  XNOR2_X1 U547 ( .A(n597), .B(n364), .ZN(n418) );
  XNOR2_X2 U548 ( .A(n411), .B(KEYINPUT109), .ZN(n771) );
  NAND2_X2 U549 ( .A1(n610), .A2(n771), .ZN(n590) );
  NOR2_X1 U550 ( .A1(n436), .A2(n361), .ZN(n415) );
  XNOR2_X1 U551 ( .A(n417), .B(n416), .ZN(n716) );
  NAND2_X1 U552 ( .A1(n713), .A2(n355), .ZN(n417) );
  NAND2_X1 U553 ( .A1(n418), .A2(n447), .ZN(n446) );
  NAND2_X1 U554 ( .A1(n640), .A2(n627), .ZN(n419) );
  NAND2_X1 U555 ( .A1(n672), .A2(n533), .ZN(n506) );
  NAND2_X1 U556 ( .A1(n768), .A2(n654), .ZN(n464) );
  NAND2_X1 U557 ( .A1(n802), .A2(KEYINPUT44), .ZN(n452) );
  XNOR2_X2 U558 ( .A(n626), .B(KEYINPUT35), .ZN(n802) );
  NAND2_X1 U559 ( .A1(n768), .A2(n577), .ZN(n578) );
  XNOR2_X2 U560 ( .A(n576), .B(KEYINPUT85), .ZN(n768) );
  NAND2_X1 U561 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U562 ( .A1(n538), .A2(n423), .ZN(n599) );
  XNOR2_X1 U563 ( .A(n446), .B(n460), .ZN(n422) );
  NAND2_X1 U564 ( .A1(n612), .A2(G234), .ZN(n421) );
  NAND2_X1 U565 ( .A1(n422), .A2(n611), .ZN(n665) );
  NAND2_X1 U566 ( .A1(n584), .A2(n424), .ZN(n766) );
  XNOR2_X2 U567 ( .A(n428), .B(n635), .ZN(n680) );
  NOR2_X1 U568 ( .A1(n633), .A2(n632), .ZN(n429) );
  XNOR2_X2 U569 ( .A(n487), .B(G128), .ZN(n504) );
  XNOR2_X2 U570 ( .A(n504), .B(n503), .ZN(n551) );
  XNOR2_X1 U571 ( .A(n643), .B(n438), .ZN(n638) );
  INV_X1 U572 ( .A(n643), .ZN(n439) );
  XNOR2_X2 U573 ( .A(n506), .B(n440), .ZN(n643) );
  INV_X1 U574 ( .A(KEYINPUT30), .ZN(n449) );
  XNOR2_X1 U575 ( .A(n450), .B(G119), .ZN(n500) );
  XNOR2_X2 U576 ( .A(G116), .B(KEYINPUT3), .ZN(n450) );
  NAND2_X1 U577 ( .A1(n660), .A2(KEYINPUT44), .ZN(n451) );
  NAND2_X1 U578 ( .A1(n360), .A2(n457), .ZN(n630) );
  NAND2_X1 U579 ( .A1(n620), .A2(n622), .ZN(n456) );
  NAND2_X1 U580 ( .A1(n621), .A2(n622), .ZN(n457) );
  NAND2_X1 U581 ( .A1(n464), .A2(n463), .ZN(n462) );
  INV_X1 U582 ( .A(n575), .ZN(n593) );
  OR2_X1 U583 ( .A1(n784), .A2(n569), .ZN(n544) );
  NOR2_X1 U584 ( .A1(n593), .A2(n648), .ZN(n465) );
  INV_X1 U585 ( .A(KEYINPUT94), .ZN(n659) );
  XNOR2_X1 U586 ( .A(n469), .B(n468), .ZN(n470) );
  INV_X1 U587 ( .A(KEYINPUT24), .ZN(n525) );
  INV_X1 U588 ( .A(G475), .ZN(n478) );
  INV_X1 U589 ( .A(n564), .ZN(n565) );
  INV_X1 U590 ( .A(n573), .ZN(n574) );
  XNOR2_X1 U591 ( .A(n689), .B(n688), .ZN(n690) );
  INV_X1 U592 ( .A(KEYINPUT63), .ZN(n678) );
  XNOR2_X1 U593 ( .A(n467), .B(n466), .ZN(n471) );
  INV_X1 U594 ( .A(KEYINPUT11), .ZN(n468) );
  XNOR2_X1 U595 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U596 ( .A(n546), .B(KEYINPUT10), .ZN(n792) );
  XNOR2_X1 U597 ( .A(n472), .B(n792), .ZN(n477) );
  NOR2_X1 U598 ( .A1(G953), .A2(G237), .ZN(n497) );
  NAND2_X1 U599 ( .A1(G214), .A2(n497), .ZN(n475) );
  XNOR2_X1 U600 ( .A(n474), .B(n473), .ZN(n502) );
  XOR2_X1 U601 ( .A(n475), .B(n502), .Z(n476) );
  XNOR2_X1 U602 ( .A(n477), .B(n476), .ZN(n692) );
  NOR2_X1 U603 ( .A1(G902), .A2(n692), .ZN(n481) );
  XNOR2_X1 U604 ( .A(KEYINPUT106), .B(KEYINPUT13), .ZN(n479) );
  INV_X1 U605 ( .A(n592), .ZN(n494) );
  XNOR2_X1 U606 ( .A(n482), .B(KEYINPUT9), .ZN(n486) );
  XNOR2_X1 U607 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U608 ( .A(n486), .B(n485), .Z(n491) );
  NAND2_X1 U609 ( .A1(G217), .A2(n528), .ZN(n489) );
  XNOR2_X2 U610 ( .A(KEYINPUT65), .B(G143), .ZN(n487) );
  INV_X1 U611 ( .A(n504), .ZN(n488) );
  XNOR2_X1 U612 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U613 ( .A(n491), .B(n490), .ZN(n689) );
  NAND2_X1 U614 ( .A1(n689), .A2(n533), .ZN(n493) );
  XOR2_X1 U615 ( .A(KEYINPUT108), .B(G478), .Z(n492) );
  XNOR2_X1 U616 ( .A(n493), .B(n492), .ZN(n591) );
  NOR2_X1 U617 ( .A1(n591), .A2(n494), .ZN(n773) );
  NOR2_X1 U618 ( .A1(n771), .A2(n773), .ZN(n722) );
  INV_X1 U619 ( .A(KEYINPUT88), .ZN(n495) );
  XNOR2_X1 U620 ( .A(n722), .B(n495), .ZN(n654) );
  NAND2_X1 U621 ( .A1(n497), .A2(G210), .ZN(n498) );
  XNOR2_X1 U622 ( .A(n500), .B(n499), .ZN(n540) );
  BUF_X1 U623 ( .A(n540), .Z(n501) );
  XNOR2_X1 U624 ( .A(n502), .B(G134), .ZN(n505) );
  NAND2_X1 U625 ( .A1(n534), .A2(G221), .ZN(n507) );
  XNOR2_X1 U626 ( .A(n507), .B(KEYINPUT21), .ZN(n509) );
  INV_X1 U627 ( .A(KEYINPUT103), .ZN(n508) );
  INV_X1 U628 ( .A(n726), .ZN(n627) );
  XNOR2_X1 U629 ( .A(n510), .B(KEYINPUT14), .ZN(n514) );
  NAND2_X1 U630 ( .A1(G952), .A2(n514), .ZN(n511) );
  XNOR2_X1 U631 ( .A(n511), .B(KEYINPUT99), .ZN(n745) );
  NAND2_X1 U632 ( .A1(n745), .A2(n795), .ZN(n513) );
  INV_X1 U633 ( .A(KEYINPUT100), .ZN(n512) );
  XNOR2_X1 U634 ( .A(n513), .B(n512), .ZN(n619) );
  INV_X1 U635 ( .A(n619), .ZN(n517) );
  NAND2_X1 U636 ( .A1(G902), .A2(n514), .ZN(n616) );
  NOR2_X1 U637 ( .A1(G900), .A2(n616), .ZN(n515) );
  NAND2_X1 U638 ( .A1(G953), .A2(n515), .ZN(n516) );
  NAND2_X1 U639 ( .A1(n517), .A2(n516), .ZN(n583) );
  NAND2_X1 U640 ( .A1(n627), .A2(n583), .ZN(n518) );
  XNOR2_X1 U641 ( .A(KEYINPUT75), .B(n518), .ZN(n538) );
  NAND2_X1 U642 ( .A1(KEYINPUT23), .A2(n519), .ZN(n522) );
  NAND2_X1 U643 ( .A1(n520), .A2(G110), .ZN(n521) );
  NAND2_X1 U644 ( .A1(n522), .A2(n521), .ZN(n524) );
  XNOR2_X1 U645 ( .A(n524), .B(n523), .ZN(n526) );
  XNOR2_X1 U646 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U647 ( .A(n527), .B(n792), .ZN(n532) );
  NAND2_X1 U648 ( .A1(G221), .A2(n528), .ZN(n530) );
  XNOR2_X1 U649 ( .A(n529), .B(G137), .ZN(n564) );
  XNOR2_X1 U650 ( .A(n530), .B(n564), .ZN(n531) );
  XNOR2_X1 U651 ( .A(n532), .B(n531), .ZN(n684) );
  NAND2_X1 U652 ( .A1(n684), .A2(n533), .ZN(n537) );
  AND2_X1 U653 ( .A1(n534), .A2(G217), .ZN(n536) );
  XNOR2_X1 U654 ( .A(KEYINPUT25), .B(KEYINPUT81), .ZN(n535) );
  XNOR2_X1 U655 ( .A(n540), .B(n539), .ZN(n784) );
  XOR2_X1 U656 ( .A(G104), .B(G110), .Z(n541) );
  XNOR2_X1 U657 ( .A(n541), .B(G107), .ZN(n786) );
  XNOR2_X1 U658 ( .A(n786), .B(n542), .ZN(n569) );
  NAND2_X1 U659 ( .A1(n784), .A2(n569), .ZN(n543) );
  NAND2_X1 U660 ( .A1(n544), .A2(n543), .ZN(n553) );
  XNOR2_X1 U661 ( .A(n546), .B(n545), .ZN(n549) );
  NAND2_X1 U662 ( .A1(n795), .A2(G224), .ZN(n547) );
  XNOR2_X1 U663 ( .A(n547), .B(KEYINPUT82), .ZN(n548) );
  XNOR2_X1 U664 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U665 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U666 ( .A(n553), .B(n552), .ZN(n704) );
  NAND2_X1 U667 ( .A1(n704), .A2(n612), .ZN(n557) );
  XNOR2_X1 U668 ( .A(n554), .B(KEYINPUT78), .ZN(n559) );
  OR2_X1 U669 ( .A1(n559), .A2(n555), .ZN(n556) );
  INV_X1 U670 ( .A(G214), .ZN(n558) );
  OR2_X1 U671 ( .A1(n559), .A2(n558), .ZN(n717) );
  INV_X1 U672 ( .A(n717), .ZN(n560) );
  INV_X1 U673 ( .A(KEYINPUT80), .ZN(n561) );
  NAND2_X1 U674 ( .A1(n795), .A2(G227), .ZN(n567) );
  XNOR2_X1 U675 ( .A(n567), .B(G146), .ZN(n568) );
  XNOR2_X1 U676 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U677 ( .A(n794), .B(n570), .ZN(n699) );
  OR2_X2 U678 ( .A1(n699), .A2(G902), .ZN(n572) );
  INV_X1 U679 ( .A(G469), .ZN(n571) );
  OR2_X1 U680 ( .A1(n621), .A2(n648), .ZN(n573) );
  INV_X1 U681 ( .A(n722), .ZN(n579) );
  OR2_X1 U682 ( .A1(KEYINPUT87), .A2(n579), .ZN(n577) );
  NAND2_X1 U683 ( .A1(n578), .A2(KEYINPUT47), .ZN(n580) );
  INV_X1 U684 ( .A(KEYINPUT113), .ZN(n581) );
  INV_X1 U685 ( .A(n602), .ZN(n607) );
  NOR2_X1 U686 ( .A1(n591), .A2(n592), .ZN(n624) );
  AND2_X1 U687 ( .A1(n607), .A2(n624), .ZN(n586) );
  XNOR2_X1 U688 ( .A(KEYINPUT92), .B(KEYINPUT39), .ZN(n589) );
  XOR2_X1 U689 ( .A(KEYINPUT77), .B(KEYINPUT38), .Z(n588) );
  NAND2_X1 U690 ( .A1(n592), .A2(n591), .ZN(n720) );
  NAND2_X1 U691 ( .A1(n594), .A2(n465), .ZN(n595) );
  XNOR2_X1 U692 ( .A(n595), .B(KEYINPUT42), .ZN(n803) );
  INV_X1 U693 ( .A(n771), .ZN(n598) );
  INV_X1 U694 ( .A(n638), .ZN(n600) );
  NAND2_X1 U695 ( .A1(n601), .A2(n600), .ZN(n605) );
  XNOR2_X1 U696 ( .A(n730), .B(KEYINPUT96), .ZN(n633) );
  OR2_X1 U697 ( .A1(n604), .A2(n633), .ZN(n682) );
  INV_X1 U698 ( .A(n730), .ZN(n644) );
  NOR2_X1 U699 ( .A1(n605), .A2(n644), .ZN(n606) );
  XNOR2_X1 U700 ( .A(n606), .B(KEYINPUT43), .ZN(n608) );
  OR2_X1 U701 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U702 ( .A(n609), .B(KEYINPUT112), .ZN(n804) );
  NAND2_X1 U703 ( .A1(n773), .A2(n610), .ZN(n776) );
  AND2_X1 U704 ( .A1(n804), .A2(n776), .ZN(n611) );
  INV_X1 U705 ( .A(n612), .ZN(n613) );
  NAND2_X1 U706 ( .A1(n714), .A2(n613), .ZN(n664) );
  NOR2_X1 U707 ( .A1(n414), .A2(n638), .ZN(n614) );
  NAND2_X1 U708 ( .A1(n614), .A2(n644), .ZN(n615) );
  XNOR2_X1 U709 ( .A(G898), .B(KEYINPUT101), .ZN(n780) );
  NAND2_X1 U710 ( .A1(G953), .A2(n780), .ZN(n787) );
  NOR2_X1 U711 ( .A1(n616), .A2(n787), .ZN(n617) );
  XNOR2_X1 U712 ( .A(n617), .B(KEYINPUT102), .ZN(n618) );
  NOR2_X1 U713 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U714 ( .A(KEYINPUT68), .B(KEYINPUT0), .ZN(n622) );
  NOR2_X1 U715 ( .A1(n748), .A2(n630), .ZN(n623) );
  XNOR2_X1 U716 ( .A(n623), .B(KEYINPUT34), .ZN(n625) );
  NAND2_X1 U717 ( .A1(n625), .A2(n624), .ZN(n626) );
  INV_X1 U718 ( .A(n720), .ZN(n628) );
  NAND2_X1 U719 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U720 ( .A(n638), .B(KEYINPUT84), .ZN(n631) );
  INV_X1 U721 ( .A(KEYINPUT83), .ZN(n634) );
  XNOR2_X1 U722 ( .A(n634), .B(KEYINPUT32), .ZN(n635) );
  INV_X1 U723 ( .A(KEYINPUT95), .ZN(n636) );
  NAND2_X1 U724 ( .A1(n637), .A2(n638), .ZN(n639) );
  XNOR2_X1 U725 ( .A(n639), .B(KEYINPUT93), .ZN(n642) );
  AND2_X1 U726 ( .A1(n640), .A2(n730), .ZN(n641) );
  AND2_X1 U727 ( .A1(n642), .A2(n641), .ZN(n755) );
  INV_X1 U728 ( .A(n630), .ZN(n646) );
  NOR2_X1 U729 ( .A1(n414), .A2(n643), .ZN(n645) );
  AND2_X1 U730 ( .A1(n645), .A2(n644), .ZN(n736) );
  NAND2_X1 U731 ( .A1(n646), .A2(n736), .ZN(n647) );
  XNOR2_X1 U732 ( .A(n647), .B(KEYINPUT31), .ZN(n774) );
  INV_X1 U733 ( .A(n648), .ZN(n649) );
  NAND2_X1 U734 ( .A1(n650), .A2(n649), .ZN(n651) );
  OR2_X1 U735 ( .A1(n630), .A2(n651), .ZN(n652) );
  INV_X1 U736 ( .A(n652), .ZN(n757) );
  INV_X1 U737 ( .A(KEYINPUT105), .ZN(n653) );
  NOR2_X1 U738 ( .A1(n755), .A2(n655), .ZN(n656) );
  INV_X1 U739 ( .A(n802), .ZN(n663) );
  INV_X1 U740 ( .A(KEYINPUT44), .ZN(n657) );
  NAND2_X1 U741 ( .A1(n657), .A2(KEYINPUT94), .ZN(n658) );
  NAND2_X1 U742 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U743 ( .A1(n664), .A2(n712), .ZN(n669) );
  BUF_X1 U744 ( .A(n665), .Z(n666) );
  INV_X1 U745 ( .A(n666), .ZN(n667) );
  NAND2_X1 U746 ( .A1(n669), .A2(n715), .ZN(n671) );
  INV_X1 U747 ( .A(KEYINPUT66), .ZN(n670) );
  XNOR2_X2 U748 ( .A(n671), .B(n670), .ZN(n703) );
  NAND2_X1 U749 ( .A1(n703), .A2(G472), .ZN(n674) );
  XOR2_X1 U750 ( .A(KEYINPUT62), .B(n672), .Z(n673) );
  XNOR2_X1 U751 ( .A(n674), .B(n673), .ZN(n677) );
  INV_X1 U752 ( .A(G952), .ZN(n675) );
  NAND2_X1 U753 ( .A1(n675), .A2(G953), .ZN(n676) );
  NOR2_X2 U754 ( .A1(n677), .A2(n709), .ZN(n679) );
  XNOR2_X1 U755 ( .A(n679), .B(n678), .ZN(G57) );
  XNOR2_X1 U756 ( .A(n680), .B(G119), .ZN(G21) );
  XOR2_X1 U757 ( .A(G125), .B(KEYINPUT37), .Z(n681) );
  XNOR2_X1 U758 ( .A(n682), .B(n681), .ZN(G27) );
  XNOR2_X1 U759 ( .A(n683), .B(G110), .ZN(G12) );
  NAND2_X1 U760 ( .A1(n697), .A2(G217), .ZN(n686) );
  XOR2_X1 U761 ( .A(n684), .B(KEYINPUT124), .Z(n685) );
  XNOR2_X1 U762 ( .A(n686), .B(n685), .ZN(n687) );
  NOR2_X1 U763 ( .A1(n687), .A2(n709), .ZN(G66) );
  NAND2_X1 U764 ( .A1(n697), .A2(G478), .ZN(n688) );
  INV_X1 U765 ( .A(n690), .ZN(n691) );
  NOR2_X1 U766 ( .A1(n691), .A2(n709), .ZN(G63) );
  NAND2_X1 U767 ( .A1(n703), .A2(G475), .ZN(n694) );
  XNOR2_X1 U768 ( .A(n694), .B(n693), .ZN(n695) );
  NOR2_X2 U769 ( .A1(n695), .A2(n709), .ZN(n696) );
  XNOR2_X1 U770 ( .A(n696), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U771 ( .A1(n697), .A2(G469), .ZN(n701) );
  XOR2_X1 U772 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n698) );
  XNOR2_X1 U773 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X1 U774 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U775 ( .A1(n702), .A2(n709), .ZN(G54) );
  NAND2_X1 U776 ( .A1(n703), .A2(G210), .ZN(n708) );
  BUF_X1 U777 ( .A(n704), .Z(n705) );
  XNOR2_X1 U778 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n706) );
  XNOR2_X1 U779 ( .A(n708), .B(n707), .ZN(n710) );
  NOR2_X2 U780 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U781 ( .A(n711), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U782 ( .A(n712), .B(KEYINPUT89), .ZN(n713) );
  AND2_X1 U783 ( .A1(n716), .A2(n715), .ZN(n753) );
  NOR2_X1 U784 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U785 ( .A1(n720), .A2(n719), .ZN(n724) );
  NOR2_X1 U786 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U787 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U788 ( .A1(n725), .A2(n748), .ZN(n741) );
  XOR2_X1 U789 ( .A(KEYINPUT120), .B(KEYINPUT49), .Z(n728) );
  XNOR2_X1 U790 ( .A(n728), .B(n727), .ZN(n733) );
  NAND2_X1 U791 ( .A1(n730), .A2(n414), .ZN(n731) );
  XNOR2_X1 U792 ( .A(n731), .B(KEYINPUT50), .ZN(n732) );
  NAND2_X1 U793 ( .A1(n733), .A2(n732), .ZN(n734) );
  NOR2_X1 U794 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U795 ( .A(n737), .B(KEYINPUT51), .ZN(n738) );
  XNOR2_X1 U796 ( .A(n738), .B(KEYINPUT121), .ZN(n739) );
  NOR2_X1 U797 ( .A1(n747), .A2(n739), .ZN(n740) );
  NOR2_X1 U798 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U799 ( .A(n742), .B(KEYINPUT52), .ZN(n744) );
  XOR2_X1 U800 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n743) );
  XOR2_X1 U801 ( .A(n744), .B(n743), .Z(n746) );
  NAND2_X1 U802 ( .A1(n746), .A2(n745), .ZN(n751) );
  NOR2_X1 U803 ( .A1(n748), .A2(n747), .ZN(n749) );
  NOR2_X1 U804 ( .A1(n749), .A2(G953), .ZN(n750) );
  NAND2_X1 U805 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U806 ( .A(n754), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U807 ( .A(G101), .B(n755), .Z(G3) );
  NAND2_X1 U808 ( .A1(n757), .A2(n771), .ZN(n756) );
  XNOR2_X1 U809 ( .A(n756), .B(G104), .ZN(G6) );
  XOR2_X1 U810 ( .A(KEYINPUT26), .B(KEYINPUT115), .Z(n759) );
  NAND2_X1 U811 ( .A1(n757), .A2(n773), .ZN(n758) );
  XNOR2_X1 U812 ( .A(n759), .B(n758), .ZN(n761) );
  XOR2_X1 U813 ( .A(G107), .B(KEYINPUT27), .Z(n760) );
  XNOR2_X1 U814 ( .A(n761), .B(n760), .ZN(G9) );
  XOR2_X1 U815 ( .A(KEYINPUT117), .B(KEYINPUT29), .Z(n763) );
  NAND2_X1 U816 ( .A1(n768), .A2(n773), .ZN(n762) );
  XNOR2_X1 U817 ( .A(n763), .B(n762), .ZN(n765) );
  XOR2_X1 U818 ( .A(G128), .B(KEYINPUT116), .Z(n764) );
  XNOR2_X1 U819 ( .A(n765), .B(n764), .ZN(G30) );
  XNOR2_X1 U820 ( .A(G143), .B(KEYINPUT118), .ZN(n767) );
  XNOR2_X1 U821 ( .A(n767), .B(n766), .ZN(G45) );
  XOR2_X1 U822 ( .A(G146), .B(KEYINPUT119), .Z(n770) );
  NAND2_X1 U823 ( .A1(n768), .A2(n771), .ZN(n769) );
  XNOR2_X1 U824 ( .A(n770), .B(n769), .ZN(G48) );
  NAND2_X1 U825 ( .A1(n774), .A2(n771), .ZN(n772) );
  XNOR2_X1 U826 ( .A(n772), .B(G113), .ZN(G15) );
  NAND2_X1 U827 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U828 ( .A(n775), .B(G116), .ZN(G18) );
  XNOR2_X1 U829 ( .A(G134), .B(n776), .ZN(G36) );
  NOR2_X1 U830 ( .A1(n777), .A2(G953), .ZN(n782) );
  NAND2_X1 U831 ( .A1(G953), .A2(G224), .ZN(n778) );
  XOR2_X1 U832 ( .A(KEYINPUT61), .B(n778), .Z(n779) );
  NOR2_X1 U833 ( .A1(n780), .A2(n779), .ZN(n781) );
  NOR2_X1 U834 ( .A1(n782), .A2(n781), .ZN(n791) );
  XNOR2_X1 U835 ( .A(G101), .B(KEYINPUT126), .ZN(n783) );
  XNOR2_X1 U836 ( .A(n784), .B(n783), .ZN(n785) );
  XNOR2_X1 U837 ( .A(n786), .B(n785), .ZN(n788) );
  NAND2_X1 U838 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U839 ( .A(n789), .B(KEYINPUT125), .ZN(n790) );
  XOR2_X1 U840 ( .A(n791), .B(n790), .Z(G69) );
  XNOR2_X1 U841 ( .A(n792), .B(KEYINPUT127), .ZN(n793) );
  XNOR2_X1 U842 ( .A(n794), .B(n793), .ZN(n797) );
  NAND2_X1 U843 ( .A1(n796), .A2(n795), .ZN(n801) );
  XNOR2_X1 U844 ( .A(G227), .B(n797), .ZN(n798) );
  NAND2_X1 U845 ( .A1(n798), .A2(G900), .ZN(n799) );
  NAND2_X1 U846 ( .A1(G953), .A2(n799), .ZN(n800) );
  NAND2_X1 U847 ( .A1(n801), .A2(n800), .ZN(G72) );
  XOR2_X1 U848 ( .A(G122), .B(n802), .Z(G24) );
  XNOR2_X1 U849 ( .A(n803), .B(G137), .ZN(G39) );
  XNOR2_X1 U850 ( .A(G140), .B(n804), .ZN(G42) );
endmodule

