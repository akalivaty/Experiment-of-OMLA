//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT1), .B1(new_n187), .B2(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G128), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n187), .A2(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n189), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n191), .A2(new_n192), .A3(new_n195), .A4(G128), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G134), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT65), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT65), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G134), .ZN(new_n201));
  AOI21_X1  g015(.A(G137), .B1(new_n199), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G137), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(G134), .ZN(new_n204));
  OAI21_X1  g018(.A(G131), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n197), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT66), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT11), .ZN(new_n209));
  NOR3_X1   g023(.A1(new_n209), .A2(new_n198), .A3(G137), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n199), .A2(new_n201), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(new_n203), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n210), .B1(new_n212), .B2(new_n209), .ZN(new_n213));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(G134), .ZN(new_n214));
  AOI21_X1  g028(.A(G131), .B1(new_n214), .B2(G137), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n208), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n210), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n217), .B1(new_n202), .B2(KEYINPUT11), .ZN(new_n218));
  INV_X1    g032(.A(G131), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n211), .B2(new_n203), .ZN(new_n220));
  NOR3_X1   g034(.A1(new_n218), .A2(KEYINPUT66), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n207), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(KEYINPUT30), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT66), .B1(new_n218), .B2(new_n220), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n209), .B1(new_n214), .B2(G137), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n226), .A2(new_n215), .A3(new_n208), .A4(new_n217), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n226), .B(new_n217), .C1(new_n203), .C2(new_n211), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n225), .A2(new_n227), .B1(new_n228), .B2(G131), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n191), .A2(new_n192), .A3(KEYINPUT0), .A4(G128), .ZN(new_n230));
  OR2_X1    g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n193), .B1(KEYINPUT64), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(KEYINPUT64), .ZN(new_n233));
  NAND2_X1  g047(.A1(KEYINPUT0), .A2(G128), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n230), .B1(new_n232), .B2(new_n235), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n222), .B(new_n224), .C1(new_n229), .C2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n206), .B1(new_n225), .B2(new_n227), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n228), .A2(G131), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n239), .B1(new_n216), .B2(new_n221), .ZN(new_n240));
  INV_X1    g054(.A(new_n236), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n238), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT67), .B(KEYINPUT30), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n237), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(G116), .B(G119), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT2), .B(G113), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n245), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n242), .A2(new_n248), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT26), .B(G101), .ZN(new_n253));
  NOR2_X1   g067(.A1(G237), .A2(G953), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G210), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n253), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n257));
  XOR2_X1   g071(.A(new_n256), .B(new_n257), .Z(new_n258));
  NAND2_X1  g072(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT29), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n222), .B1(new_n229), .B2(new_n236), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n249), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n251), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT28), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT28), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n251), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n258), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n259), .A2(new_n260), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT70), .ZN(new_n270));
  INV_X1    g084(.A(G902), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n271), .B1(new_n268), .B2(new_n260), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT71), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n274), .B(new_n271), .C1(new_n268), .C2(new_n260), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n259), .A2(new_n268), .A3(new_n276), .A4(new_n260), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n270), .A2(new_n273), .A3(new_n275), .A4(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G472), .ZN(new_n279));
  INV_X1    g093(.A(G472), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT69), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n261), .A2(new_n249), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n282), .B1(new_n245), .B2(new_n249), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n281), .B1(new_n283), .B2(new_n267), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n225), .A2(new_n227), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n236), .B1(new_n285), .B2(new_n239), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n243), .B1(new_n286), .B2(new_n238), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n248), .B1(new_n287), .B2(new_n237), .ZN(new_n288));
  NOR4_X1   g102(.A1(new_n288), .A2(KEYINPUT69), .A3(new_n282), .A4(new_n258), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT31), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n284), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n265), .B1(new_n251), .B2(new_n262), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n282), .A2(KEYINPUT28), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n258), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n250), .A2(new_n251), .A3(new_n267), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n294), .B1(new_n295), .B2(KEYINPUT31), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n280), .B(new_n271), .C1(new_n291), .C2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n297), .A2(KEYINPUT32), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT32), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n295), .A2(KEYINPUT69), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n283), .A2(new_n281), .A3(new_n267), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(KEYINPUT31), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n267), .B1(new_n264), .B2(new_n266), .ZN(new_n303));
  NOR4_X1   g117(.A1(new_n288), .A2(KEYINPUT31), .A3(new_n282), .A4(new_n258), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(G902), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n299), .B1(new_n306), .B2(new_n280), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n279), .B1(new_n298), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G217), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n309), .B1(G234), .B2(new_n271), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(KEYINPUT74), .A2(G125), .ZN(new_n312));
  INV_X1    g126(.A(G140), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(KEYINPUT74), .A2(G125), .A3(G140), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(KEYINPUT16), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT16), .ZN(new_n317));
  INV_X1    g131(.A(G125), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n317), .B1(new_n318), .B2(G140), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n316), .A2(new_n190), .A3(new_n319), .ZN(new_n320));
  OR2_X1    g134(.A1(new_n320), .A2(KEYINPUT75), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n316), .A2(new_n319), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G146), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n320), .A2(KEYINPUT75), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n321), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G128), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G119), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT72), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT23), .ZN(new_n330));
  INV_X1    g144(.A(G119), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G128), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT23), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n327), .A2(new_n328), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n330), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT73), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n330), .A2(new_n334), .A3(KEYINPUT73), .A4(new_n332), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n337), .A2(G110), .A3(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n327), .A2(new_n332), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  XOR2_X1   g155(.A(KEYINPUT24), .B(G110), .Z(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n325), .B(new_n339), .C1(new_n341), .C2(new_n343), .ZN(new_n344));
  OAI22_X1  g158(.A1(new_n335), .A2(G110), .B1(new_n340), .B2(new_n342), .ZN(new_n345));
  XNOR2_X1  g159(.A(G125), .B(G140), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n190), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(new_n323), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT22), .B(G137), .ZN(new_n350));
  INV_X1    g164(.A(G953), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(G221), .A3(G234), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n350), .B(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n344), .A2(new_n348), .A3(new_n353), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n271), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT25), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT25), .A4(new_n271), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n311), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  AND2_X1   g175(.A1(new_n355), .A2(new_n356), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n311), .A2(new_n271), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(KEYINPUT76), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n197), .A2(new_n318), .ZN(new_n368));
  OAI211_X1 g182(.A(G125), .B(new_n230), .C1(new_n232), .C2(new_n235), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n351), .A2(G224), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT7), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n374), .B(KEYINPUT82), .ZN(new_n375));
  XOR2_X1   g189(.A(G116), .B(G119), .Z(new_n376));
  INV_X1    g190(.A(KEYINPUT5), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n331), .A3(G116), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G113), .ZN(new_n380));
  OAI22_X1  g194(.A1(new_n378), .A2(new_n380), .B1(new_n376), .B2(new_n247), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n382));
  INV_X1    g196(.A(G104), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n382), .B1(new_n383), .B2(G107), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(G107), .ZN(new_n385));
  INV_X1    g199(.A(G107), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(KEYINPUT80), .A3(G104), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n385), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G101), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT3), .B1(new_n383), .B2(G107), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT3), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(new_n386), .A3(G104), .ZN(new_n392));
  INV_X1    g206(.A(G101), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n390), .A2(new_n392), .A3(new_n393), .A4(new_n385), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n381), .B(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(G110), .B(G122), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(KEYINPUT8), .ZN(new_n398));
  AOI22_X1  g212(.A1(new_n396), .A2(new_n398), .B1(new_n370), .B2(new_n373), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n375), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT78), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n390), .A2(new_n392), .A3(new_n385), .ZN(new_n402));
  AND2_X1   g216(.A1(new_n402), .A2(G101), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n394), .A2(KEYINPUT4), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n401), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(G101), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n406), .A2(KEYINPUT78), .A3(KEYINPUT4), .A4(new_n394), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n402), .A2(new_n409), .A3(G101), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT79), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT79), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n402), .A2(new_n412), .A3(new_n409), .A4(G101), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n248), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n381), .A2(new_n395), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n397), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n271), .B1(new_n400), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n418), .A2(new_n419), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT6), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n416), .B1(new_n408), .B2(new_n414), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n423), .B1(new_n424), .B2(new_n397), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n418), .A2(new_n423), .A3(new_n419), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n370), .B(new_n371), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT81), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT81), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n426), .A2(new_n431), .A3(new_n427), .A4(new_n428), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n421), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(G210), .B1(G237), .B2(G902), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n434), .B(KEYINPUT83), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n435), .B1(new_n437), .B2(new_n433), .ZN(new_n438));
  INV_X1    g252(.A(G469), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT12), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n395), .B(new_n197), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n440), .B1(new_n441), .B2(new_n229), .ZN(new_n442));
  INV_X1    g256(.A(new_n196), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n188), .A2(G128), .B1(new_n191), .B2(new_n192), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n395), .B(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n240), .A2(new_n446), .A3(KEYINPUT12), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(G110), .B(G140), .ZN(new_n449));
  INV_X1    g263(.A(G227), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(G953), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n449), .B(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n236), .B1(new_n411), .B2(new_n413), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT10), .B1(new_n395), .B2(new_n445), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT10), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n197), .A2(new_n455), .A3(new_n394), .A4(new_n389), .ZN(new_n456));
  AOI22_X1  g270(.A1(new_n408), .A2(new_n453), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n452), .B1(new_n457), .B2(new_n229), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n448), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n452), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n408), .A2(new_n453), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n454), .A2(new_n456), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n240), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n457), .A2(new_n229), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n439), .B(new_n271), .C1(new_n459), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(G469), .A2(G902), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n458), .A2(new_n464), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n442), .A2(new_n447), .B1(new_n457), .B2(new_n229), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n469), .B(G469), .C1(new_n460), .C2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n467), .A2(new_n468), .A3(new_n471), .ZN(new_n472));
  XOR2_X1   g286(.A(KEYINPUT9), .B(G234), .Z(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT77), .ZN(new_n474));
  OAI21_X1  g288(.A(G221), .B1(new_n474), .B2(G902), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  XOR2_X1   g290(.A(G113), .B(G122), .Z(new_n477));
  XOR2_X1   g291(.A(KEYINPUT86), .B(G104), .Z(new_n478));
  XOR2_X1   g292(.A(new_n477), .B(new_n478), .Z(new_n479));
  AND2_X1   g293(.A1(new_n314), .A2(new_n315), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT19), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT19), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n346), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n314), .A2(new_n315), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT85), .B1(new_n485), .B2(new_n483), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(G146), .ZN(new_n488));
  INV_X1    g302(.A(G237), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(new_n351), .A3(G214), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(new_n187), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n254), .A2(G143), .A3(G214), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G131), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n491), .A2(new_n219), .A3(new_n492), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n323), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n488), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT84), .ZN(new_n499));
  NAND2_X1  g313(.A1(KEYINPUT18), .A2(G131), .ZN(new_n500));
  OR3_X1    g314(.A1(new_n493), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n500), .B1(new_n493), .B2(new_n499), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n480), .A2(G146), .ZN(new_n503));
  AOI22_X1  g317(.A1(new_n501), .A2(new_n502), .B1(new_n347), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n479), .B1(new_n498), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n501), .A2(new_n502), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n503), .A2(new_n347), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n479), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n493), .A2(KEYINPUT17), .A3(G131), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(new_n496), .B2(KEYINPUT17), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n508), .B(new_n509), .C1(new_n325), .C2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n505), .A2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT20), .ZN(new_n514));
  NOR2_X1   g328(.A1(G475), .A2(G902), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT87), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n513), .A2(KEYINPUT87), .A3(new_n514), .A4(new_n515), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n513), .A2(new_n515), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT20), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  OR2_X1    g336(.A1(new_n511), .A2(new_n325), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n509), .B1(new_n523), .B2(new_n508), .ZN(new_n524));
  INV_X1    g338(.A(new_n512), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n271), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G475), .ZN(new_n527));
  NAND2_X1  g341(.A1(G234), .A2(G237), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(G952), .A3(new_n351), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(G902), .A3(G953), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  XNOR2_X1  g346(.A(KEYINPUT21), .B(G898), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n187), .A2(G128), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n326), .A2(KEYINPUT89), .A3(G143), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT89), .B1(new_n326), .B2(G143), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n211), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n214), .B(new_n536), .C1(new_n537), .C2(new_n538), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(G116), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(G122), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT88), .B(G122), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n544), .B1(new_n545), .B2(new_n543), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT14), .B1(new_n545), .B2(new_n543), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n547), .A3(G107), .ZN(new_n548));
  OAI221_X1 g362(.A(new_n544), .B1(KEYINPUT14), .B2(new_n386), .C1(new_n545), .C2(new_n543), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n542), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  OR2_X1    g364(.A1(new_n541), .A2(KEYINPUT91), .ZN(new_n551));
  OR2_X1    g365(.A1(new_n546), .A2(new_n386), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n541), .A2(KEYINPUT91), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n546), .A2(new_n386), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n551), .A2(new_n552), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT13), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n536), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n187), .A2(KEYINPUT13), .A3(G128), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n557), .B(new_n558), .C1(new_n537), .C2(new_n538), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n559), .A2(KEYINPUT90), .A3(G134), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT90), .B1(new_n559), .B2(G134), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n550), .B1(new_n555), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n351), .A2(G217), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n474), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n565), .B(new_n550), .C1(new_n555), .C2(new_n562), .ZN(new_n568));
  AOI21_X1  g382(.A(G902), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(G478), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(KEYINPUT15), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  AOI211_X1 g387(.A(G902), .B(new_n571), .C1(new_n567), .C2(new_n568), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n522), .A2(new_n527), .A3(new_n535), .A4(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n476), .A2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(G214), .B1(G237), .B2(G902), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n438), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n308), .A2(new_n367), .A3(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(G101), .ZN(G3));
  NOR2_X1   g396(.A1(new_n284), .A2(new_n289), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n296), .B1(new_n583), .B2(KEYINPUT31), .ZN(new_n584));
  OAI21_X1  g398(.A(G472), .B1(new_n584), .B2(G902), .ZN(new_n585));
  INV_X1    g399(.A(new_n476), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n585), .A2(new_n297), .A3(new_n367), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n567), .A2(new_n568), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n566), .A2(KEYINPUT33), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT33), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n588), .A2(KEYINPUT92), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n591), .B1(new_n588), .B2(KEYINPUT92), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n570), .A2(G902), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  OAI22_X1  g410(.A1(new_n594), .A2(new_n596), .B1(G478), .B2(new_n569), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n522), .A2(new_n527), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n598), .A2(new_n599), .A3(new_n534), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n433), .A2(new_n434), .ZN(new_n602));
  INV_X1    g416(.A(new_n434), .ZN(new_n603));
  AOI211_X1 g417(.A(new_n603), .B(new_n421), .C1(new_n430), .C2(new_n432), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n578), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n587), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(KEYINPUT93), .ZN(new_n607));
  XNOR2_X1  g421(.A(KEYINPUT34), .B(G104), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G6));
  INV_X1    g423(.A(new_n578), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n430), .A2(new_n432), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n603), .B1(new_n611), .B2(new_n421), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n610), .B1(new_n612), .B2(new_n435), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n521), .A2(new_n516), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n527), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n534), .B(KEYINPUT94), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NOR3_X1   g431(.A1(new_n615), .A2(new_n575), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n587), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT35), .B(G107), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G9));
  NAND2_X1  g436(.A1(new_n585), .A2(new_n297), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n354), .A2(KEYINPUT36), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n349), .B(new_n624), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n625), .A2(new_n365), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n361), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n438), .A2(new_n577), .A3(new_n578), .A4(new_n628), .ZN(new_n629));
  OR2_X1    g443(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(KEYINPUT37), .B(G110), .Z(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G12));
  NOR2_X1   g446(.A1(new_n476), .A2(new_n627), .ZN(new_n633));
  INV_X1    g447(.A(G900), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n532), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n529), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR3_X1   g451(.A1(new_n615), .A2(new_n575), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n613), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n308), .A2(new_n633), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G128), .ZN(G30));
  XNOR2_X1  g456(.A(new_n636), .B(KEYINPUT39), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n586), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n644), .A2(KEYINPUT40), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n644), .A2(KEYINPUT40), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n599), .A2(new_n575), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(new_n578), .A3(new_n627), .ZN(new_n648));
  NOR3_X1   g462(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n297), .A2(KEYINPUT32), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n306), .A2(new_n299), .A3(new_n280), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n583), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n267), .B1(new_n251), .B2(new_n262), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n271), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(G472), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n438), .B(new_n658), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n649), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(new_n187), .ZN(G45));
  NAND2_X1  g475(.A1(new_n522), .A2(new_n527), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n597), .A2(new_n662), .A3(new_n636), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n663), .B(new_n578), .C1(new_n604), .C2(new_n602), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n308), .A2(new_n633), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT96), .B(G146), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G48));
  INV_X1    g482(.A(new_n367), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n669), .B1(new_n652), .B2(new_n279), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n439), .A2(KEYINPUT97), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n464), .A2(new_n465), .ZN(new_n672));
  AOI22_X1  g486(.A1(new_n672), .A2(new_n452), .B1(new_n448), .B2(new_n458), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n671), .B1(new_n673), .B2(G902), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n457), .A2(new_n229), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n461), .A2(new_n229), .A3(new_n462), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n452), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n448), .A2(new_n458), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n671), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n679), .A2(new_n271), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n674), .A2(new_n681), .A3(new_n475), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT98), .ZN(new_n683));
  NOR3_X1   g497(.A1(new_n601), .A2(new_n683), .A3(new_n605), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n670), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT41), .B(G113), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT99), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n685), .B(new_n687), .ZN(G15));
  INV_X1    g502(.A(KEYINPUT100), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT98), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n682), .B(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n613), .A3(new_n618), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n689), .B1(new_n670), .B2(new_n693), .ZN(new_n694));
  AOI22_X1  g508(.A1(new_n650), .A2(new_n651), .B1(new_n278), .B2(G472), .ZN(new_n695));
  NOR4_X1   g509(.A1(new_n695), .A2(new_n692), .A3(KEYINPUT100), .A4(new_n669), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(new_n543), .ZN(G18));
  INV_X1    g512(.A(KEYINPUT101), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n699), .B1(new_n683), .B2(new_n605), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n691), .A2(new_n613), .A3(KEYINPUT101), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n627), .A2(new_n576), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n308), .A2(new_n700), .A3(new_n701), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G119), .ZN(G21));
  OAI211_X1 g518(.A(new_n647), .B(new_n578), .C1(new_n602), .C2(new_n604), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n705), .A2(new_n683), .A3(new_n617), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT102), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n707), .B1(new_n584), .B2(G902), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n302), .A2(new_n305), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n280), .B1(new_n709), .B2(new_n271), .ZN(new_n710));
  AOI211_X1 g524(.A(G472), .B(G902), .C1(new_n302), .C2(new_n305), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n708), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n707), .B(new_n280), .C1(new_n584), .C2(G902), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n706), .A2(new_n367), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G122), .ZN(G24));
  NAND4_X1  g529(.A1(new_n712), .A2(new_n628), .A3(new_n663), .A4(new_n713), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n700), .A2(new_n701), .ZN(new_n717));
  OR2_X1    g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G125), .ZN(G27));
  INV_X1    g533(.A(KEYINPUT104), .ZN(new_n720));
  INV_X1    g534(.A(new_n475), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n721), .B1(new_n472), .B2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n467), .A2(KEYINPUT103), .A3(new_n468), .A4(new_n471), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n720), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n435), .B(new_n578), .C1(new_n437), .C2(new_n433), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n723), .A2(new_n720), .A3(new_n724), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT105), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n472), .A2(new_n722), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n730), .A2(new_n475), .A3(new_n724), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(KEYINPUT104), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n433), .A2(new_n437), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n733), .A2(new_n604), .A3(new_n610), .ZN(new_n734));
  AND4_X1   g548(.A1(KEYINPUT105), .A2(new_n732), .A3(new_n734), .A4(new_n728), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n670), .B(new_n663), .C1(new_n729), .C2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT42), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n732), .A2(new_n734), .A3(new_n728), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT105), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n727), .A2(KEYINPUT105), .A3(new_n728), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(KEYINPUT42), .A3(new_n670), .A4(new_n663), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n738), .A2(KEYINPUT106), .A3(new_n744), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT106), .B1(new_n738), .B2(new_n744), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G131), .ZN(G33));
  XNOR2_X1  g562(.A(new_n638), .B(KEYINPUT107), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n670), .B(new_n749), .C1(new_n729), .C2(new_n735), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G134), .ZN(G36));
  OR2_X1    g565(.A1(new_n470), .A2(new_n460), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(KEYINPUT45), .A3(new_n469), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n753), .A2(KEYINPUT108), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(KEYINPUT108), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT45), .B1(new_n752), .B2(new_n469), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n439), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n468), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT46), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n758), .A2(KEYINPUT46), .A3(new_n468), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(new_n467), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n475), .A3(new_n643), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n598), .A2(new_n662), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT43), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n766), .B1(new_n662), .B2(KEYINPUT109), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n765), .B(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n768), .A2(new_n623), .A3(new_n628), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT44), .ZN(new_n770));
  AOI211_X1 g584(.A(new_n726), .B(new_n764), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n771), .B1(new_n770), .B2(new_n769), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G137), .ZN(G39));
  AND3_X1   g587(.A1(new_n763), .A2(KEYINPUT47), .A3(new_n475), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT47), .B1(new_n763), .B2(new_n475), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n695), .A2(new_n669), .A3(new_n663), .A4(new_n734), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G140), .ZN(G42));
  NOR3_X1   g593(.A1(new_n669), .A2(new_n610), .A3(new_n721), .ZN(new_n780));
  INV_X1    g594(.A(new_n674), .ZN(new_n781));
  INV_X1    g595(.A(new_n681), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n784), .A2(KEYINPUT49), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n780), .A2(new_n785), .A3(new_n765), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT110), .ZN(new_n787));
  INV_X1    g601(.A(new_n659), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n788), .B1(KEYINPUT49), .B2(new_n784), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n787), .A2(new_n789), .A3(new_n657), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT111), .ZN(new_n791));
  AND4_X1   g605(.A1(new_n628), .A2(new_n712), .A3(new_n663), .A4(new_n713), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n743), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n575), .A2(new_n636), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n726), .A2(new_n615), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n308), .A2(new_n633), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n793), .A2(new_n750), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n714), .A2(new_n685), .A3(new_n703), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n797), .A2(new_n697), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n738), .A2(new_n744), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT106), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n738), .A2(KEYINPUT106), .A3(new_n744), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n662), .A2(new_n575), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n438), .A2(new_n578), .A3(new_n616), .A4(new_n804), .ZN(new_n805));
  OAI22_X1  g619(.A1(new_n587), .A2(new_n805), .B1(new_n623), .B2(new_n629), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT113), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n808));
  OAI221_X1 g622(.A(new_n808), .B1(new_n623), .B2(new_n629), .C1(new_n587), .C2(new_n805), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n695), .A2(new_n669), .A3(new_n579), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n598), .A2(new_n599), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(new_n438), .A3(new_n578), .A4(new_n616), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n587), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT112), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT112), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n581), .B(new_n816), .C1(new_n587), .C2(new_n813), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n810), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n799), .A2(new_n802), .A3(new_n803), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT114), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n308), .B(new_n633), .C1(new_n640), .C2(new_n665), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT115), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n823), .B1(new_n628), .B2(new_n637), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n627), .A2(KEYINPUT115), .A3(new_n636), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n731), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n657), .A2(new_n613), .A3(new_n647), .A4(new_n826), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n822), .B(new_n827), .C1(new_n717), .C2(new_n716), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n718), .A2(KEYINPUT52), .A3(new_n822), .A4(new_n827), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n830), .A2(KEYINPUT116), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT116), .B1(new_n830), .B2(new_n831), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n832), .A2(new_n833), .A3(KEYINPUT53), .ZN(new_n834));
  INV_X1    g648(.A(new_n798), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n308), .A2(new_n367), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT100), .B1(new_n836), .B2(new_n692), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n670), .A2(new_n689), .A3(new_n693), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n840), .A2(new_n818), .A3(new_n797), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n841), .A2(new_n747), .A3(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n821), .A2(new_n834), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n830), .A2(new_n831), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n841), .A2(new_n747), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT53), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n844), .A2(KEYINPUT54), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n849));
  INV_X1    g663(.A(new_n845), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n849), .B1(new_n820), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n845), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n830), .A2(KEYINPUT116), .A3(new_n831), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n849), .B1(new_n738), .B2(new_n744), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n841), .A2(new_n854), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n851), .A2(new_n852), .A3(new_n857), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n848), .A2(KEYINPUT117), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT117), .B1(new_n848), .B2(new_n858), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n768), .A2(new_n530), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n683), .A2(new_n726), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n863), .A2(new_n836), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n864), .B(KEYINPUT48), .Z(new_n865));
  INV_X1    g679(.A(G952), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n862), .A2(new_n367), .A3(new_n530), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(new_n657), .ZN(new_n868));
  AOI211_X1 g682(.A(new_n866), .B(G953), .C1(new_n868), .C2(new_n812), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n712), .A2(new_n713), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n870), .A2(new_n367), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n861), .ZN(new_n872));
  OAI211_X1 g686(.A(new_n865), .B(new_n869), .C1(new_n717), .C2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n788), .A2(new_n610), .A3(new_n691), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT50), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n870), .A2(new_n628), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n863), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n868), .A2(new_n599), .A3(new_n598), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n871), .A2(new_n734), .A3(new_n861), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n783), .A2(new_n721), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n882), .B1(new_n776), .B2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT51), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n873), .B1(new_n881), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n776), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n888), .A2(KEYINPUT118), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n883), .B(KEYINPUT119), .Z(new_n890));
  AOI21_X1  g704(.A(new_n890), .B1(new_n888), .B2(KEYINPUT118), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n882), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n885), .B1(new_n880), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n887), .A2(new_n893), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n859), .A2(new_n860), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(G952), .A2(G953), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n791), .B1(new_n895), .B2(new_n896), .ZN(G75));
  NAND2_X1  g711(.A1(new_n866), .A2(G953), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT123), .Z(new_n899));
  NAND2_X1  g713(.A1(new_n851), .A2(new_n857), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(G902), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT56), .B1(new_n902), .B2(G210), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n426), .A2(new_n427), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(new_n428), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT55), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n899), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n907), .A2(KEYINPUT122), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(KEYINPUT122), .ZN(new_n910));
  XOR2_X1   g724(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n911));
  NAND3_X1  g725(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n902), .A2(KEYINPUT120), .A3(new_n436), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n914), .B1(new_n901), .B2(new_n437), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n912), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n908), .A2(new_n916), .ZN(G51));
  INV_X1    g731(.A(new_n899), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n468), .B(KEYINPUT57), .Z(new_n919));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n851), .A2(new_n920), .A3(new_n852), .A4(new_n857), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n832), .A2(new_n833), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n799), .A2(new_n819), .A3(new_n856), .ZN(new_n923));
  AOI22_X1  g737(.A1(new_n846), .A2(new_n849), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n921), .B1(new_n852), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n920), .B1(new_n924), .B2(new_n852), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n919), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n679), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n901), .A2(new_n758), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n918), .B1(new_n928), .B2(new_n929), .ZN(G54));
  NAND2_X1  g744(.A1(KEYINPUT58), .A2(G475), .ZN(new_n931));
  OR3_X1    g745(.A1(new_n901), .A2(new_n513), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n513), .B1(new_n901), .B2(new_n931), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n918), .B1(new_n932), .B2(new_n933), .ZN(G60));
  NAND2_X1  g748(.A1(G478), .A2(G902), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT59), .Z(new_n936));
  NOR2_X1   g750(.A1(new_n594), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(new_n925), .B2(new_n926), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n899), .ZN(new_n939));
  INV_X1    g753(.A(new_n936), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(new_n859), .B2(new_n860), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n939), .B1(new_n594), .B2(new_n941), .ZN(G63));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n943));
  XNOR2_X1  g757(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n944));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n924), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n625), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n899), .B1(new_n947), .B2(new_n362), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n943), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OR2_X1    g765(.A1(new_n947), .A2(new_n362), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n952), .A2(KEYINPUT61), .A3(new_n899), .A4(new_n948), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(new_n953), .ZN(G66));
  NAND2_X1  g768(.A1(G224), .A2(G953), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n533), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n840), .A2(new_n818), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n956), .B1(new_n957), .B2(new_n351), .ZN(new_n958));
  INV_X1    g772(.A(G898), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n904), .B1(new_n959), .B2(G953), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n958), .B(new_n960), .Z(G69));
  NAND2_X1  g775(.A1(new_n772), .A2(new_n778), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n764), .A2(new_n836), .A3(new_n705), .ZN(new_n963));
  INV_X1    g777(.A(new_n750), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n718), .A2(new_n822), .ZN(new_n965));
  NOR4_X1   g779(.A1(new_n962), .A2(new_n963), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n966), .A2(new_n351), .A3(new_n747), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n245), .B(new_n487), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(G900), .B2(G953), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n967), .A2(KEYINPUT127), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(KEYINPUT127), .B1(new_n967), .B2(new_n969), .ZN(new_n971));
  INV_X1    g785(.A(new_n968), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n812), .A2(new_n804), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n973), .A2(new_n644), .A3(new_n726), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n962), .B1(new_n670), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(KEYINPUT62), .B1(new_n965), .B2(new_n660), .ZN(new_n976));
  OR3_X1    g790(.A1(new_n965), .A2(KEYINPUT62), .A3(new_n660), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n972), .B1(new_n978), .B2(new_n351), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n970), .A2(new_n971), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g794(.A(G953), .B1(new_n450), .B2(new_n634), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n967), .A2(new_n969), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(KEYINPUT126), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  OAI22_X1  g798(.A1(new_n980), .A2(new_n981), .B1(new_n982), .B2(new_n984), .ZN(G72));
  NAND2_X1  g799(.A1(G472), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT63), .Z(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n978), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n988), .B1(new_n989), .B2(new_n957), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n252), .A2(new_n267), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n899), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n844), .A2(new_n847), .ZN(new_n993));
  AOI211_X1 g807(.A(new_n988), .B(new_n993), .C1(new_n259), .C2(new_n583), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n966), .A2(new_n747), .A3(new_n957), .ZN(new_n995));
  AOI211_X1 g809(.A(new_n267), .B(new_n252), .C1(new_n995), .C2(new_n987), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n992), .A2(new_n994), .A3(new_n996), .ZN(G57));
endmodule


