//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n205), .B(new_n206), .Z(new_n207));
  NAND2_X1  g006(.A1(G229gat), .A2(G233gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(KEYINPUT14), .B(G29gat), .ZN(new_n210));
  INV_X1    g009(.A(G36gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G43gat), .B(G50gat), .ZN(new_n213));
  INV_X1    g012(.A(G29gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n212), .A2(KEYINPUT15), .A3(new_n213), .A4(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n216), .A2(KEYINPUT84), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(KEYINPUT84), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n212), .A2(new_n215), .ZN(new_n220));
  XOR2_X1   g019(.A(new_n213), .B(KEYINPUT15), .Z(new_n221));
  AOI22_X1  g020(.A1(new_n218), .A2(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT16), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n223), .B1(new_n224), .B2(G1gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G1gat), .B2(new_n223), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(G8gat), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n222), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT85), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n222), .A2(new_n230), .A3(KEYINPUT17), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n221), .A2(new_n220), .ZN(new_n232));
  INV_X1    g031(.A(new_n219), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n232), .B1(new_n233), .B2(new_n217), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT17), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT85), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n227), .B1(new_n234), .B2(new_n235), .ZN(new_n238));
  AOI211_X1 g037(.A(new_n209), .B(new_n229), .C1(new_n237), .C2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT18), .B1(new_n239), .B2(KEYINPUT86), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n234), .B(new_n227), .ZN(new_n241));
  XOR2_X1   g040(.A(new_n208), .B(KEYINPUT13), .Z(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n229), .B1(new_n237), .B2(new_n238), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(new_n208), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT86), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT18), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n246), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n207), .B1(new_n244), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n207), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n240), .A2(new_n249), .A3(new_n252), .A4(new_n243), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(G197gat), .ZN(new_n255));
  INV_X1    g054(.A(G204gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G197gat), .A2(G204gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT22), .ZN(new_n259));
  NAND2_X1  g058(.A1(G211gat), .A2(G218gat), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n257), .A2(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(G211gat), .B(G218gat), .Z(new_n262));
  OR3_X1    g061(.A1(new_n261), .A2(new_n262), .A3(KEYINPUT70), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n262), .B1(new_n261), .B2(KEYINPUT70), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT25), .ZN(new_n267));
  INV_X1    g066(.A(G169gat), .ZN(new_n268));
  INV_X1    g067(.A(G176gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT23), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT24), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n271), .A2(G183gat), .A3(G190gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT24), .ZN(new_n274));
  NOR2_X1   g073(.A1(G183gat), .A2(G190gat), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n270), .B(new_n272), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G169gat), .A2(G176gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n277), .B1(new_n278), .B2(KEYINPUT23), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n267), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n273), .ZN(new_n281));
  AOI22_X1  g080(.A1(new_n281), .A2(new_n271), .B1(new_n278), .B2(KEYINPUT23), .ZN(new_n282));
  NAND3_X1  g081(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n268), .A2(new_n269), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT23), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n267), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G183gat), .ZN(new_n290));
  INV_X1    g089(.A(G190gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n292), .A2(KEYINPUT24), .A3(new_n273), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n282), .A2(new_n286), .A3(new_n289), .A4(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n280), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n290), .A2(KEYINPUT27), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT27), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G183gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(new_n298), .A3(new_n291), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT28), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(KEYINPUT27), .B(G183gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n302), .A2(KEYINPUT28), .A3(new_n291), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n305));
  AND2_X1   g104(.A1(new_n305), .A2(new_n277), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT26), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n278), .A2(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n281), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G226gat), .ZN(new_n312));
  INV_X1    g111(.A(G233gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n314), .B1(new_n311), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n266), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n280), .A2(new_n294), .B1(new_n304), .B2(new_n309), .ZN(new_n320));
  OAI22_X1  g119(.A1(new_n320), .A2(KEYINPUT29), .B1(new_n312), .B2(new_n313), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n321), .A2(new_n265), .A3(new_n315), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  XOR2_X1   g122(.A(G8gat), .B(G36gat), .Z(new_n324));
  XOR2_X1   g123(.A(G64gat), .B(G92gat), .Z(new_n325));
  XOR2_X1   g124(.A(new_n324), .B(new_n325), .Z(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(KEYINPUT71), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n326), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n329), .B1(new_n319), .B2(new_n322), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT30), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  OR2_X1    g130(.A1(new_n330), .A2(KEYINPUT30), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(G225gat), .A2(G233gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT73), .ZN(new_n337));
  AND2_X1   g136(.A1(G141gat), .A2(G148gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(G141gat), .A2(G148gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(G141gat), .ZN(new_n341));
  INV_X1    g140(.A(G148gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G141gat), .A2(G148gat), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n343), .A2(KEYINPUT73), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT2), .ZN(new_n347));
  INV_X1    g146(.A(G155gat), .ZN(new_n348));
  INV_X1    g147(.A(G162gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n340), .A2(new_n345), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(G155gat), .B(G162gat), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n338), .A2(new_n339), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT72), .B(KEYINPUT2), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT74), .B1(new_n351), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n350), .A2(new_n346), .ZN(new_n357));
  NOR3_X1   g156(.A1(new_n338), .A2(new_n339), .A3(new_n337), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT73), .B1(new_n343), .B2(new_n344), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT74), .ZN(new_n361));
  XOR2_X1   g160(.A(G155gat), .B(G162gat), .Z(new_n362));
  XOR2_X1   g161(.A(KEYINPUT72), .B(KEYINPUT2), .Z(new_n363));
  NAND2_X1  g162(.A1(new_n343), .A2(new_n344), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n360), .A2(new_n361), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n356), .A2(new_n366), .A3(KEYINPUT3), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n340), .A2(new_n345), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n354), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n368), .A2(new_n357), .B1(new_n369), .B2(new_n362), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT3), .ZN(new_n371));
  INV_X1    g170(.A(G120gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G113gat), .ZN(new_n373));
  INV_X1    g172(.A(G113gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G120gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT1), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G127gat), .B(G134gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n373), .A2(new_n375), .A3(KEYINPUT65), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT65), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n383), .A2(new_n374), .A3(G120gat), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n382), .A2(new_n377), .A3(new_n379), .A4(new_n384), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n370), .A2(new_n371), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  AOI211_X1 g185(.A(KEYINPUT5), .B(new_n336), .C1(new_n367), .C2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(G134gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n388), .A2(G127gat), .ZN(new_n389));
  INV_X1    g188(.A(G127gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(G134gat), .ZN(new_n391));
  AND4_X1   g190(.A1(new_n377), .A2(new_n384), .A3(new_n389), .A4(new_n391), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n392), .A2(new_n382), .B1(new_n378), .B2(new_n380), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT4), .B1(new_n393), .B2(new_n370), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT75), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n360), .A2(new_n365), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n385), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n395), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n393), .A2(new_n370), .A3(KEYINPUT75), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n394), .B1(new_n400), .B2(KEYINPUT4), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n387), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n398), .A2(new_n403), .A3(new_n399), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n367), .A2(new_n386), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n393), .A2(new_n370), .A3(KEYINPUT4), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n404), .A2(new_n405), .A3(new_n335), .A4(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT5), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n356), .A2(new_n366), .A3(new_n397), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT76), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT76), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n356), .A2(new_n366), .A3(new_n411), .A4(new_n397), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n400), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n335), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n402), .B1(new_n408), .B2(new_n415), .ZN(new_n416));
  XOR2_X1   g215(.A(G1gat), .B(G29gat), .Z(new_n417));
  XNOR2_X1  g216(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n418));
  XNOR2_X1  g217(.A(new_n417), .B(new_n418), .ZN(new_n419));
  XNOR2_X1  g218(.A(G57gat), .B(G85gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n400), .B1(new_n410), .B2(new_n412), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n407), .B(KEYINPUT5), .C1(new_n423), .C2(new_n335), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n421), .B1(new_n387), .B2(new_n401), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT6), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n422), .A2(KEYINPUT81), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n421), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n428), .B1(new_n424), .B2(new_n402), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT6), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT81), .B1(new_n422), .B2(new_n426), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n334), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT82), .ZN(new_n434));
  AND2_X1   g233(.A1(G169gat), .A2(G176gat), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n435), .B1(new_n287), .B2(new_n288), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n282), .A2(new_n436), .A3(new_n293), .ZN(new_n437));
  INV_X1    g236(.A(new_n276), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT64), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n277), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n283), .ZN(new_n441));
  OAI21_X1  g240(.A(KEYINPUT25), .B1(new_n278), .B2(KEYINPUT23), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n267), .A2(new_n437), .B1(new_n438), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n308), .A2(new_n277), .A3(new_n305), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n273), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n446), .B1(new_n301), .B2(new_n303), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n397), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(G227gat), .A2(G233gat), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n295), .A2(new_n310), .A3(new_n393), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n449), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT34), .B1(new_n452), .B2(KEYINPUT69), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n451), .B(new_n453), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n295), .A2(new_n393), .A3(new_n310), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n393), .B1(new_n295), .B2(new_n310), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n452), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  XOR2_X1   g256(.A(G71gat), .B(G99gat), .Z(new_n458));
  XNOR2_X1  g257(.A(G15gat), .B(G43gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(new_n458), .B(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT33), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n457), .A2(KEYINPUT32), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT67), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n457), .A2(KEYINPUT67), .A3(KEYINPUT32), .A4(new_n461), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n457), .A2(KEYINPUT32), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT33), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n457), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n467), .A2(new_n469), .A3(KEYINPUT66), .A4(new_n460), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT66), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n449), .B1(new_n448), .B2(new_n450), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n460), .B1(new_n472), .B2(KEYINPUT33), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT32), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n471), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  AND4_X1   g275(.A1(new_n454), .A2(new_n466), .A3(new_n470), .A4(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(KEYINPUT31), .B(G50gat), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n317), .B1(new_n396), .B2(KEYINPUT3), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(new_n265), .ZN(new_n481));
  NAND2_X1  g280(.A1(G228gat), .A2(G233gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT79), .ZN(new_n484));
  AND2_X1   g283(.A1(new_n257), .A2(new_n258), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n261), .A2(KEYINPUT79), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n262), .A3(new_n488), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n489), .B(new_n317), .C1(new_n262), .C2(new_n487), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n370), .B1(new_n490), .B2(new_n371), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n483), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n371), .B1(new_n265), .B2(KEYINPUT29), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n356), .A2(new_n366), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n482), .B1(new_n495), .B2(new_n481), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n479), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n479), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n493), .A2(new_n494), .B1(new_n480), .B2(new_n265), .ZN(new_n499));
  OAI221_X1 g298(.A(new_n498), .B1(new_n483), .B2(new_n491), .C1(new_n499), .C2(new_n482), .ZN(new_n500));
  XNOR2_X1  g299(.A(G78gat), .B(G106gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(G22gat), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n497), .A2(new_n500), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n502), .B1(new_n497), .B2(new_n500), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n466), .A2(new_n470), .A3(new_n476), .ZN(new_n506));
  INV_X1    g305(.A(new_n454), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT35), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n478), .A2(new_n505), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT82), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n512), .B(new_n334), .C1(new_n431), .C2(new_n432), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n434), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT68), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n454), .B1(new_n506), .B2(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n466), .A2(new_n476), .A3(KEYINPUT68), .A4(new_n470), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n477), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT78), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n422), .B1(new_n426), .B2(new_n519), .ZN(new_n520));
  AOI211_X1 g319(.A(KEYINPUT78), .B(KEYINPUT6), .C1(new_n424), .C2(new_n425), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n430), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n518), .A2(new_n505), .A3(new_n522), .A4(new_n334), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT35), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n514), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n506), .A2(new_n515), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n526), .A2(new_n507), .A3(new_n517), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n527), .A2(KEYINPUT36), .A3(new_n478), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT36), .ZN(new_n529));
  INV_X1    g328(.A(new_n508), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n529), .B1(new_n530), .B2(new_n477), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n505), .ZN(new_n533));
  INV_X1    g332(.A(new_n430), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n424), .A2(new_n425), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT6), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n429), .B1(new_n537), .B2(KEYINPUT78), .ZN(new_n538));
  INV_X1    g337(.A(new_n521), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n534), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n533), .B1(new_n540), .B2(new_n333), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT38), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT37), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n326), .B1(new_n323), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n319), .A2(KEYINPUT37), .A3(new_n322), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n321), .A2(new_n265), .A3(new_n315), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n265), .B1(new_n321), .B2(new_n315), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n543), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n327), .A2(KEYINPUT38), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n549), .A2(new_n545), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n330), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n546), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT81), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n537), .B2(new_n429), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n554), .A2(new_n556), .A3(new_n430), .A4(new_n427), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n429), .B1(new_n331), .B2(new_n332), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT39), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n401), .A2(new_n405), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n559), .B1(new_n560), .B2(new_n336), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n423), .A2(KEYINPUT80), .A3(new_n335), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n423), .A2(new_n335), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT80), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n561), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT40), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n335), .B1(new_n401), .B2(new_n405), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n421), .B1(new_n568), .B2(new_n559), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n567), .B1(new_n566), .B2(new_n569), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n558), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n557), .A2(new_n572), .A3(new_n505), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n532), .A2(new_n541), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n254), .B1(new_n525), .B2(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(KEYINPUT91), .B(KEYINPUT19), .Z(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT92), .ZN(new_n577));
  XOR2_X1   g376(.A(G127gat), .B(G155gat), .Z(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G183gat), .B(G211gat), .Z(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT20), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT87), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(G71gat), .B(G78gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(G64gat), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n589), .A2(G57gat), .ZN(new_n590));
  XOR2_X1   g389(.A(KEYINPUT89), .B(G57gat), .Z(new_n591));
  AOI21_X1  g390(.A(new_n590), .B1(new_n591), .B2(G64gat), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT90), .ZN(new_n594));
  XOR2_X1   g393(.A(G57gat), .B(G64gat), .Z(new_n595));
  AOI21_X1  g394(.A(new_n587), .B1(new_n586), .B2(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n596), .B(KEYINPUT88), .Z(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT21), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n600), .A2(G231gat), .A3(G233gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n598), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n583), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n598), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n227), .B1(new_n606), .B2(KEYINPUT21), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n601), .A2(new_n583), .A3(new_n603), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n605), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n608), .B1(new_n605), .B2(new_n609), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n582), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n612), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n614), .A2(new_n610), .A3(new_n581), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g415(.A1(G232gat), .A2(G233gat), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n617), .A2(KEYINPUT41), .ZN(new_n618));
  XNOR2_X1  g417(.A(G134gat), .B(G162gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G190gat), .B(G218gat), .Z(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT94), .ZN(new_n624));
  NAND2_X1  g423(.A1(G85gat), .A2(G92gat), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n625), .A2(KEYINPUT93), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT7), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G99gat), .A2(G106gat), .ZN(new_n629));
  INV_X1    g428(.A(G85gat), .ZN(new_n630));
  INV_X1    g429(.A(G92gat), .ZN(new_n631));
  AOI22_X1  g430(.A1(KEYINPUT8), .A2(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(KEYINPUT7), .B1(new_n625), .B2(KEYINPUT93), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n628), .B(new_n632), .C1(new_n626), .C2(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(G99gat), .B(G106gat), .Z(new_n635));
  XOR2_X1   g434(.A(new_n634), .B(new_n635), .Z(new_n636));
  AOI21_X1  g435(.A(new_n636), .B1(new_n234), .B2(new_n235), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n624), .B1(new_n237), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n237), .A2(new_n624), .A3(new_n637), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n617), .A2(KEYINPUT41), .ZN(new_n642));
  INV_X1    g441(.A(new_n636), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n642), .B1(new_n643), .B2(new_n222), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n623), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  AOI211_X1 g445(.A(new_n622), .B(new_n644), .C1(new_n639), .C2(new_n640), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n621), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n640), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n645), .B1(new_n649), .B2(new_n638), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n622), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n641), .A2(new_n623), .A3(new_n645), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n651), .A2(new_n652), .A3(new_n620), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n648), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n616), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n598), .A2(new_n643), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT10), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n594), .A2(new_n597), .A3(new_n636), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n658), .A2(new_n657), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(G230gat), .A2(G233gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n662), .B1(new_n656), .B2(new_n658), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G120gat), .B(G148gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(G176gat), .B(G204gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n666), .B(new_n667), .Z(new_n668));
  NAND3_X1  g467(.A1(new_n663), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n668), .ZN(new_n670));
  INV_X1    g469(.A(new_n662), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n671), .B1(new_n659), .B2(new_n660), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n672), .B2(new_n664), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n655), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n575), .A2(new_n675), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n522), .A2(KEYINPUT95), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n522), .A2(KEYINPUT95), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT96), .B(G1gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1324gat));
  XNOR2_X1  g482(.A(KEYINPUT16), .B(G8gat), .ZN(new_n684));
  OR3_X1    g483(.A1(new_n676), .A2(new_n334), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n676), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n333), .ZN(new_n688));
  AOI22_X1  g487(.A1(new_n686), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n688), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n686), .A2(KEYINPUT97), .A3(KEYINPUT42), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT97), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT42), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n691), .B1(new_n685), .B2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n689), .B1(new_n690), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT98), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT98), .ZN(new_n696));
  OAI211_X1 g495(.A(new_n696), .B(new_n689), .C1(new_n690), .C2(new_n693), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(G1325gat));
  NAND2_X1  g497(.A1(new_n478), .A2(new_n508), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(G15gat), .B1(new_n687), .B2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT99), .ZN(new_n702));
  INV_X1    g501(.A(new_n532), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n703), .A2(G15gat), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n702), .B1(new_n687), .B2(new_n704), .ZN(G1326gat));
  NOR2_X1   g504(.A1(new_n676), .A2(new_n505), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT43), .B(G22gat), .Z(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  INV_X1    g507(.A(KEYINPUT100), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n616), .A2(new_n674), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n648), .A2(new_n653), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NOR4_X1   g511(.A1(new_n616), .A2(new_n654), .A3(KEYINPUT100), .A4(new_n674), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(new_n575), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n716), .A2(new_n214), .A3(new_n679), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT45), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT102), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(KEYINPUT44), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n510), .B1(new_n433), .B2(KEYINPUT82), .ZN(new_n721));
  AOI22_X1  g520(.A1(new_n721), .A2(new_n513), .B1(KEYINPUT35), .B2(new_n523), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n532), .A2(new_n541), .A3(new_n573), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n711), .B(new_n720), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n654), .B1(new_n525), .B2(new_n574), .ZN(new_n725));
  XNOR2_X1  g524(.A(KEYINPUT102), .B(KEYINPUT44), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n616), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n674), .B(KEYINPUT101), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n251), .A2(new_n253), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n728), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n727), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n734), .A2(KEYINPUT103), .A3(new_n679), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT103), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(new_n733), .B2(new_n680), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n735), .A2(G29gat), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n718), .A2(new_n738), .ZN(G1328gat));
  NOR3_X1   g538(.A1(new_n715), .A2(G36gat), .A3(new_n334), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT46), .ZN(new_n741));
  OAI21_X1  g540(.A(G36gat), .B1(new_n733), .B2(new_n334), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(G1329gat));
  NOR3_X1   g542(.A1(new_n715), .A2(G43gat), .A3(new_n699), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n727), .A2(new_n703), .A3(new_n732), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G43gat), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n745), .A2(KEYINPUT47), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n744), .B1(new_n747), .B2(KEYINPUT104), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT104), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n746), .A2(new_n750), .A3(G43gat), .ZN(new_n751));
  AOI211_X1 g550(.A(KEYINPUT105), .B(KEYINPUT47), .C1(new_n749), .C2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT105), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n711), .B1(new_n722), .B2(new_n723), .ZN(new_n754));
  INV_X1    g553(.A(new_n726), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI211_X1 g555(.A(new_n532), .B(new_n731), .C1(new_n756), .C2(new_n724), .ZN(new_n757));
  INV_X1    g556(.A(G43gat), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT104), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n759), .A2(new_n751), .A3(new_n745), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT47), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n753), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n748), .B1(new_n752), .B2(new_n762), .ZN(G1330gat));
  NOR3_X1   g562(.A1(new_n715), .A2(G50gat), .A3(new_n505), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n734), .A2(new_n533), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n764), .B1(new_n765), .B2(G50gat), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g566(.A(new_n729), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n254), .ZN(new_n769));
  AOI211_X1 g568(.A(new_n655), .B(new_n769), .C1(new_n574), .C2(new_n525), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n679), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(new_n591), .Z(G1332gat));
  INV_X1    g571(.A(KEYINPUT49), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n333), .B1(new_n773), .B2(new_n589), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT106), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n773), .A2(new_n589), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1333gat));
  NAND2_X1  g577(.A1(new_n770), .A2(new_n703), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n699), .A2(G71gat), .ZN(new_n780));
  AOI22_X1  g579(.A1(new_n779), .A2(G71gat), .B1(new_n770), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g581(.A1(new_n770), .A2(new_n533), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G78gat), .ZN(G1335gat));
  INV_X1    g583(.A(KEYINPUT108), .ZN(new_n785));
  OR3_X1    g584(.A1(new_n616), .A2(new_n730), .A3(KEYINPUT107), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT107), .B1(new_n616), .B2(new_n730), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n727), .A2(new_n674), .A3(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n785), .B1(new_n789), .B2(new_n680), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n674), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n791), .B1(new_n756), .B2(new_n724), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n792), .A2(KEYINPUT108), .A3(new_n679), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n790), .A2(G85gat), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n725), .A2(new_n788), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT51), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n725), .A2(KEYINPUT51), .A3(new_n788), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n679), .A2(new_n630), .A3(new_n674), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n794), .B1(new_n799), .B2(new_n800), .ZN(G1336gat));
  OAI21_X1  g600(.A(G92gat), .B1(new_n789), .B2(new_n334), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT110), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n729), .A2(G92gat), .A3(new_n334), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n802), .B(new_n803), .C1(new_n799), .C2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT109), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n807), .B1(new_n802), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n631), .B1(new_n792), .B2(new_n333), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n805), .B1(new_n797), .B2(new_n798), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT110), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n806), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n809), .B1(new_n806), .B2(new_n812), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n813), .A2(new_n814), .ZN(G1337gat));
  INV_X1    g614(.A(G99gat), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n792), .A2(new_n703), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n816), .B1(new_n817), .B2(KEYINPUT111), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(KEYINPUT111), .B2(new_n817), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n700), .A2(new_n816), .A3(new_n674), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(new_n799), .B2(new_n820), .ZN(G1338gat));
  OAI21_X1  g620(.A(G106gat), .B1(new_n789), .B2(new_n505), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n729), .A2(G106gat), .A3(new_n505), .ZN(new_n823));
  XOR2_X1   g622(.A(new_n823), .B(KEYINPUT112), .Z(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n799), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g625(.A1(new_n730), .A2(new_n374), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT116), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n659), .A2(new_n660), .A3(new_n671), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n663), .A2(KEYINPUT54), .A3(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n668), .B1(new_n672), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(KEYINPUT55), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n669), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT55), .B1(new_n830), .B2(new_n832), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n245), .A2(new_n208), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n241), .A2(new_n242), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n205), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n253), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n836), .A2(new_n711), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(KEYINPUT113), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT113), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n836), .A2(new_n711), .A3(new_n844), .A4(new_n841), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT114), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n674), .A2(new_n253), .A3(new_n839), .ZN(new_n848));
  AOI22_X1  g647(.A1(new_n836), .A2(new_n730), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n674), .A2(new_n253), .A3(KEYINPUT114), .A4(new_n839), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n711), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n728), .B1(new_n846), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n675), .A2(new_n254), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n505), .A3(new_n679), .ZN(new_n855));
  INV_X1    g654(.A(new_n518), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n855), .A2(new_n856), .A3(new_n333), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n857), .A2(KEYINPUT115), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n859));
  NOR4_X1   g658(.A1(new_n855), .A2(new_n859), .A3(new_n856), .A4(new_n333), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n828), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n655), .A2(new_n730), .A3(new_n674), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n848), .A2(new_n847), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n830), .A2(new_n832), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT55), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n669), .A3(new_n833), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n863), .B(new_n850), .C1(new_n254), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n654), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(new_n843), .A3(new_n845), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n862), .B1(new_n870), .B2(new_n728), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(new_n533), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n872), .A2(new_n700), .A3(new_n334), .A4(new_n679), .ZN(new_n873));
  OAI21_X1  g672(.A(G113gat), .B1(new_n873), .B2(new_n254), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n861), .A2(new_n874), .ZN(G1340gat));
  AOI21_X1  g674(.A(G120gat), .B1(new_n669), .B2(new_n673), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n876), .B1(new_n858), .B2(new_n860), .ZN(new_n877));
  OAI21_X1  g676(.A(G120gat), .B1(new_n873), .B2(new_n729), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(G1341gat));
  NAND3_X1  g678(.A1(new_n857), .A2(new_n390), .A3(new_n616), .ZN(new_n880));
  OAI21_X1  g679(.A(G127gat), .B1(new_n873), .B2(new_n728), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(G1342gat));
  NAND2_X1  g681(.A1(new_n711), .A2(new_n334), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(G134gat), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n872), .A2(new_n518), .A3(new_n679), .A4(new_n884), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n885), .A2(KEYINPUT56), .ZN(new_n886));
  OAI21_X1  g685(.A(G134gat), .B1(new_n873), .B2(new_n654), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(KEYINPUT56), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(G1343gat));
  NOR3_X1   g688(.A1(new_n680), .A2(new_n703), .A3(new_n333), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT57), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n892), .B1(new_n871), .B2(new_n505), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n505), .A2(new_n892), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n843), .A2(new_n845), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n848), .A2(KEYINPUT117), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n674), .A2(new_n253), .A3(new_n897), .A4(new_n839), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n896), .B(new_n898), .C1(new_n254), .C2(new_n867), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n654), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n616), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n894), .B1(new_n901), .B2(new_n862), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n891), .B1(new_n893), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n341), .B1(new_n903), .B2(new_n730), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT118), .B1(new_n703), .B2(new_n505), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT118), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n532), .A2(new_n906), .A3(new_n533), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n905), .A2(new_n679), .A3(new_n907), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n871), .A2(new_n333), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n341), .A3(new_n730), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT58), .B1(new_n904), .B2(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT58), .ZN(new_n913));
  AOI211_X1 g712(.A(new_n254), .B(new_n891), .C1(new_n893), .C2(new_n902), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n913), .B(new_n910), .C1(new_n914), .C2(new_n341), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n912), .A2(new_n915), .ZN(G1344gat));
  INV_X1    g715(.A(new_n894), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n917), .B1(new_n852), .B2(new_n853), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n867), .A2(new_n654), .A3(new_n840), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n919), .B1(new_n899), .B2(new_n654), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n853), .B1(new_n920), .B2(new_n616), .ZN(new_n921));
  AOI21_X1  g720(.A(KEYINPUT57), .B1(new_n921), .B2(new_n533), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n674), .A3(new_n890), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT59), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n903), .A2(new_n926), .A3(new_n674), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n926), .B1(new_n909), .B2(new_n674), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n925), .B(new_n927), .C1(G148gat), .C2(new_n928), .ZN(G1345gat));
  NOR2_X1   g728(.A1(new_n728), .A2(new_n348), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT57), .B1(new_n854), .B2(new_n533), .ZN(new_n931));
  INV_X1    g730(.A(new_n900), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n728), .B1(new_n932), .B2(new_n846), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n917), .B1(new_n933), .B2(new_n853), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n890), .B(new_n930), .C1(new_n931), .C2(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n908), .B1(new_n852), .B2(new_n853), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT119), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n936), .A2(new_n937), .A3(new_n334), .A4(new_n616), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(new_n348), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n937), .B1(new_n909), .B2(new_n616), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n935), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT120), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT120), .ZN(new_n943));
  OAI211_X1 g742(.A(new_n935), .B(new_n943), .C1(new_n939), .C2(new_n940), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(G1346gat));
  NOR4_X1   g744(.A1(new_n871), .A2(G162gat), .A3(new_n883), .A4(new_n908), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT121), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n903), .A2(new_n711), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n948), .B2(new_n349), .ZN(G1347gat));
  NOR2_X1   g748(.A1(new_n871), .A2(new_n679), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n518), .A2(new_n505), .A3(new_n333), .ZN(new_n951));
  XNOR2_X1  g750(.A(new_n951), .B(KEYINPUT122), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n953), .A2(new_n268), .A3(new_n730), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n680), .A2(new_n333), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n955), .A2(new_n699), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n872), .A2(new_n730), .A3(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n957), .A2(new_n958), .A3(G169gat), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n958), .B1(new_n957), .B2(G169gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n954), .B1(new_n959), .B2(new_n960), .ZN(G1348gat));
  AND2_X1   g760(.A1(new_n872), .A2(new_n956), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n729), .A2(new_n269), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n962), .A2(KEYINPUT124), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g763(.A(G176gat), .B1(new_n953), .B2(new_n674), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT124), .B1(new_n962), .B2(new_n963), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(G1349gat));
  NAND2_X1  g766(.A1(new_n872), .A2(new_n956), .ZN(new_n968));
  OAI21_X1  g767(.A(G183gat), .B1(new_n968), .B2(new_n728), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n950), .A2(new_n302), .A3(new_n616), .A4(new_n952), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(KEYINPUT60), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT60), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n969), .A2(new_n973), .A3(new_n970), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n974), .ZN(G1350gat));
  NAND3_X1  g774(.A1(new_n953), .A2(new_n291), .A3(new_n711), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n872), .A2(new_n711), .A3(new_n956), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT61), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n977), .A2(new_n978), .A3(G190gat), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n978), .B1(new_n977), .B2(G190gat), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n976), .B1(new_n979), .B2(new_n980), .ZN(G1351gat));
  NOR3_X1   g780(.A1(new_n703), .A2(new_n505), .A3(new_n334), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n950), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g782(.A(G197gat), .B1(new_n983), .B2(new_n730), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n955), .A2(new_n703), .ZN(new_n985));
  AND2_X1   g784(.A1(new_n923), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n254), .A2(new_n255), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(G1352gat));
  NAND3_X1  g787(.A1(new_n983), .A2(new_n256), .A3(new_n674), .ZN(new_n989));
  XNOR2_X1  g788(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n923), .A2(new_n768), .A3(new_n985), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(G204gat), .ZN(new_n993));
  AND2_X1   g792(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n994));
  OAI211_X1 g793(.A(new_n991), .B(new_n993), .C1(new_n994), .C2(new_n989), .ZN(G1353gat));
  OAI211_X1 g794(.A(new_n616), .B(new_n985), .C1(new_n918), .C2(new_n922), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(G211gat), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT63), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n996), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n999), .A2(KEYINPUT126), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g800(.A(KEYINPUT63), .B1(new_n996), .B2(G211gat), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT126), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n728), .A2(G211gat), .ZN(new_n1004));
  AOI22_X1  g803(.A1(new_n1002), .A2(new_n1003), .B1(new_n983), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1001), .A2(new_n1005), .ZN(G1354gat));
  AOI21_X1  g805(.A(G218gat), .B1(new_n983), .B2(new_n711), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n711), .A2(G218gat), .ZN(new_n1008));
  XNOR2_X1  g807(.A(new_n1008), .B(KEYINPUT127), .ZN(new_n1009));
  AOI21_X1  g808(.A(new_n1007), .B1(new_n986), .B2(new_n1009), .ZN(G1355gat));
endmodule


