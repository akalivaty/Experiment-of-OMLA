//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1241, new_n1242, new_n1243,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n206));
  INV_X1    g0006(.A(G68), .ZN(new_n207));
  INV_X1    g0007(.A(G238), .ZN(new_n208));
  INV_X1    g0008(.A(G77), .ZN(new_n209));
  INV_X1    g0009(.A(G244), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(KEYINPUT66), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n214));
  NAND3_X1  g0014(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n211), .A2(KEYINPUT66), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n205), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT67), .ZN(new_n218));
  INV_X1    g0018(.A(KEYINPUT1), .ZN(new_n219));
  OR2_X1    g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n218), .A2(new_n219), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n205), .A2(G13), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT64), .Z(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT0), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n229), .A2(G50), .A3(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n225), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  AND3_X1   g0033(.A1(new_n220), .A2(new_n221), .A3(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT68), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n238), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G58), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(G107), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G97), .ZN(new_n249));
  INV_X1    g0049(.A(G97), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G107), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G87), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n247), .B(new_n254), .ZN(G351));
  OR2_X1    g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G1698), .ZN(new_n259));
  INV_X1    g0059(.A(G223), .ZN(new_n260));
  OAI22_X1  g0060(.A1(new_n259), .A2(new_n260), .B1(new_n209), .B2(new_n258), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT72), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT72), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G1698), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n263), .B(new_n265), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G222), .ZN(new_n269));
  OR3_X1    g0069(.A1(new_n268), .A2(KEYINPUT73), .A3(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(KEYINPUT73), .B1(new_n268), .B2(new_n269), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n261), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(new_n226), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  OR2_X1    g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G179), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT69), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT69), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G41), .ZN(new_n281));
  INV_X1    g0081(.A(G45), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n279), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT70), .B1(new_n273), .B2(new_n226), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G33), .A2(G41), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT70), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n285), .A2(new_n286), .A3(G1), .A4(G13), .ZN(new_n287));
  INV_X1    g0087(.A(G274), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(G1), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n283), .A2(new_n284), .A3(new_n287), .A4(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G1), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(G41), .B2(G45), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n284), .A2(new_n287), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT71), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT71), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n284), .A2(new_n295), .A3(new_n287), .A4(new_n292), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G226), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n276), .A2(new_n277), .A3(new_n290), .A4(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G50), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n227), .B1(new_n201), .B2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT75), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n301), .B(new_n302), .ZN(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT8), .B(G58), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G33), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n306), .A2(G20), .ZN(new_n307));
  NOR2_X1   g0107(.A1(G20), .A2(G33), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n305), .A2(new_n307), .B1(G150), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT74), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g0113(.A1(KEYINPUT74), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(new_n226), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G13), .ZN(new_n316));
  NOR3_X1   g0116(.A1(new_n316), .A2(new_n227), .A3(G1), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n310), .A2(new_n315), .B1(new_n300), .B2(new_n317), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n315), .A2(new_n317), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n291), .A2(G20), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(G50), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G169), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n290), .B1(new_n272), .B2(new_n275), .ZN(new_n324));
  INV_X1    g0124(.A(new_n298), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n323), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n299), .A2(new_n322), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n276), .A2(G190), .A3(new_n290), .A4(new_n298), .ZN(new_n329));
  AOI21_X1  g0129(.A(KEYINPUT9), .B1(new_n318), .B2(new_n321), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(G200), .B1(new_n324), .B2(new_n325), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n318), .A2(KEYINPUT9), .A3(new_n321), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n329), .A2(new_n331), .A3(new_n332), .A4(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT10), .ZN(new_n335));
  INV_X1    g0135(.A(new_n333), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n336), .A2(new_n330), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT10), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n337), .A2(new_n338), .A3(new_n329), .A4(new_n332), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n328), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n284), .A2(G232), .A3(new_n287), .A4(new_n292), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n290), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g0142(.A(G226), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G33), .A2(G87), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n343), .B(new_n344), .C1(new_n268), .C2(new_n260), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n274), .ZN(new_n346));
  INV_X1    g0146(.A(G190), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n342), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n290), .A2(new_n341), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(new_n274), .B2(new_n345), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n348), .B1(new_n350), .B2(G200), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n304), .B1(new_n291), .B2(G20), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n319), .A2(new_n352), .B1(new_n317), .B2(new_n304), .ZN(new_n353));
  INV_X1    g0153(.A(G58), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n354), .A2(new_n207), .ZN(new_n355));
  OAI21_X1  g0155(.A(G20), .B1(new_n355), .B2(new_n201), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n308), .A2(G159), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n266), .A2(new_n267), .ZN(new_n359));
  AOI21_X1  g0159(.A(KEYINPUT7), .B1(new_n359), .B2(new_n227), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT7), .ZN(new_n361));
  NOR4_X1   g0161(.A1(new_n266), .A2(new_n267), .A3(new_n361), .A4(G20), .ZN(new_n362));
  OAI21_X1  g0162(.A(G68), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT82), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n358), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n256), .A2(new_n227), .A3(new_n257), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n361), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n256), .A2(KEYINPUT7), .A3(new_n227), .A4(new_n257), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n207), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT82), .ZN(new_n370));
  AOI21_X1  g0170(.A(KEYINPUT16), .B1(new_n365), .B2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n358), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n363), .A2(KEYINPUT16), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n315), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n351), .B(new_n353), .C1(new_n371), .C2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT17), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n353), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT16), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n372), .B1(new_n369), .B2(KEYINPUT82), .ZN(new_n380));
  AOI211_X1 g0180(.A(new_n364), .B(new_n207), .C1(new_n367), .C2(new_n368), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n313), .A2(new_n226), .A3(new_n314), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n369), .A2(new_n358), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n383), .B1(new_n384), .B2(KEYINPUT16), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n378), .B1(new_n382), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n342), .A2(new_n346), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G169), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n342), .A2(new_n346), .A3(G179), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g0190(.A(KEYINPUT18), .B1(new_n386), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n353), .B1(new_n371), .B2(new_n374), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT18), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n388), .A2(new_n389), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n386), .A2(KEYINPUT17), .A3(new_n351), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n377), .A2(new_n391), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n359), .A2(G107), .ZN(new_n399));
  OAI221_X1 g0199(.A(new_n399), .B1(new_n268), .B2(new_n240), .C1(new_n259), .C2(new_n208), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n290), .B1(new_n401), .B2(new_n275), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n210), .B1(new_n294), .B2(new_n296), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(G190), .ZN(new_n405));
  XOR2_X1   g0205(.A(KEYINPUT15), .B(G87), .Z(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n307), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n227), .A2(new_n209), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n407), .B1(KEYINPUT77), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n304), .B(KEYINPUT76), .ZN(new_n410));
  INV_X1    g0210(.A(new_n308), .ZN(new_n411));
  OAI221_X1 g0211(.A(new_n409), .B1(KEYINPUT77), .B2(new_n407), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n315), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n319), .A2(G77), .A3(new_n320), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n317), .A2(new_n209), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(G200), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n405), .B(new_n416), .C1(new_n404), .C2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n404), .A2(new_n277), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n323), .B1(new_n402), .B2(new_n403), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AND2_X1   g0222(.A1(new_n418), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n340), .A2(new_n398), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n290), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n263), .A2(new_n265), .A3(G226), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G232), .A2(G1698), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n258), .ZN(new_n429));
  AND3_X1   g0229(.A1(KEYINPUT78), .A2(G33), .A3(G97), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT78), .B1(G33), .B2(G97), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n425), .B1(new_n433), .B2(new_n274), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n297), .A2(G238), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT13), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n432), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n438), .B1(new_n428), .B2(new_n258), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n290), .B1(new_n439), .B2(new_n275), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n208), .B1(new_n294), .B2(new_n296), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT13), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G169), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT14), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT80), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n434), .A2(new_n435), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(KEYINPUT80), .B1(new_n440), .B2(new_n441), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT13), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n449), .A2(G179), .A3(new_n437), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT14), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n443), .A2(new_n451), .A3(G169), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n445), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n308), .A2(G50), .B1(G20), .B2(new_n207), .ZN(new_n454));
  INV_X1    g0254(.A(new_n307), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n454), .B1(new_n455), .B2(new_n209), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n315), .ZN(new_n457));
  XNOR2_X1  g0257(.A(new_n457), .B(KEYINPUT81), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT11), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT81), .ZN(new_n461));
  XNOR2_X1  g0261(.A(new_n457), .B(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT11), .ZN(new_n463));
  INV_X1    g0263(.A(new_n317), .ZN(new_n464));
  OR3_X1    g0264(.A1(new_n464), .A2(KEYINPUT12), .A3(G68), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT12), .B1(new_n464), .B2(G68), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n207), .B1(new_n291), .B2(G20), .ZN(new_n467));
  AOI22_X1  g0267(.A1(new_n465), .A2(new_n466), .B1(new_n319), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n460), .A2(new_n463), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n453), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n469), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n449), .A2(G190), .A3(new_n437), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT79), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n473), .B1(new_n443), .B2(G200), .ZN(new_n474));
  AOI211_X1 g0274(.A(KEYINPUT79), .B(new_n417), .C1(new_n437), .C2(new_n442), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n471), .B(new_n472), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n424), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n288), .B1(KEYINPUT5), .B2(new_n278), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n284), .A2(new_n287), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT84), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT5), .B1(new_n279), .B2(new_n281), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n282), .A2(G1), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n481), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  XNOR2_X1  g0285(.A(KEYINPUT69), .B(G41), .ZN(new_n486));
  OAI211_X1 g0286(.A(KEYINPUT84), .B(new_n483), .C1(new_n486), .C2(KEYINPUT5), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n480), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  OAI211_X1 g0288(.A(G264), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n256), .A2(G303), .A3(new_n257), .ZN(new_n490));
  OAI21_X1  g0290(.A(G257), .B1(new_n266), .B2(new_n267), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n263), .A2(new_n265), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n489), .B(new_n490), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n493), .A2(new_n274), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n284), .A2(new_n287), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n278), .A2(KEYINPUT5), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n483), .B(new_n496), .C1(new_n486), .C2(KEYINPUT5), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n497), .A3(G270), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n488), .A2(new_n494), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n291), .A2(G33), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n383), .A2(G116), .A3(new_n464), .A4(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(G116), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n317), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(G20), .B1(G33), .B2(G283), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n306), .A2(G97), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n504), .A2(new_n505), .B1(G20), .B2(new_n502), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n315), .A2(KEYINPUT20), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT20), .B1(new_n315), .B2(new_n506), .ZN(new_n508));
  OAI211_X1 g0308(.A(new_n501), .B(new_n503), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n499), .A2(new_n509), .A3(G169), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT21), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT90), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n510), .A2(KEYINPUT90), .A3(new_n511), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n499), .A2(KEYINPUT21), .A3(G169), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n488), .A2(new_n494), .A3(new_n498), .A4(G179), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(new_n509), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n509), .B1(new_n499), .B2(G200), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n347), .B2(new_n499), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n516), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n464), .A2(new_n406), .ZN(new_n525));
  AOI21_X1  g0325(.A(G20), .B1(new_n256), .B2(new_n257), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G68), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT19), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n455), .B2(new_n250), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(G87), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT87), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT87), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G87), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n533), .A2(new_n535), .A3(new_n250), .A4(new_n248), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G97), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT78), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(KEYINPUT78), .A2(G33), .A3(G97), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n528), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(KEYINPUT88), .B(new_n536), .C1(new_n541), .C2(G20), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(KEYINPUT19), .B1(new_n430), .B2(new_n431), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n227), .ZN(new_n545));
  AOI21_X1  g0345(.A(KEYINPUT88), .B1(new_n545), .B2(new_n536), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n531), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n525), .B1(new_n547), .B2(new_n315), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G116), .ZN(new_n549));
  OAI211_X1 g0349(.A(G244), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n549), .B(new_n550), .C1(new_n268), .C2(new_n208), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n289), .A2(G45), .ZN(new_n552));
  INV_X1    g0352(.A(G250), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n552), .B1(new_n553), .B2(new_n483), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n551), .A2(new_n274), .B1(new_n495), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n347), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n556), .B1(G200), .B2(new_n555), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n319), .A2(new_n500), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(new_n532), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n548), .A2(new_n557), .A3(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n551), .A2(new_n274), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n495), .A2(new_n554), .ZN(new_n563));
  AOI21_X1  g0363(.A(G169), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n277), .B2(new_n555), .ZN(new_n565));
  INV_X1    g0365(.A(new_n525), .ZN(new_n566));
  AND2_X1   g0366(.A1(new_n319), .A2(new_n500), .ZN(new_n567));
  XNOR2_X1  g0367(.A(KEYINPUT15), .B(G87), .ZN(new_n568));
  XNOR2_X1  g0368(.A(new_n568), .B(KEYINPUT89), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n536), .B1(new_n541), .B2(G20), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT88), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n530), .B1(new_n573), .B2(new_n542), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n566), .B(new_n570), .C1(new_n574), .C2(new_n383), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n565), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n561), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n495), .A2(new_n497), .A3(G257), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n488), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT4), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n268), .B2(new_n210), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT83), .ZN(new_n582));
  XNOR2_X1  g0382(.A(KEYINPUT72), .B(G1698), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n258), .A2(new_n583), .A3(G244), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT83), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n585), .A3(new_n580), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n258), .A2(new_n583), .A3(KEYINPUT4), .A4(G244), .ZN(new_n587));
  INV_X1    g0387(.A(G283), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n306), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n359), .A2(new_n262), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n589), .B1(new_n590), .B2(G250), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n582), .A2(new_n586), .A3(new_n587), .A4(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n579), .B1(new_n592), .B2(new_n274), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G190), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT6), .ZN(new_n595));
  NOR3_X1   g0395(.A1(new_n595), .A2(new_n250), .A3(G107), .ZN(new_n596));
  XNOR2_X1  g0396(.A(G97), .B(G107), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n596), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  OAI22_X1  g0398(.A1(new_n598), .A2(new_n227), .B1(new_n209), .B2(new_n411), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n248), .B1(new_n367), .B2(new_n368), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n315), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n567), .A2(G97), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n464), .A2(G97), .ZN(new_n603));
  INV_X1    g0403(.A(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n601), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n579), .A2(KEYINPUT85), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT85), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n488), .A2(new_n607), .A3(new_n578), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n606), .A2(new_n608), .B1(new_n274), .B2(new_n592), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n594), .B(new_n605), .C1(new_n609), .C2(new_n417), .ZN(new_n610));
  INV_X1    g0410(.A(new_n589), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n587), .B(new_n611), .C1(new_n553), .C2(new_n259), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n585), .B1(new_n584), .B2(new_n580), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n275), .B1(new_n614), .B2(new_n586), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n323), .B1(new_n615), .B2(new_n579), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n601), .A2(new_n602), .A3(new_n604), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n592), .A2(new_n274), .ZN(new_n618));
  INV_X1    g0418(.A(new_n608), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n607), .B1(new_n488), .B2(new_n578), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n618), .B(new_n277), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n616), .A2(new_n617), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n610), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n577), .B1(new_n623), .B2(KEYINPUT86), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n317), .A2(new_n248), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT25), .ZN(new_n626));
  XNOR2_X1  g0426(.A(new_n625), .B(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(new_n558), .B2(new_n248), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT23), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n227), .B2(G107), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n248), .A2(KEYINPUT23), .A3(G20), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n227), .A2(G33), .A3(G116), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT22), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n526), .B2(G87), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n227), .B(G87), .C1(new_n266), .C2(new_n267), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n638), .A2(KEYINPUT22), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n635), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT24), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n638), .A2(KEYINPUT22), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n258), .A2(new_n636), .A3(new_n227), .A4(G87), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT24), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n644), .A2(new_n645), .A3(new_n635), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n628), .B1(new_n647), .B2(new_n315), .ZN(new_n648));
  OAI211_X1 g0448(.A(G257), .B(G1698), .C1(new_n266), .C2(new_n267), .ZN(new_n649));
  NAND2_X1  g0449(.A1(G33), .A2(G294), .ZN(new_n650));
  OAI211_X1 g0450(.A(new_n649), .B(new_n650), .C1(new_n268), .C2(new_n553), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n274), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n495), .A2(new_n497), .A3(G264), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n488), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n323), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n488), .A2(new_n652), .A3(new_n277), .A4(new_n653), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT91), .B1(new_n648), .B2(new_n657), .ZN(new_n658));
  AOI211_X1 g0458(.A(KEYINPUT24), .B(new_n634), .C1(new_n642), .C2(new_n643), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n645), .B1(new_n644), .B2(new_n635), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n315), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n628), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT91), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n663), .A2(new_n664), .A3(new_n656), .A4(new_n655), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n654), .A2(new_n347), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n654), .A2(G200), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n648), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n658), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n579), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n618), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n605), .B1(new_n323), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(G200), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n617), .B1(new_n593), .B2(G190), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n672), .A2(new_n621), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT86), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n669), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  AND4_X1   g0478(.A1(new_n478), .A2(new_n524), .A3(new_n624), .A4(new_n678), .ZN(G372));
  NAND2_X1  g0479(.A1(new_n335), .A2(new_n339), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n377), .A2(new_n396), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n476), .A2(new_n420), .A3(new_n419), .A4(new_n421), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n681), .B1(new_n682), .B2(new_n470), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n391), .A2(new_n395), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n680), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AND2_X1   g0485(.A1(new_n685), .A2(new_n327), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n610), .A2(new_n622), .A3(new_n668), .ZN(new_n687));
  AOI211_X1 g0487(.A(new_n525), .B(new_n559), .C1(new_n547), .C2(new_n315), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n688), .A2(new_n557), .B1(new_n575), .B2(new_n565), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n383), .B1(new_n641), .B2(new_n646), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n656), .B(new_n655), .C1(new_n690), .C2(new_n628), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n510), .A2(KEYINPUT90), .A3(new_n511), .ZN(new_n692));
  AOI21_X1  g0492(.A(KEYINPUT90), .B1(new_n510), .B2(new_n511), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n520), .B(new_n691), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n687), .A2(KEYINPUT92), .A3(new_n689), .A4(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT92), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n689), .A2(new_n610), .A3(new_n622), .A4(new_n668), .ZN(new_n697));
  INV_X1    g0497(.A(new_n694), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n576), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT26), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n622), .B2(new_n577), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n689), .A2(KEYINPUT26), .A3(new_n621), .A4(new_n672), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n700), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n695), .A2(new_n699), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n478), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n686), .A2(new_n706), .ZN(G369));
  AND2_X1   g0507(.A1(new_n516), .A2(new_n520), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n291), .A2(new_n227), .A3(G13), .ZN(new_n709));
  OR2_X1    g0509(.A1(new_n709), .A2(KEYINPUT27), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(KEYINPUT27), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n710), .A2(G213), .A3(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(G343), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n509), .A2(new_n714), .ZN(new_n715));
  MUX2_X1   g0515(.A(new_n708), .B(new_n523), .S(new_n715), .Z(new_n716));
  XNOR2_X1  g0516(.A(new_n716), .B(KEYINPUT93), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G330), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n669), .ZN(new_n720));
  INV_X1    g0520(.A(new_n714), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n720), .B1(new_n648), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(new_n691), .B2(new_n721), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  OR2_X1    g0524(.A1(new_n691), .A2(new_n714), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n708), .A2(new_n714), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n720), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(G399));
  INV_X1    g0528(.A(new_n486), .ZN(new_n729));
  INV_X1    g0529(.A(new_n222), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n536), .A2(G116), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n732), .A2(G1), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(new_n231), .B2(new_n732), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT28), .ZN(new_n736));
  INV_X1    g0536(.A(G330), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n678), .A2(new_n624), .A3(new_n524), .A4(new_n721), .ZN(new_n738));
  INV_X1    g0538(.A(new_n518), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n555), .A2(new_n653), .A3(new_n652), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n593), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT30), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n593), .A2(new_n739), .A3(new_n740), .A4(KEYINPUT30), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n555), .A2(G179), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n745), .A2(new_n654), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n673), .A2(new_n746), .A3(new_n499), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n743), .A2(new_n744), .A3(new_n747), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n748), .A2(KEYINPUT31), .A3(new_n714), .ZN(new_n749));
  AOI21_X1  g0549(.A(KEYINPUT31), .B1(new_n748), .B2(new_n714), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n737), .B1(new_n738), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n705), .A2(new_n721), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT29), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n516), .A2(new_n520), .A3(new_n658), .A4(new_n665), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n687), .A2(new_n689), .A3(new_n756), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n754), .B(new_n714), .C1(new_n704), .C2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n752), .B1(new_n755), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n736), .B1(new_n760), .B2(G1), .ZN(G364));
  AOI21_X1  g0561(.A(new_n226), .B1(G20), .B2(new_n323), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n227), .A2(new_n277), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G190), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT32), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n227), .A2(G179), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G190), .A2(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(G159), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n767), .A2(new_n207), .B1(new_n768), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(new_n768), .B2(new_n773), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n764), .A2(G190), .A3(new_n417), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n258), .B1(new_n776), .B2(new_n354), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n764), .A2(new_n770), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n777), .B1(G77), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n769), .A2(G190), .A3(G200), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(new_n533), .B2(new_n535), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n347), .A2(G179), .A3(G200), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n227), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n782), .B1(G97), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n769), .A2(new_n347), .A3(G200), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n248), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n765), .A2(new_n347), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n788), .B1(G50), .B2(new_n789), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n775), .A2(new_n780), .A3(new_n786), .A4(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n776), .ZN(new_n792));
  INV_X1    g0592(.A(new_n771), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n792), .A2(G322), .B1(new_n793), .B2(G329), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n258), .B1(new_n779), .B2(G311), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n789), .A2(G326), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT33), .B(G317), .ZN(new_n798));
  INV_X1    g0598(.A(new_n781), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n766), .A2(new_n798), .B1(new_n799), .B2(G303), .ZN(new_n800));
  INV_X1    g0600(.A(new_n787), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n785), .A2(G294), .B1(new_n801), .B2(G283), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n796), .A2(new_n797), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n763), .B1(new_n791), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(G13), .A2(G33), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n806), .A2(G20), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n762), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n730), .A2(new_n258), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n811), .B1(new_n232), .B2(new_n282), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n282), .B2(new_n247), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n258), .A2(new_n222), .ZN(new_n814));
  INV_X1    g0614(.A(G355), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n814), .A2(new_n815), .B1(G116), .B2(new_n222), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT94), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n809), .B1(new_n813), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n316), .A2(G20), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n291), .B1(new_n819), .B2(G45), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n732), .A2(new_n820), .ZN(new_n821));
  NOR3_X1   g0621(.A1(new_n804), .A2(new_n818), .A3(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n807), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n822), .B1(new_n717), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n718), .A2(new_n821), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n717), .A2(G330), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n824), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g0627(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n827), .B(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(G396));
  NAND2_X1  g0630(.A1(new_n420), .A2(new_n714), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n418), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n422), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n422), .A2(new_n714), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n753), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n835), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n705), .A2(new_n837), .A3(new_n721), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n752), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(new_n732), .B2(new_n820), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n836), .A2(new_n752), .A3(new_n838), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n792), .A2(G143), .B1(new_n779), .B2(G159), .ZN(new_n843));
  INV_X1    g0643(.A(G150), .ZN(new_n844));
  INV_X1    g0644(.A(G137), .ZN(new_n845));
  INV_X1    g0645(.A(new_n789), .ZN(new_n846));
  OAI221_X1 g0646(.A(new_n843), .B1(new_n767), .B2(new_n844), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT34), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(G132), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n258), .B1(new_n771), .B2(new_n850), .C1(new_n207), .C2(new_n787), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n784), .A2(new_n354), .B1(new_n781), .B2(new_n300), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n849), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n848), .B2(new_n847), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n787), .A2(new_n532), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n781), .A2(new_n248), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n855), .B(new_n856), .C1(G303), .C2(new_n789), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n258), .B1(new_n792), .B2(G294), .ZN(new_n858));
  AOI22_X1  g0658(.A1(G116), .A2(new_n779), .B1(new_n793), .B2(G311), .ZN(new_n859));
  AOI22_X1  g0659(.A1(G97), .A2(new_n785), .B1(new_n766), .B2(G283), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n857), .A2(new_n858), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n763), .B1(new_n854), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n762), .A2(new_n805), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n821), .B(new_n862), .C1(new_n209), .C2(new_n863), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT97), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n806), .B2(new_n837), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n842), .A2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(G384));
  INV_X1    g0668(.A(new_n598), .ZN(new_n869));
  OR2_X1    g0669(.A1(new_n869), .A2(KEYINPUT35), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(KEYINPUT35), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n870), .A2(new_n871), .A3(G116), .A4(new_n228), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT36), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n231), .A2(new_n209), .A3(new_n355), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT98), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n874), .A2(new_n875), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n300), .A2(G68), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT99), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n316), .A2(G1), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT40), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n738), .A2(new_n751), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n474), .A2(new_n475), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n472), .A2(new_n471), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n469), .B(new_n714), .C1(new_n886), .C2(new_n453), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n469), .A2(new_n714), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n470), .A2(new_n476), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n835), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n379), .B1(new_n369), .B2(new_n358), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(new_n373), .A3(new_n315), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n712), .B1(new_n892), .B2(new_n353), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n397), .A2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT100), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n392), .A2(new_n394), .ZN(new_n896));
  INV_X1    g0696(.A(new_n712), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n392), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT37), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n896), .A2(new_n898), .A3(new_n899), .A4(new_n375), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n892), .A2(new_n353), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n901), .B1(new_n394), .B2(new_n897), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n375), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT37), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n894), .A2(new_n895), .A3(KEYINPUT38), .A4(new_n905), .ZN(new_n906));
  AOI22_X1  g0706(.A1(new_n397), .A2(new_n893), .B1(new_n900), .B2(new_n904), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n906), .B1(KEYINPUT38), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n895), .B1(new_n907), .B2(KEYINPUT38), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n883), .B(new_n890), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n887), .A2(new_n889), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n883), .A2(new_n837), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n896), .A2(new_n898), .A3(new_n375), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(KEYINPUT37), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n900), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n397), .A2(new_n392), .A3(new_n897), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g0717(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n905), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n882), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n882), .A2(new_n910), .B1(new_n912), .B2(new_n921), .ZN(new_n922));
  AND3_X1   g0722(.A1(new_n922), .A2(new_n478), .A3(new_n883), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n922), .B1(new_n478), .B2(new_n883), .ZN(new_n924));
  OR3_X1    g0724(.A1(new_n923), .A2(new_n924), .A3(new_n737), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n887), .A2(new_n889), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n838), .B2(new_n834), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n909), .B2(new_n908), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n920), .A2(KEYINPUT100), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n894), .A2(new_n905), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT38), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n929), .A2(new_n932), .A3(KEYINPUT39), .A4(new_n906), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT39), .ZN(new_n934));
  INV_X1    g0734(.A(new_n920), .ZN(new_n935));
  INV_X1    g0735(.A(new_n918), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n936), .B1(new_n915), .B2(new_n916), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n934), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n470), .A2(new_n714), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n933), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n684), .A2(new_n712), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n928), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n755), .A2(new_n478), .A3(new_n759), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n686), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n942), .B(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n925), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n291), .B2(new_n819), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n925), .A2(new_n945), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n873), .B1(new_n880), .B2(new_n881), .C1(new_n947), .C2(new_n948), .ZN(G367));
  NOR2_X1   g0749(.A1(new_n688), .A2(new_n721), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n700), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n577), .B2(new_n950), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n952), .A2(KEYINPUT102), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n952), .A2(KEYINPUT102), .ZN(new_n954));
  NOR3_X1   g0754(.A1(new_n953), .A2(new_n954), .A3(KEYINPUT43), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(KEYINPUT43), .B2(new_n952), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n676), .B1(new_n605), .B2(new_n721), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n672), .A2(new_n621), .A3(new_n714), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OR3_X1    g0759(.A1(new_n959), .A2(new_n727), .A3(KEYINPUT42), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n658), .A2(new_n665), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n622), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n721), .ZN(new_n963));
  OAI21_X1  g0763(.A(KEYINPUT42), .B1(new_n959), .B2(new_n727), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n960), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT103), .ZN(new_n966));
  MUX2_X1   g0766(.A(new_n955), .B(new_n956), .S(new_n966), .Z(new_n967));
  OR2_X1    g0767(.A1(new_n724), .A2(new_n959), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n967), .A2(new_n968), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n731), .B(KEYINPUT41), .Z(new_n971));
  INV_X1    g0771(.A(new_n724), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n727), .A2(new_n725), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n959), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n974), .B(KEYINPUT44), .Z(new_n975));
  NOR2_X1   g0775(.A1(new_n973), .A2(new_n959), .ZN(new_n976));
  XNOR2_X1  g0776(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n976), .B(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n972), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n724), .A2(new_n975), .A3(new_n978), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n727), .B1(new_n723), .B2(new_n726), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n718), .B(new_n983), .Z(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n760), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n971), .B1(new_n986), .B2(new_n760), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n820), .B(KEYINPUT105), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  OAI211_X1 g0789(.A(new_n969), .B(new_n970), .C1(new_n987), .C2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n821), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n238), .A2(new_n810), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n808), .B1(new_n222), .B2(new_n568), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n991), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(G311), .ZN(new_n995));
  INV_X1    g0795(.A(G303), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n846), .A2(new_n995), .B1(new_n996), .B2(new_n776), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT106), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n787), .A2(new_n250), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n784), .A2(new_n248), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(G294), .C2(new_n766), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n359), .B1(new_n778), .B2(new_n588), .ZN(new_n1002));
  AOI21_X1  g0802(.A(KEYINPUT46), .B1(new_n799), .B2(G116), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n1002), .B(new_n1003), .C1(G317), .C2(new_n793), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n799), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT107), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n998), .A2(new_n1001), .A3(new_n1004), .A4(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n784), .A2(new_n207), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(G150), .B2(new_n792), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n1009), .A2(KEYINPUT108), .B1(new_n789), .B2(G143), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(KEYINPUT108), .B2(new_n1009), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT109), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n258), .B1(new_n300), .B2(new_n778), .C1(new_n767), .C2(new_n772), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n799), .A2(G58), .B1(new_n793), .B2(G137), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n1014), .A2(KEYINPUT110), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n787), .A2(new_n209), .ZN(new_n1016));
  NOR3_X1   g0816(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(KEYINPUT110), .B2(new_n1014), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1007), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT47), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n994), .B1(new_n1020), .B2(new_n762), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n823), .B2(new_n952), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n990), .A2(new_n1022), .ZN(G387));
  OR2_X1    g0823(.A1(new_n723), .A2(new_n823), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n733), .A2(new_n814), .B1(G107), .B2(new_n222), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT111), .Z(new_n1026));
  NOR2_X1   g0826(.A1(new_n410), .A2(G50), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT50), .ZN(new_n1028));
  AOI21_X1  g0828(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1028), .A2(new_n733), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n811), .B1(new_n243), .B2(G45), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1026), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n991), .B1(new_n1032), .B2(new_n809), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n792), .A2(G317), .B1(new_n779), .B2(G303), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(KEYINPUT113), .B(G322), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1034), .B1(new_n767), .B2(new_n995), .C1(new_n846), .C2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT48), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n785), .A2(G283), .B1(new_n799), .B2(G294), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT49), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n787), .A2(new_n502), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n258), .B(new_n1045), .C1(G326), .C2(new_n793), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1043), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G159), .A2(new_n789), .B1(new_n766), .B2(new_n305), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n569), .A2(new_n785), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n776), .A2(new_n300), .B1(new_n778), .B2(new_n207), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(KEYINPUT112), .B(G150), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n258), .B1(new_n771), .B2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n999), .B1(G77), .B2(new_n799), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1048), .A2(new_n1049), .A3(new_n1053), .A4(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1047), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1033), .B1(new_n1056), .B2(new_n762), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n984), .A2(new_n989), .B1(new_n1024), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n985), .A2(new_n731), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n984), .A2(new_n760), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(G393));
  NAND2_X1  g0861(.A1(new_n982), .A2(new_n985), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n986), .A2(new_n1062), .A3(new_n731), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n982), .A2(new_n988), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n959), .A2(new_n807), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n808), .B1(new_n250), .B2(new_n222), .C1(new_n254), .C2(new_n811), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n991), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n846), .A2(new_n844), .B1(new_n772), .B2(new_n776), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT51), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n781), .A2(new_n207), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n784), .A2(new_n209), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(G50), .C2(new_n766), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n410), .A2(new_n778), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n359), .B(new_n855), .C1(G143), .C2(new_n793), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1069), .A2(new_n1072), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(G317), .A2(new_n789), .B1(new_n792), .B2(G311), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT114), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT52), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n785), .A2(G116), .B1(new_n779), .B2(G294), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n996), .B2(new_n767), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT115), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n359), .B1(new_n771), .B2(new_n1035), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n788), .B(new_n1082), .C1(G283), .C2(new_n799), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1075), .B1(new_n1078), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1067), .B1(new_n1085), .B2(new_n762), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1064), .B1(new_n1065), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1063), .A2(new_n1087), .ZN(G390));
  NAND2_X1  g0888(.A1(new_n933), .A2(new_n938), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n927), .B2(new_n939), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n939), .B1(new_n919), .B2(new_n920), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n834), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n714), .B1(new_n704), .B2(new_n757), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1092), .B1(new_n1093), .B2(new_n833), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1091), .B1(new_n1094), .B2(new_n926), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1090), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n752), .A2(new_n837), .A3(new_n911), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1090), .A2(new_n1097), .A3(new_n1095), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n752), .A2(new_n478), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n943), .A2(new_n686), .A3(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n883), .A2(G330), .A3(new_n837), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n926), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n1097), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n838), .A2(new_n834), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1104), .A2(new_n1097), .A3(new_n1094), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1102), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT116), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1099), .B(new_n1100), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(KEYINPUT29), .B1(new_n705), .B2(new_n721), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n477), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1113), .A2(new_n340), .A3(new_n398), .A4(new_n423), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n1112), .A2(new_n1114), .A3(new_n758), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n685), .A2(new_n327), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n752), .A2(new_n478), .ZN(new_n1117));
  NOR3_X1   g0917(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n1104), .A2(new_n1097), .A3(new_n1094), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n1104), .A2(new_n1097), .B1(new_n834), .B2(new_n838), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n1090), .A2(new_n1097), .A3(new_n1095), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1097), .B1(new_n1090), .B2(new_n1095), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1121), .B(KEYINPUT116), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1111), .A2(new_n1124), .A3(new_n731), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n863), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n258), .B1(new_n793), .B2(G294), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n1127), .B1(new_n250), .B2(new_n778), .C1(new_n502), .C2(new_n776), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1071), .B(new_n1128), .C1(G68), .C2(new_n801), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n248), .A2(new_n767), .B1(new_n846), .B2(new_n588), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(G87), .B2(new_n799), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n359), .B1(new_n793), .B2(G125), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT54), .B(G143), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1132), .B1(new_n850), .B2(new_n776), .C1(new_n778), .C2(new_n1133), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n767), .A2(new_n845), .B1(new_n787), .B2(new_n300), .ZN(new_n1135));
  INV_X1    g0935(.A(G128), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n846), .A2(new_n1136), .B1(new_n772), .B2(new_n784), .ZN(new_n1137));
  NOR3_X1   g0937(.A1(new_n1134), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n781), .A2(new_n1051), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT53), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1129), .A2(new_n1131), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n991), .B1(new_n305), .B2(new_n1126), .C1(new_n1141), .C2(new_n763), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n1089), .B2(new_n805), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1143), .B1(new_n1144), .B2(new_n989), .ZN(new_n1145));
  AND2_X1   g0945(.A1(new_n1145), .A2(KEYINPUT117), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1145), .A2(KEYINPUT117), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1125), .B1(new_n1146), .B2(new_n1147), .ZN(G378));
  NAND2_X1  g0948(.A1(new_n910), .A2(new_n882), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT120), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n921), .A2(new_n883), .A3(new_n890), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1149), .A2(new_n1150), .A3(G330), .A4(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n322), .A2(new_n897), .ZN(new_n1153));
  XOR2_X1   g0953(.A(new_n340), .B(new_n1153), .Z(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1154), .B(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1152), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1150), .B1(new_n922), .B2(G330), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1149), .A2(G330), .A3(new_n1151), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1161), .A2(KEYINPUT120), .A3(new_n1156), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n942), .B1(new_n1160), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1161), .A2(KEYINPUT120), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1165), .A2(new_n1152), .A3(new_n1157), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n942), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1166), .A2(new_n1167), .A3(new_n1162), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1099), .A2(new_n1100), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n1118), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1164), .A2(new_n1168), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT57), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n731), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1164), .A2(new_n989), .A3(new_n1168), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n991), .B1(G50), .B2(new_n1126), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(G33), .A2(G41), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT118), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n300), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n359), .B2(new_n486), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n258), .B(new_n729), .C1(G283), .C2(new_n793), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n248), .B2(new_n776), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n569), .B2(new_n779), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n787), .A2(new_n354), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT119), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1008), .B1(G77), .B2(new_n799), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(G97), .A2(new_n766), .B1(new_n789), .B2(G116), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1185), .A2(new_n1187), .A3(new_n1188), .A4(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT58), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1182), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1180), .B1(G124), .B2(new_n793), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n789), .A2(G125), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n767), .B2(new_n850), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n792), .A2(G128), .B1(new_n779), .B2(G137), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n781), .B2(new_n1133), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1195), .B(new_n1197), .C1(G150), .C2(new_n785), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT59), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1193), .B1(new_n772), .B2(new_n787), .C1(new_n1198), .C2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1198), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1201), .A2(KEYINPUT59), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n1192), .B1(new_n1191), .B2(new_n1190), .C1(new_n1200), .C2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1178), .B1(new_n1203), .B2(new_n762), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n1156), .B2(new_n806), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1177), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1176), .A2(new_n1206), .ZN(G375));
  NAND3_X1  g1007(.A1(new_n1107), .A2(new_n1102), .A3(new_n1108), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1121), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n971), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT121), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n911), .A2(new_n806), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT122), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n991), .B1(G68), .B2(new_n1126), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n778), .A2(new_n844), .B1(new_n771), .B2(new_n1136), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n359), .B(new_n1216), .C1(G137), .C2(new_n792), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1133), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G132), .A2(new_n789), .B1(new_n766), .B2(new_n1218), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n785), .A2(G50), .B1(new_n799), .B2(G159), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1217), .A2(new_n1187), .A3(new_n1219), .A4(new_n1220), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n789), .A2(G294), .B1(new_n779), .B2(G107), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n502), .B2(new_n767), .ZN(new_n1223));
  XNOR2_X1  g1023(.A(new_n1223), .B(KEYINPUT123), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n359), .B1(new_n776), .B2(new_n588), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G303), .B2(new_n793), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1016), .B1(G97), .B2(new_n799), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1226), .A2(new_n1049), .A3(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1221), .B1(new_n1224), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1215), .B1(new_n1229), .B2(new_n762), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1169), .A2(new_n989), .B1(new_n1214), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1212), .A2(new_n1231), .ZN(G381));
  OR4_X1    g1032(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(new_n1233), .A2(G387), .A3(G381), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT124), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1125), .A2(new_n1235), .A3(new_n1145), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1235), .B1(new_n1125), .B2(new_n1145), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1234), .A2(new_n1206), .A3(new_n1176), .A4(new_n1239), .ZN(G407));
  NAND2_X1  g1040(.A1(new_n713), .A2(G213), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(G375), .A2(new_n1238), .A3(new_n1241), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(new_n1242), .B(KEYINPUT125), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(G213), .A3(G407), .ZN(G409));
  NAND4_X1  g1044(.A1(new_n1164), .A2(new_n1171), .A3(new_n1210), .A4(new_n1168), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1245), .A2(new_n1177), .A3(new_n1205), .ZN(new_n1246));
  OAI21_X1  g1046(.A(KEYINPUT126), .B1(new_n1238), .B2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G378), .B(new_n1206), .C1(new_n1174), .C2(new_n1175), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1245), .A2(new_n1177), .A3(new_n1205), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT126), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1249), .B(new_n1250), .C1(new_n1236), .C2(new_n1237), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1247), .A2(new_n1248), .A3(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT60), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1209), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1208), .A2(new_n1253), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n731), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1231), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1257));
  OR2_X1    g1057(.A1(new_n1257), .A2(new_n867), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n867), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1252), .A2(new_n1241), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(KEYINPUT62), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1252), .A2(new_n1241), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n713), .A2(G213), .A3(G2897), .ZN(new_n1265));
  XNOR2_X1  g1065(.A(new_n1260), .B(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT61), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT62), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1252), .A2(new_n1269), .A3(new_n1241), .A4(new_n1261), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1263), .A2(new_n1267), .A3(new_n1268), .A4(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(G390), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(G387), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n990), .A2(new_n1022), .A3(G390), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(G393), .B(new_n829), .ZN(new_n1276));
  AOI21_X1  g1076(.A(G390), .B1(new_n990), .B2(new_n1022), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1276), .B1(new_n1277), .B2(KEYINPUT127), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1273), .A2(new_n1276), .A3(KEYINPUT127), .A4(new_n1274), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1271), .A2(new_n1281), .ZN(new_n1282));
  AND2_X1   g1082(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1283));
  AOI21_X1  g1083(.A(KEYINPUT61), .B1(new_n1264), .B2(new_n1266), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT63), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1262), .A2(new_n1285), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1252), .A2(KEYINPUT63), .A3(new_n1241), .A4(new_n1261), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1283), .A2(new_n1284), .A3(new_n1286), .A4(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1282), .A2(new_n1288), .ZN(G405));
  NAND2_X1  g1089(.A1(G375), .A2(new_n1239), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(new_n1260), .A3(new_n1248), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1260), .B1(new_n1290), .B2(new_n1248), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1283), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1281), .B1(new_n1292), .B2(new_n1293), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(G402));
endmodule


