

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U555 ( .A1(G8), .A2(n772), .ZN(n821) );
  NOR2_X1 U556 ( .A1(n642), .A2(n547), .ZN(n668) );
  NOR2_X2 U557 ( .A1(n532), .A2(n531), .ZN(G160) );
  NOR2_X1 U558 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U559 ( .A1(n522), .A2(G2104), .ZN(n563) );
  NAND2_X1 U560 ( .A1(n794), .A2(n786), .ZN(n788) );
  INV_X1 U561 ( .A(KEYINPUT105), .ZN(n787) );
  INV_X1 U562 ( .A(n986), .ZN(n789) );
  XNOR2_X1 U563 ( .A(n592), .B(KEYINPUT73), .ZN(n595) );
  OR2_X1 U564 ( .A1(n821), .A2(n802), .ZN(n520) );
  INV_X1 U565 ( .A(KEYINPUT102), .ZN(n731) );
  NOR2_X1 U566 ( .A1(n724), .A2(n723), .ZN(n736) );
  NOR2_X1 U567 ( .A1(n758), .A2(n757), .ZN(n759) );
  INV_X1 U568 ( .A(KEYINPUT29), .ZN(n749) );
  AND2_X1 U569 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U570 ( .A(n788), .B(n787), .ZN(n791) );
  AND2_X1 U571 ( .A1(n791), .A2(n790), .ZN(n793) );
  OR2_X1 U572 ( .A1(n827), .A2(n826), .ZN(n828) );
  INV_X1 U573 ( .A(G2105), .ZN(n522) );
  AND2_X1 U574 ( .A1(n522), .A2(G2104), .ZN(n619) );
  BUF_X1 U575 ( .A(n619), .Z(n912) );
  NOR2_X1 U576 ( .A1(G651), .A2(n642), .ZN(n665) );
  NAND2_X1 U577 ( .A1(n563), .A2(G125), .ZN(n521) );
  XNOR2_X1 U578 ( .A(KEYINPUT65), .B(n521), .ZN(n525) );
  NAND2_X1 U579 ( .A1(n619), .A2(G101), .ZN(n523) );
  XNOR2_X1 U580 ( .A(KEYINPUT23), .B(n523), .ZN(n524) );
  NOR2_X1 U581 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U582 ( .A(n526), .B(KEYINPUT66), .Z(n532) );
  XNOR2_X1 U583 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n528) );
  NOR2_X1 U584 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  XNOR2_X1 U585 ( .A(n528), .B(n527), .ZN(n622) );
  NAND2_X1 U586 ( .A1(G137), .A2(n622), .ZN(n530) );
  AND2_X1 U587 ( .A1(G2104), .A2(G2105), .ZN(n909) );
  NAND2_X1 U588 ( .A1(G113), .A2(n909), .ZN(n529) );
  NAND2_X1 U589 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U590 ( .A(G2427), .B(KEYINPUT109), .ZN(n542) );
  XOR2_X1 U591 ( .A(G2443), .B(G2438), .Z(n534) );
  XNOR2_X1 U592 ( .A(KEYINPUT108), .B(G2454), .ZN(n533) );
  XNOR2_X1 U593 ( .A(n534), .B(n533), .ZN(n538) );
  XOR2_X1 U594 ( .A(G2430), .B(G2435), .Z(n536) );
  XNOR2_X1 U595 ( .A(G1341), .B(G1348), .ZN(n535) );
  XNOR2_X1 U596 ( .A(n536), .B(n535), .ZN(n537) );
  XOR2_X1 U597 ( .A(n538), .B(n537), .Z(n540) );
  XNOR2_X1 U598 ( .A(G2451), .B(G2446), .ZN(n539) );
  XNOR2_X1 U599 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U600 ( .A(n542), .B(n541), .ZN(n543) );
  AND2_X1 U601 ( .A1(n543), .A2(G14), .ZN(G401) );
  INV_X1 U602 ( .A(G651), .ZN(n547) );
  NOR2_X1 U603 ( .A1(G543), .A2(n547), .ZN(n544) );
  XOR2_X1 U604 ( .A(KEYINPUT1), .B(n544), .Z(n596) );
  BUF_X1 U605 ( .A(n596), .Z(n664) );
  NAND2_X1 U606 ( .A1(G64), .A2(n664), .ZN(n546) );
  XOR2_X1 U607 ( .A(KEYINPUT0), .B(G543), .Z(n642) );
  NAND2_X1 U608 ( .A1(G52), .A2(n665), .ZN(n545) );
  NAND2_X1 U609 ( .A1(n546), .A2(n545), .ZN(n553) );
  NAND2_X1 U610 ( .A1(G77), .A2(n668), .ZN(n549) );
  NOR2_X1 U611 ( .A1(G651), .A2(G543), .ZN(n672) );
  NAND2_X1 U612 ( .A1(G90), .A2(n672), .ZN(n548) );
  NAND2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U614 ( .A(KEYINPUT9), .B(n550), .ZN(n551) );
  XNOR2_X1 U615 ( .A(KEYINPUT69), .B(n551), .ZN(n552) );
  NOR2_X1 U616 ( .A1(n553), .A2(n552), .ZN(G171) );
  AND2_X1 U617 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U618 ( .A1(G65), .A2(n664), .ZN(n555) );
  NAND2_X1 U619 ( .A1(G53), .A2(n665), .ZN(n554) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n559) );
  NAND2_X1 U621 ( .A1(G78), .A2(n668), .ZN(n557) );
  NAND2_X1 U622 ( .A1(G91), .A2(n672), .ZN(n556) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  NOR2_X1 U624 ( .A1(n559), .A2(n558), .ZN(n737) );
  INV_X1 U625 ( .A(n737), .ZN(G299) );
  INV_X1 U626 ( .A(G132), .ZN(G219) );
  INV_X1 U627 ( .A(G82), .ZN(G220) );
  INV_X1 U628 ( .A(G57), .ZN(G237) );
  INV_X1 U629 ( .A(G120), .ZN(G236) );
  INV_X1 U630 ( .A(G108), .ZN(G238) );
  NAND2_X1 U631 ( .A1(n619), .A2(G102), .ZN(n560) );
  XNOR2_X1 U632 ( .A(n560), .B(KEYINPUT90), .ZN(n562) );
  NAND2_X1 U633 ( .A1(G138), .A2(n622), .ZN(n561) );
  NAND2_X1 U634 ( .A1(n562), .A2(n561), .ZN(n568) );
  INV_X1 U635 ( .A(n563), .ZN(n564) );
  INV_X1 U636 ( .A(n564), .ZN(n908) );
  NAND2_X1 U637 ( .A1(G126), .A2(n908), .ZN(n566) );
  NAND2_X1 U638 ( .A1(G114), .A2(n909), .ZN(n565) );
  NAND2_X1 U639 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U640 ( .A1(n568), .A2(n567), .ZN(G164) );
  NAND2_X1 U641 ( .A1(n672), .A2(G89), .ZN(n569) );
  XNOR2_X1 U642 ( .A(n569), .B(KEYINPUT4), .ZN(n571) );
  NAND2_X1 U643 ( .A1(G76), .A2(n668), .ZN(n570) );
  NAND2_X1 U644 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U645 ( .A(KEYINPUT5), .B(n572), .ZN(n578) );
  NAND2_X1 U646 ( .A1(G63), .A2(n664), .ZN(n574) );
  NAND2_X1 U647 ( .A1(G51), .A2(n665), .ZN(n573) );
  NAND2_X1 U648 ( .A1(n574), .A2(n573), .ZN(n576) );
  XOR2_X1 U649 ( .A(KEYINPUT6), .B(KEYINPUT78), .Z(n575) );
  XNOR2_X1 U650 ( .A(n576), .B(n575), .ZN(n577) );
  NAND2_X1 U651 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U652 ( .A(KEYINPUT7), .B(n579), .ZN(G168) );
  XOR2_X1 U653 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U654 ( .A1(G7), .A2(G661), .ZN(n580) );
  XNOR2_X1 U655 ( .A(n580), .B(KEYINPUT10), .ZN(n581) );
  XNOR2_X1 U656 ( .A(KEYINPUT70), .B(n581), .ZN(G223) );
  INV_X1 U657 ( .A(G223), .ZN(n849) );
  NAND2_X1 U658 ( .A1(n849), .A2(G567), .ZN(n582) );
  XOR2_X1 U659 ( .A(KEYINPUT11), .B(n582), .Z(G234) );
  NAND2_X1 U660 ( .A1(n672), .A2(G81), .ZN(n583) );
  XNOR2_X1 U661 ( .A(n583), .B(KEYINPUT12), .ZN(n585) );
  NAND2_X1 U662 ( .A1(G68), .A2(n668), .ZN(n584) );
  NAND2_X1 U663 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U664 ( .A(n586), .B(KEYINPUT13), .ZN(n591) );
  NAND2_X1 U665 ( .A1(G56), .A2(n596), .ZN(n588) );
  XOR2_X1 U666 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n587) );
  XNOR2_X1 U667 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U668 ( .A(KEYINPUT71), .B(n589), .ZN(n590) );
  NAND2_X1 U669 ( .A1(n591), .A2(n590), .ZN(n592) );
  NAND2_X1 U670 ( .A1(n665), .A2(G43), .ZN(n593) );
  XNOR2_X1 U671 ( .A(KEYINPUT74), .B(n593), .ZN(n594) );
  NAND2_X1 U672 ( .A1(n595), .A2(n594), .ZN(n998) );
  INV_X1 U673 ( .A(G860), .ZN(n638) );
  OR2_X1 U674 ( .A1(n998), .A2(n638), .ZN(G153) );
  XNOR2_X1 U675 ( .A(G171), .B(KEYINPUT75), .ZN(G301) );
  NAND2_X1 U676 ( .A1(n665), .A2(G54), .ZN(n603) );
  NAND2_X1 U677 ( .A1(G79), .A2(n668), .ZN(n598) );
  NAND2_X1 U678 ( .A1(G66), .A2(n596), .ZN(n597) );
  NAND2_X1 U679 ( .A1(n598), .A2(n597), .ZN(n601) );
  NAND2_X1 U680 ( .A1(n672), .A2(G92), .ZN(n599) );
  XOR2_X1 U681 ( .A(KEYINPUT76), .B(n599), .Z(n600) );
  NOR2_X1 U682 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U683 ( .A1(n603), .A2(n602), .ZN(n604) );
  XOR2_X1 U684 ( .A(KEYINPUT15), .B(n604), .Z(n984) );
  INV_X1 U685 ( .A(n984), .ZN(n636) );
  NOR2_X1 U686 ( .A1(n636), .A2(G868), .ZN(n605) );
  XNOR2_X1 U687 ( .A(n605), .B(KEYINPUT77), .ZN(n607) );
  NAND2_X1 U688 ( .A1(G868), .A2(G301), .ZN(n606) );
  NAND2_X1 U689 ( .A1(n607), .A2(n606), .ZN(G284) );
  XNOR2_X1 U690 ( .A(KEYINPUT79), .B(G868), .ZN(n608) );
  NOR2_X1 U691 ( .A1(G286), .A2(n608), .ZN(n609) );
  XNOR2_X1 U692 ( .A(n609), .B(KEYINPUT80), .ZN(n611) );
  NOR2_X1 U693 ( .A1(G299), .A2(G868), .ZN(n610) );
  NOR2_X1 U694 ( .A1(n611), .A2(n610), .ZN(G297) );
  NAND2_X1 U695 ( .A1(n638), .A2(G559), .ZN(n612) );
  NAND2_X1 U696 ( .A1(n612), .A2(n636), .ZN(n613) );
  XNOR2_X1 U697 ( .A(n613), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U698 ( .A1(G868), .A2(n998), .ZN(n616) );
  NAND2_X1 U699 ( .A1(G868), .A2(n636), .ZN(n614) );
  NOR2_X1 U700 ( .A1(G559), .A2(n614), .ZN(n615) );
  NOR2_X1 U701 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U702 ( .A(KEYINPUT81), .B(n617), .Z(G282) );
  NAND2_X1 U703 ( .A1(G123), .A2(n908), .ZN(n618) );
  XNOR2_X1 U704 ( .A(n618), .B(KEYINPUT18), .ZN(n621) );
  NAND2_X1 U705 ( .A1(n912), .A2(G99), .ZN(n620) );
  NAND2_X1 U706 ( .A1(n621), .A2(n620), .ZN(n626) );
  BUF_X1 U707 ( .A(n622), .Z(n913) );
  NAND2_X1 U708 ( .A1(G135), .A2(n913), .ZN(n624) );
  NAND2_X1 U709 ( .A1(G111), .A2(n909), .ZN(n623) );
  NAND2_X1 U710 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U711 ( .A1(n626), .A2(n625), .ZN(n942) );
  XNOR2_X1 U712 ( .A(G2096), .B(n942), .ZN(n628) );
  INV_X1 U713 ( .A(G2100), .ZN(n627) );
  NAND2_X1 U714 ( .A1(n628), .A2(n627), .ZN(G156) );
  NAND2_X1 U715 ( .A1(G80), .A2(n668), .ZN(n630) );
  NAND2_X1 U716 ( .A1(G93), .A2(n672), .ZN(n629) );
  NAND2_X1 U717 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U718 ( .A(KEYINPUT82), .B(n631), .ZN(n635) );
  NAND2_X1 U719 ( .A1(G67), .A2(n664), .ZN(n633) );
  NAND2_X1 U720 ( .A1(G55), .A2(n665), .ZN(n632) );
  NAND2_X1 U721 ( .A1(n633), .A2(n632), .ZN(n634) );
  OR2_X1 U722 ( .A1(n635), .A2(n634), .ZN(n684) );
  NAND2_X1 U723 ( .A1(G559), .A2(n636), .ZN(n637) );
  XOR2_X1 U724 ( .A(n998), .B(n637), .Z(n681) );
  NAND2_X1 U725 ( .A1(n638), .A2(n681), .ZN(n639) );
  XNOR2_X1 U726 ( .A(n639), .B(KEYINPUT83), .ZN(n640) );
  XOR2_X1 U727 ( .A(n684), .B(n640), .Z(G145) );
  NAND2_X1 U728 ( .A1(G49), .A2(n665), .ZN(n641) );
  XNOR2_X1 U729 ( .A(n641), .B(KEYINPUT84), .ZN(n647) );
  NAND2_X1 U730 ( .A1(G87), .A2(n642), .ZN(n644) );
  NAND2_X1 U731 ( .A1(G74), .A2(G651), .ZN(n643) );
  NAND2_X1 U732 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U733 ( .A1(n664), .A2(n645), .ZN(n646) );
  NAND2_X1 U734 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U735 ( .A(KEYINPUT85), .B(n648), .Z(G288) );
  NAND2_X1 U736 ( .A1(G62), .A2(n664), .ZN(n650) );
  NAND2_X1 U737 ( .A1(G88), .A2(n672), .ZN(n649) );
  NAND2_X1 U738 ( .A1(n650), .A2(n649), .ZN(n653) );
  NAND2_X1 U739 ( .A1(G50), .A2(n665), .ZN(n651) );
  XNOR2_X1 U740 ( .A(KEYINPUT87), .B(n651), .ZN(n652) );
  NOR2_X1 U741 ( .A1(n653), .A2(n652), .ZN(n655) );
  NAND2_X1 U742 ( .A1(n668), .A2(G75), .ZN(n654) );
  NAND2_X1 U743 ( .A1(n655), .A2(n654), .ZN(G303) );
  INV_X1 U744 ( .A(G303), .ZN(G166) );
  NAND2_X1 U745 ( .A1(G61), .A2(n664), .ZN(n657) );
  NAND2_X1 U746 ( .A1(G86), .A2(n672), .ZN(n656) );
  NAND2_X1 U747 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U748 ( .A(KEYINPUT86), .B(n658), .ZN(n661) );
  NAND2_X1 U749 ( .A1(n668), .A2(G73), .ZN(n659) );
  XOR2_X1 U750 ( .A(KEYINPUT2), .B(n659), .Z(n660) );
  NOR2_X1 U751 ( .A1(n661), .A2(n660), .ZN(n663) );
  NAND2_X1 U752 ( .A1(n665), .A2(G48), .ZN(n662) );
  NAND2_X1 U753 ( .A1(n663), .A2(n662), .ZN(G305) );
  NAND2_X1 U754 ( .A1(G60), .A2(n664), .ZN(n667) );
  NAND2_X1 U755 ( .A1(G47), .A2(n665), .ZN(n666) );
  NAND2_X1 U756 ( .A1(n667), .A2(n666), .ZN(n671) );
  NAND2_X1 U757 ( .A1(G72), .A2(n668), .ZN(n669) );
  XOR2_X1 U758 ( .A(KEYINPUT68), .B(n669), .Z(n670) );
  NOR2_X1 U759 ( .A1(n671), .A2(n670), .ZN(n674) );
  NAND2_X1 U760 ( .A1(n672), .A2(G85), .ZN(n673) );
  NAND2_X1 U761 ( .A1(n674), .A2(n673), .ZN(G290) );
  INV_X1 U762 ( .A(G868), .ZN(n683) );
  XOR2_X1 U763 ( .A(KEYINPUT19), .B(KEYINPUT88), .Z(n675) );
  XNOR2_X1 U764 ( .A(G305), .B(n675), .ZN(n676) );
  XNOR2_X1 U765 ( .A(G166), .B(n676), .ZN(n678) );
  XNOR2_X1 U766 ( .A(G290), .B(n737), .ZN(n677) );
  XNOR2_X1 U767 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U768 ( .A(n684), .B(n679), .ZN(n680) );
  XNOR2_X1 U769 ( .A(G288), .B(n680), .ZN(n858) );
  XOR2_X1 U770 ( .A(n858), .B(n681), .Z(n682) );
  NOR2_X1 U771 ( .A1(n683), .A2(n682), .ZN(n686) );
  NOR2_X1 U772 ( .A1(G868), .A2(n684), .ZN(n685) );
  NOR2_X1 U773 ( .A1(n686), .A2(n685), .ZN(G295) );
  NAND2_X1 U774 ( .A1(G2078), .A2(G2084), .ZN(n687) );
  XOR2_X1 U775 ( .A(KEYINPUT20), .B(n687), .Z(n688) );
  NAND2_X1 U776 ( .A1(G2090), .A2(n688), .ZN(n689) );
  XNOR2_X1 U777 ( .A(KEYINPUT21), .B(n689), .ZN(n690) );
  NAND2_X1 U778 ( .A1(n690), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U779 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U780 ( .A1(G238), .A2(G236), .ZN(n691) );
  NAND2_X1 U781 ( .A1(G69), .A2(n691), .ZN(n692) );
  NOR2_X1 U782 ( .A1(n692), .A2(G237), .ZN(n693) );
  XNOR2_X1 U783 ( .A(n693), .B(KEYINPUT89), .ZN(n854) );
  NAND2_X1 U784 ( .A1(n854), .A2(G567), .ZN(n698) );
  NOR2_X1 U785 ( .A1(G220), .A2(G219), .ZN(n694) );
  XOR2_X1 U786 ( .A(KEYINPUT22), .B(n694), .Z(n695) );
  NOR2_X1 U787 ( .A1(G218), .A2(n695), .ZN(n696) );
  NAND2_X1 U788 ( .A1(G96), .A2(n696), .ZN(n855) );
  NAND2_X1 U789 ( .A1(n855), .A2(G2106), .ZN(n697) );
  NAND2_X1 U790 ( .A1(n698), .A2(n697), .ZN(n931) );
  NAND2_X1 U791 ( .A1(G483), .A2(G661), .ZN(n699) );
  NOR2_X1 U792 ( .A1(n931), .A2(n699), .ZN(n851) );
  NAND2_X1 U793 ( .A1(n851), .A2(G36), .ZN(G176) );
  NAND2_X1 U794 ( .A1(G107), .A2(n909), .ZN(n700) );
  XNOR2_X1 U795 ( .A(n700), .B(KEYINPUT94), .ZN(n707) );
  NAND2_X1 U796 ( .A1(G119), .A2(n908), .ZN(n702) );
  NAND2_X1 U797 ( .A1(G131), .A2(n913), .ZN(n701) );
  NAND2_X1 U798 ( .A1(n702), .A2(n701), .ZN(n705) );
  NAND2_X1 U799 ( .A1(G95), .A2(n912), .ZN(n703) );
  XNOR2_X1 U800 ( .A(KEYINPUT95), .B(n703), .ZN(n704) );
  NOR2_X1 U801 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U802 ( .A1(n707), .A2(n706), .ZN(n898) );
  XNOR2_X1 U803 ( .A(KEYINPUT96), .B(G1991), .ZN(n961) );
  NAND2_X1 U804 ( .A1(n898), .A2(n961), .ZN(n717) );
  NAND2_X1 U805 ( .A1(G105), .A2(n912), .ZN(n708) );
  XNOR2_X1 U806 ( .A(n708), .B(KEYINPUT38), .ZN(n715) );
  NAND2_X1 U807 ( .A1(G129), .A2(n908), .ZN(n710) );
  NAND2_X1 U808 ( .A1(G141), .A2(n913), .ZN(n709) );
  NAND2_X1 U809 ( .A1(n710), .A2(n709), .ZN(n713) );
  NAND2_X1 U810 ( .A1(G117), .A2(n909), .ZN(n711) );
  XNOR2_X1 U811 ( .A(KEYINPUT97), .B(n711), .ZN(n712) );
  NOR2_X1 U812 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U813 ( .A1(n715), .A2(n714), .ZN(n919) );
  NAND2_X1 U814 ( .A1(G1996), .A2(n919), .ZN(n716) );
  NAND2_X1 U815 ( .A1(n717), .A2(n716), .ZN(n949) );
  NOR2_X1 U816 ( .A1(G164), .A2(G1384), .ZN(n720) );
  NAND2_X1 U817 ( .A1(G160), .A2(G40), .ZN(n718) );
  NOR2_X1 U818 ( .A1(n720), .A2(n718), .ZN(n844) );
  NAND2_X1 U819 ( .A1(n949), .A2(n844), .ZN(n719) );
  XOR2_X1 U820 ( .A(KEYINPUT98), .B(n719), .Z(n835) );
  AND2_X1 U821 ( .A1(n720), .A2(G40), .ZN(n721) );
  NAND2_X2 U822 ( .A1(G160), .A2(n721), .ZN(n772) );
  NOR2_X1 U823 ( .A1(G2084), .A2(n772), .ZN(n758) );
  NAND2_X1 U824 ( .A1(G8), .A2(n758), .ZN(n769) );
  INV_X1 U825 ( .A(n772), .ZN(n733) );
  NAND2_X1 U826 ( .A1(n733), .A2(G2072), .ZN(n722) );
  XNOR2_X1 U827 ( .A(n722), .B(KEYINPUT27), .ZN(n724) );
  AND2_X1 U828 ( .A1(G1956), .A2(n772), .ZN(n723) );
  NOR2_X1 U829 ( .A1(n737), .A2(n736), .ZN(n725) );
  XOR2_X1 U830 ( .A(n725), .B(KEYINPUT28), .Z(n748) );
  NAND2_X1 U831 ( .A1(G1341), .A2(n772), .ZN(n726) );
  XNOR2_X1 U832 ( .A(KEYINPUT101), .B(n726), .ZN(n727) );
  NOR2_X1 U833 ( .A1(n998), .A2(n727), .ZN(n730) );
  NAND2_X1 U834 ( .A1(G1996), .A2(n733), .ZN(n728) );
  XNOR2_X1 U835 ( .A(n728), .B(KEYINPUT26), .ZN(n729) );
  NAND2_X1 U836 ( .A1(n730), .A2(n729), .ZN(n742) );
  NOR2_X1 U837 ( .A1(n742), .A2(n984), .ZN(n732) );
  XNOR2_X1 U838 ( .A(n732), .B(n731), .ZN(n740) );
  NOR2_X1 U839 ( .A1(n733), .A2(G1348), .ZN(n735) );
  NOR2_X1 U840 ( .A1(G2067), .A2(n772), .ZN(n734) );
  NOR2_X1 U841 ( .A1(n735), .A2(n734), .ZN(n738) );
  NAND2_X1 U842 ( .A1(n737), .A2(n736), .ZN(n741) );
  AND2_X1 U843 ( .A1(n738), .A2(n741), .ZN(n739) );
  NAND2_X1 U844 ( .A1(n740), .A2(n739), .ZN(n746) );
  INV_X1 U845 ( .A(n741), .ZN(n744) );
  NAND2_X1 U846 ( .A1(n742), .A2(n984), .ZN(n743) );
  OR2_X1 U847 ( .A1(n744), .A2(n743), .ZN(n745) );
  AND2_X1 U848 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U849 ( .A1(n748), .A2(n747), .ZN(n750) );
  XNOR2_X1 U850 ( .A(n750), .B(n749), .ZN(n755) );
  NOR2_X1 U851 ( .A1(n733), .A2(G1961), .ZN(n751) );
  XOR2_X1 U852 ( .A(KEYINPUT100), .B(n751), .Z(n753) );
  XNOR2_X1 U853 ( .A(G2078), .B(KEYINPUT25), .ZN(n966) );
  NAND2_X1 U854 ( .A1(n733), .A2(n966), .ZN(n752) );
  NAND2_X1 U855 ( .A1(n753), .A2(n752), .ZN(n761) );
  NAND2_X1 U856 ( .A1(n761), .A2(G171), .ZN(n754) );
  NAND2_X1 U857 ( .A1(n755), .A2(n754), .ZN(n766) );
  NOR2_X1 U858 ( .A1(n821), .A2(G1966), .ZN(n756) );
  XNOR2_X1 U859 ( .A(n756), .B(KEYINPUT99), .ZN(n767) );
  NAND2_X1 U860 ( .A1(G8), .A2(n767), .ZN(n757) );
  XOR2_X1 U861 ( .A(KEYINPUT30), .B(n759), .Z(n760) );
  NOR2_X1 U862 ( .A1(G168), .A2(n760), .ZN(n763) );
  NOR2_X1 U863 ( .A1(G171), .A2(n761), .ZN(n762) );
  XOR2_X1 U864 ( .A(KEYINPUT31), .B(n764), .Z(n765) );
  NAND2_X1 U865 ( .A1(n766), .A2(n765), .ZN(n771) );
  AND2_X1 U866 ( .A1(n771), .A2(n767), .ZN(n768) );
  NAND2_X1 U867 ( .A1(n769), .A2(n768), .ZN(n784) );
  AND2_X1 U868 ( .A1(G286), .A2(G8), .ZN(n770) );
  NAND2_X1 U869 ( .A1(n771), .A2(n770), .ZN(n781) );
  INV_X1 U870 ( .A(G8), .ZN(n779) );
  NOR2_X1 U871 ( .A1(G2090), .A2(n772), .ZN(n773) );
  XOR2_X1 U872 ( .A(KEYINPUT103), .B(n773), .Z(n775) );
  NOR2_X1 U873 ( .A1(G1971), .A2(n821), .ZN(n774) );
  NOR2_X1 U874 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U875 ( .A(n776), .B(KEYINPUT104), .ZN(n777) );
  NAND2_X1 U876 ( .A1(n777), .A2(G303), .ZN(n778) );
  OR2_X1 U877 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U878 ( .A(n782), .B(KEYINPUT32), .ZN(n783) );
  NAND2_X1 U879 ( .A1(n784), .A2(n783), .ZN(n794) );
  NOR2_X1 U880 ( .A1(G1976), .A2(G288), .ZN(n990) );
  NOR2_X1 U881 ( .A1(G1971), .A2(G303), .ZN(n785) );
  NOR2_X1 U882 ( .A1(n990), .A2(n785), .ZN(n786) );
  NAND2_X1 U883 ( .A1(G1976), .A2(G288), .ZN(n986) );
  NOR2_X1 U884 ( .A1(n789), .A2(n821), .ZN(n790) );
  INV_X1 U885 ( .A(KEYINPUT64), .ZN(n792) );
  XNOR2_X1 U886 ( .A(n793), .B(n792), .ZN(n819) );
  INV_X1 U887 ( .A(KEYINPUT33), .ZN(n817) );
  INV_X1 U888 ( .A(n794), .ZN(n797) );
  NAND2_X1 U889 ( .A1(G166), .A2(G8), .ZN(n795) );
  NOR2_X1 U890 ( .A1(G2090), .A2(n795), .ZN(n796) );
  NOR2_X1 U891 ( .A1(n797), .A2(n796), .ZN(n799) );
  INV_X1 U892 ( .A(n821), .ZN(n798) );
  NOR2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n800) );
  INV_X1 U894 ( .A(n800), .ZN(n803) );
  NOR2_X1 U895 ( .A1(G1981), .A2(G305), .ZN(n801) );
  XOR2_X1 U896 ( .A(n801), .B(KEYINPUT24), .Z(n802) );
  NAND2_X1 U897 ( .A1(n803), .A2(n520), .ZN(n816) );
  XNOR2_X1 U898 ( .A(G2067), .B(KEYINPUT37), .ZN(n842) );
  XNOR2_X1 U899 ( .A(KEYINPUT93), .B(KEYINPUT36), .ZN(n815) );
  NAND2_X1 U900 ( .A1(n909), .A2(G116), .ZN(n804) );
  XNOR2_X1 U901 ( .A(n804), .B(KEYINPUT92), .ZN(n806) );
  NAND2_X1 U902 ( .A1(G128), .A2(n908), .ZN(n805) );
  NAND2_X1 U903 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U904 ( .A(n807), .B(KEYINPUT35), .ZN(n813) );
  XNOR2_X1 U905 ( .A(KEYINPUT91), .B(KEYINPUT34), .ZN(n811) );
  NAND2_X1 U906 ( .A1(G104), .A2(n912), .ZN(n809) );
  NAND2_X1 U907 ( .A1(G140), .A2(n913), .ZN(n808) );
  NAND2_X1 U908 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U909 ( .A(n811), .B(n810), .ZN(n812) );
  NAND2_X1 U910 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U911 ( .A(n815), .B(n814), .ZN(n894) );
  NOR2_X1 U912 ( .A1(n842), .A2(n894), .ZN(n945) );
  NAND2_X1 U913 ( .A1(n844), .A2(n945), .ZN(n840) );
  NAND2_X1 U914 ( .A1(n816), .A2(n840), .ZN(n820) );
  AND2_X1 U915 ( .A1(n817), .A2(n820), .ZN(n818) );
  NAND2_X1 U916 ( .A1(n819), .A2(n818), .ZN(n829) );
  INV_X1 U917 ( .A(n820), .ZN(n827) );
  NAND2_X1 U918 ( .A1(n990), .A2(KEYINPUT33), .ZN(n822) );
  NOR2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n824) );
  XOR2_X1 U920 ( .A(G1981), .B(G305), .Z(n980) );
  INV_X1 U921 ( .A(n980), .ZN(n823) );
  NOR2_X1 U922 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U923 ( .A1(n825), .A2(n840), .ZN(n826) );
  NAND2_X1 U924 ( .A1(n829), .A2(n828), .ZN(n830) );
  NOR2_X1 U925 ( .A1(n835), .A2(n830), .ZN(n831) );
  XNOR2_X1 U926 ( .A(n831), .B(KEYINPUT106), .ZN(n833) );
  XNOR2_X1 U927 ( .A(G1986), .B(G290), .ZN(n988) );
  NAND2_X1 U928 ( .A1(n988), .A2(n844), .ZN(n832) );
  NAND2_X1 U929 ( .A1(n833), .A2(n832), .ZN(n847) );
  XOR2_X1 U930 ( .A(KEYINPUT39), .B(KEYINPUT107), .Z(n839) );
  NOR2_X1 U931 ( .A1(G1996), .A2(n919), .ZN(n937) );
  NOR2_X1 U932 ( .A1(n961), .A2(n898), .ZN(n943) );
  NOR2_X1 U933 ( .A1(G1986), .A2(G290), .ZN(n834) );
  NOR2_X1 U934 ( .A1(n943), .A2(n834), .ZN(n836) );
  NOR2_X1 U935 ( .A1(n836), .A2(n835), .ZN(n837) );
  NOR2_X1 U936 ( .A1(n937), .A2(n837), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n841) );
  NAND2_X1 U938 ( .A1(n841), .A2(n840), .ZN(n843) );
  NAND2_X1 U939 ( .A1(n842), .A2(n894), .ZN(n952) );
  NAND2_X1 U940 ( .A1(n843), .A2(n952), .ZN(n845) );
  NAND2_X1 U941 ( .A1(n845), .A2(n844), .ZN(n846) );
  NAND2_X1 U942 ( .A1(n847), .A2(n846), .ZN(n848) );
  XNOR2_X1 U943 ( .A(KEYINPUT40), .B(n848), .ZN(G329) );
  NAND2_X1 U944 ( .A1(G2106), .A2(n849), .ZN(G217) );
  AND2_X1 U945 ( .A1(G15), .A2(G2), .ZN(n850) );
  NAND2_X1 U946 ( .A1(G661), .A2(n850), .ZN(G259) );
  NAND2_X1 U947 ( .A1(G1), .A2(G3), .ZN(n852) );
  NAND2_X1 U948 ( .A1(n852), .A2(n851), .ZN(n853) );
  XNOR2_X1 U949 ( .A(n853), .B(KEYINPUT110), .ZN(G188) );
  XNOR2_X1 U950 ( .A(G69), .B(KEYINPUT111), .ZN(G235) );
  INV_X1 U952 ( .A(G96), .ZN(G221) );
  NOR2_X1 U953 ( .A1(n855), .A2(n854), .ZN(G325) );
  INV_X1 U954 ( .A(G325), .ZN(G261) );
  XOR2_X1 U955 ( .A(G171), .B(KEYINPUT119), .Z(n856) );
  XNOR2_X1 U956 ( .A(n984), .B(n856), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n860) );
  XNOR2_X1 U958 ( .A(n998), .B(G286), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n861) );
  NOR2_X1 U960 ( .A1(G37), .A2(n861), .ZN(G397) );
  XOR2_X1 U961 ( .A(G2474), .B(G1981), .Z(n863) );
  XNOR2_X1 U962 ( .A(G1966), .B(G1956), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U964 ( .A(n864), .B(KEYINPUT113), .Z(n866) );
  XNOR2_X1 U965 ( .A(G1996), .B(G1991), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U967 ( .A(G1976), .B(G1971), .Z(n868) );
  XNOR2_X1 U968 ( .A(G1986), .B(G1961), .ZN(n867) );
  XNOR2_X1 U969 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U970 ( .A(n870), .B(n869), .Z(n872) );
  XNOR2_X1 U971 ( .A(KEYINPUT114), .B(KEYINPUT41), .ZN(n871) );
  XNOR2_X1 U972 ( .A(n872), .B(n871), .ZN(G229) );
  XOR2_X1 U973 ( .A(G2096), .B(KEYINPUT43), .Z(n874) );
  XNOR2_X1 U974 ( .A(G2072), .B(G2678), .ZN(n873) );
  XNOR2_X1 U975 ( .A(n874), .B(n873), .ZN(n875) );
  XOR2_X1 U976 ( .A(n875), .B(KEYINPUT42), .Z(n877) );
  XNOR2_X1 U977 ( .A(G2067), .B(G2090), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n877), .B(n876), .ZN(n881) );
  XOR2_X1 U979 ( .A(KEYINPUT112), .B(G2100), .Z(n879) );
  XNOR2_X1 U980 ( .A(G2078), .B(G2084), .ZN(n878) );
  XNOR2_X1 U981 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U982 ( .A(n881), .B(n880), .ZN(G227) );
  NAND2_X1 U983 ( .A1(G100), .A2(n912), .ZN(n883) );
  NAND2_X1 U984 ( .A1(G112), .A2(n909), .ZN(n882) );
  NAND2_X1 U985 ( .A1(n883), .A2(n882), .ZN(n890) );
  NAND2_X1 U986 ( .A1(G136), .A2(n913), .ZN(n884) );
  XNOR2_X1 U987 ( .A(n884), .B(KEYINPUT116), .ZN(n888) );
  XOR2_X1 U988 ( .A(KEYINPUT44), .B(KEYINPUT115), .Z(n886) );
  NAND2_X1 U989 ( .A1(G124), .A2(n908), .ZN(n885) );
  XNOR2_X1 U990 ( .A(n886), .B(n885), .ZN(n887) );
  NAND2_X1 U991 ( .A1(n888), .A2(n887), .ZN(n889) );
  NOR2_X1 U992 ( .A1(n890), .A2(n889), .ZN(G162) );
  XOR2_X1 U993 ( .A(KEYINPUT48), .B(KEYINPUT118), .Z(n892) );
  XNOR2_X1 U994 ( .A(KEYINPUT46), .B(KEYINPUT117), .ZN(n891) );
  XNOR2_X1 U995 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U996 ( .A(G162), .B(n893), .ZN(n896) );
  XNOR2_X1 U997 ( .A(n894), .B(n942), .ZN(n895) );
  XNOR2_X1 U998 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U999 ( .A(n898), .B(n897), .ZN(n900) );
  XNOR2_X1 U1000 ( .A(G164), .B(G160), .ZN(n899) );
  XNOR2_X1 U1001 ( .A(n900), .B(n899), .ZN(n923) );
  NAND2_X1 U1002 ( .A1(G103), .A2(n912), .ZN(n902) );
  NAND2_X1 U1003 ( .A1(G139), .A2(n913), .ZN(n901) );
  NAND2_X1 U1004 ( .A1(n902), .A2(n901), .ZN(n907) );
  NAND2_X1 U1005 ( .A1(G127), .A2(n908), .ZN(n904) );
  NAND2_X1 U1006 ( .A1(G115), .A2(n909), .ZN(n903) );
  NAND2_X1 U1007 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1008 ( .A(KEYINPUT47), .B(n905), .Z(n906) );
  NOR2_X1 U1009 ( .A1(n907), .A2(n906), .ZN(n932) );
  NAND2_X1 U1010 ( .A1(G130), .A2(n908), .ZN(n911) );
  NAND2_X1 U1011 ( .A1(G118), .A2(n909), .ZN(n910) );
  NAND2_X1 U1012 ( .A1(n911), .A2(n910), .ZN(n918) );
  NAND2_X1 U1013 ( .A1(G106), .A2(n912), .ZN(n915) );
  NAND2_X1 U1014 ( .A1(G142), .A2(n913), .ZN(n914) );
  NAND2_X1 U1015 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1016 ( .A(n916), .B(KEYINPUT45), .Z(n917) );
  NOR2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n920) );
  XNOR2_X1 U1018 ( .A(n920), .B(n919), .ZN(n921) );
  XNOR2_X1 U1019 ( .A(n932), .B(n921), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(n923), .B(n922), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(G37), .A2(n924), .ZN(G395) );
  NOR2_X1 U1022 ( .A1(G401), .A2(n931), .ZN(n928) );
  NOR2_X1 U1023 ( .A1(G229), .A2(G227), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(KEYINPUT49), .B(n925), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(G397), .A2(n926), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1027 ( .A1(n929), .A2(G395), .ZN(n930) );
  XNOR2_X1 U1028 ( .A(n930), .B(KEYINPUT120), .ZN(G308) );
  INV_X1 U1029 ( .A(G308), .ZN(G225) );
  INV_X1 U1030 ( .A(n931), .ZN(G319) );
  XOR2_X1 U1031 ( .A(G2072), .B(n932), .Z(n934) );
  XOR2_X1 U1032 ( .A(G164), .B(G2078), .Z(n933) );
  NOR2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(KEYINPUT50), .B(n935), .ZN(n941) );
  XOR2_X1 U1035 ( .A(G2090), .B(G162), .Z(n936) );
  NOR2_X1 U1036 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1037 ( .A(KEYINPUT51), .B(n938), .Z(n939) );
  XNOR2_X1 U1038 ( .A(KEYINPUT122), .B(n939), .ZN(n940) );
  NAND2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n954) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n947) );
  XOR2_X1 U1041 ( .A(G160), .B(G2084), .Z(n944) );
  NOR2_X1 U1042 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  NOR2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1045 ( .A(KEYINPUT121), .B(n950), .Z(n951) );
  NAND2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  NOR2_X1 U1047 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1048 ( .A(KEYINPUT52), .B(n955), .ZN(n956) );
  INV_X1 U1049 ( .A(KEYINPUT55), .ZN(n976) );
  NAND2_X1 U1050 ( .A1(n956), .A2(n976), .ZN(n957) );
  NAND2_X1 U1051 ( .A1(n957), .A2(G29), .ZN(n1035) );
  XNOR2_X1 U1052 ( .A(G2090), .B(G35), .ZN(n971) );
  XNOR2_X1 U1053 ( .A(G1996), .B(G32), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(G33), .B(G2072), .ZN(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n965) );
  XOR2_X1 U1056 ( .A(G2067), .B(G26), .Z(n960) );
  NAND2_X1 U1057 ( .A1(n960), .A2(G28), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(G25), .B(n961), .ZN(n962) );
  NOR2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n968) );
  XOR2_X1 U1061 ( .A(G27), .B(n966), .Z(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(KEYINPUT53), .B(n969), .ZN(n970) );
  NOR2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n974) );
  XOR2_X1 U1065 ( .A(G2084), .B(G34), .Z(n972) );
  XNOR2_X1 U1066 ( .A(KEYINPUT54), .B(n972), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n976), .B(n975), .ZN(n978) );
  INV_X1 U1069 ( .A(G29), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(G11), .A2(n979), .ZN(n1033) );
  XNOR2_X1 U1072 ( .A(G16), .B(KEYINPUT56), .ZN(n1004) );
  XNOR2_X1 U1073 ( .A(G1966), .B(G168), .ZN(n981) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(n982), .B(KEYINPUT57), .ZN(n1002) );
  XNOR2_X1 U1076 ( .A(G1971), .B(KEYINPUT123), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(n983), .B(G303), .ZN(n996) );
  XOR2_X1 U1078 ( .A(G1348), .B(n984), .Z(n985) );
  NAND2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n994) );
  XNOR2_X1 U1080 ( .A(G1956), .B(G299), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n992) );
  XOR2_X1 U1082 ( .A(G1961), .B(G171), .Z(n989) );
  NOR2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(KEYINPUT124), .B(n997), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(G1341), .B(n998), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1031) );
  INV_X1 U1092 ( .A(G16), .ZN(n1029) );
  XNOR2_X1 U1093 ( .A(KEYINPUT125), .B(G1956), .ZN(n1005) );
  XNOR2_X1 U1094 ( .A(n1005), .B(G20), .ZN(n1011) );
  XNOR2_X1 U1095 ( .A(KEYINPUT59), .B(KEYINPUT127), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(n1006), .B(G4), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(G1348), .B(n1007), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(G1981), .B(G6), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1014) );
  XNOR2_X1 U1101 ( .A(KEYINPUT126), .B(G1341), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(G19), .B(n1012), .ZN(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1104 ( .A(KEYINPUT60), .B(n1015), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(G1966), .B(G21), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(G1961), .B(G5), .ZN(n1016) );
  NOR2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1026) );
  XNOR2_X1 U1109 ( .A(G1971), .B(G22), .ZN(n1021) );
  XNOR2_X1 U1110 ( .A(G23), .B(G1976), .ZN(n1020) );
  NOR2_X1 U1111 ( .A1(n1021), .A2(n1020), .ZN(n1023) );
  XOR2_X1 U1112 ( .A(G1986), .B(G24), .Z(n1022) );
  NAND2_X1 U1113 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1114 ( .A(KEYINPUT58), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1116 ( .A(KEYINPUT61), .B(n1027), .ZN(n1028) );
  NAND2_X1 U1117 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1119 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1120 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XOR2_X1 U1121 ( .A(KEYINPUT62), .B(n1036), .Z(G311) );
  INV_X1 U1122 ( .A(G311), .ZN(G150) );
endmodule

