//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1274, new_n1275, new_n1276, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0003(.A1(G97), .A2(G107), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n205), .A2(G87), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT67), .B(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G58), .A2(G232), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n212), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  NAND3_X1  g0024(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(KEYINPUT65), .B1(G1), .B2(G13), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(new_n210), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n202), .A2(G50), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT66), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n215), .B1(KEYINPUT1), .B2(new_n224), .C1(new_n230), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G50), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G68), .ZN(new_n247));
  INV_X1    g0047(.A(G68), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G50), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n245), .B(new_n252), .ZN(G351));
  XNOR2_X1  g0053(.A(KEYINPUT3), .B(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(G222), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G77), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(G1698), .ZN(new_n258));
  INV_X1    g0058(.A(G223), .ZN(new_n259));
  OAI221_X1 g0059(.A(new_n256), .B1(new_n257), .B2(new_n254), .C1(new_n258), .C2(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n228), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G274), .ZN(new_n264));
  AND2_X1   g0064(.A1(G1), .A2(G13), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT68), .B(G45), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n267), .B(new_n209), .C1(new_n268), .C2(G41), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT69), .B(G1), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n270), .A2(G45), .B1(new_n265), .B2(new_n266), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n209), .A2(KEYINPUT69), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT69), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G1), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(new_n274), .A3(G41), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G226), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n263), .A2(new_n269), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G190), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n280), .B1(G200), .B2(new_n278), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n272), .A2(new_n274), .A3(G13), .A4(G20), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G1), .A2(G13), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT65), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g0085(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n286));
  AND3_X1   g0086(.A1(new_n285), .A2(new_n225), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n270), .A2(G20), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  MUX2_X1   g0089(.A(new_n282), .B(new_n289), .S(G50), .Z(new_n290));
  NAND3_X1  g0090(.A1(new_n285), .A2(new_n225), .A3(new_n286), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n210), .B1(new_n201), .B2(new_n246), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT71), .ZN(new_n293));
  INV_X1    g0093(.A(G33), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n210), .A2(new_n294), .A3(KEYINPUT70), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT70), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n296), .B1(G20), .B2(G33), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G150), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n210), .A2(G33), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT8), .B(G58), .ZN(new_n301));
  OAI22_X1  g0101(.A1(new_n298), .A2(new_n299), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n291), .B1(new_n293), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n290), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(KEYINPUT73), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT73), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n306), .B1(new_n290), .B2(new_n303), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n308), .A2(new_n309), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n281), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT10), .ZN(new_n314));
  INV_X1    g0114(.A(new_n312), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n310), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT10), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(new_n317), .A3(new_n281), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n298), .A2(new_n246), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n248), .A2(KEYINPUT67), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT67), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G68), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n324), .A2(new_n210), .B1(new_n257), .B2(new_n300), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n291), .B1(new_n320), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n326), .B(KEYINPUT11), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT12), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(new_n282), .B2(G68), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n287), .A2(new_n288), .A3(G68), .ZN(new_n330));
  INV_X1    g0130(.A(new_n282), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(KEYINPUT12), .A3(new_n216), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n327), .A2(new_n329), .A3(new_n330), .A4(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(KEYINPUT75), .A2(G169), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n294), .A2(KEYINPUT3), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT3), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G33), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n335), .A2(new_n337), .A3(G226), .A4(new_n255), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT74), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT74), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n254), .A2(new_n340), .A3(G226), .A4(new_n255), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G33), .A2(G97), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n254), .A2(G232), .A3(G1698), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n339), .A2(new_n341), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n262), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n272), .A2(new_n274), .A3(G45), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n265), .A2(new_n266), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n346), .A2(new_n275), .A3(G238), .A4(new_n347), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n348), .A2(new_n269), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT13), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT13), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n345), .A2(new_n352), .A3(new_n349), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n334), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT14), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n351), .A2(new_n353), .ZN(new_n356));
  INV_X1    g0156(.A(G179), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n354), .A2(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n334), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n356), .A2(new_n355), .A3(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n333), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n278), .A2(G179), .ZN(new_n363));
  INV_X1    g0163(.A(G169), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n278), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n363), .A2(new_n304), .A3(new_n365), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n351), .A2(new_n353), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n333), .B1(new_n367), .B2(G190), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n356), .A2(G200), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n254), .A2(G232), .A3(new_n255), .ZN(new_n371));
  INV_X1    g0171(.A(G107), .ZN(new_n372));
  OAI221_X1 g0172(.A(new_n371), .B1(new_n372), .B2(new_n254), .C1(new_n258), .C2(new_n217), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n262), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n276), .A2(G244), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n374), .A2(new_n269), .A3(new_n375), .ZN(new_n376));
  OR2_X1    g0176(.A1(new_n376), .A2(G179), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n298), .A2(new_n301), .ZN(new_n378));
  XNOR2_X1  g0178(.A(KEYINPUT15), .B(G87), .ZN(new_n379));
  OAI22_X1  g0179(.A1(new_n379), .A2(new_n300), .B1(new_n210), .B2(new_n257), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n291), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g0181(.A(new_n381), .B(KEYINPUT72), .ZN(new_n382));
  MUX2_X1   g0182(.A(new_n282), .B(new_n289), .S(G77), .Z(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n376), .A2(new_n364), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n377), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  OR2_X1    g0186(.A1(new_n376), .A2(new_n279), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n376), .A2(G200), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n387), .A2(new_n382), .A3(new_n383), .A4(new_n388), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n370), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n319), .A2(new_n362), .A3(new_n366), .A4(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT16), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n201), .B1(new_n324), .B2(G58), .ZN(new_n393));
  INV_X1    g0193(.A(G159), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n393), .A2(new_n210), .B1(new_n298), .B2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT7), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n254), .B2(G20), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n336), .A2(G33), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n294), .A2(KEYINPUT3), .ZN(new_n399));
  OAI211_X1 g0199(.A(KEYINPUT7), .B(new_n210), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n216), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n392), .B1(new_n395), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n335), .A2(new_n337), .ZN(new_n403));
  AOI21_X1  g0203(.A(KEYINPUT7), .B1(new_n403), .B2(new_n210), .ZN(new_n404));
  AOI211_X1 g0204(.A(new_n396), .B(G20), .C1(new_n335), .C2(new_n337), .ZN(new_n405));
  OAI21_X1  g0205(.A(G68), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(G58), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n202), .B1(new_n216), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n295), .A2(new_n297), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n408), .A2(G20), .B1(G159), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n406), .A2(new_n410), .A3(KEYINPUT16), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n402), .A2(new_n411), .A3(new_n291), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n287), .A2(new_n282), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n301), .B1(G20), .B2(new_n270), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n413), .B1(new_n414), .B2(KEYINPUT76), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n414), .A2(KEYINPUT76), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n415), .A2(new_n417), .B1(new_n331), .B2(new_n301), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n412), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT18), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n346), .A2(new_n275), .A3(G232), .A4(new_n347), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n269), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n335), .A2(new_n337), .A3(G226), .A4(G1698), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n335), .A2(new_n337), .A3(G223), .A4(new_n255), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G33), .A2(G87), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n262), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n423), .A2(G179), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n428), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(new_n422), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n429), .B1(new_n431), .B2(new_n364), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n419), .A2(new_n420), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n420), .B1(new_n419), .B2(new_n432), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT77), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n414), .A2(KEYINPUT76), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n331), .A2(new_n291), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n301), .ZN(new_n439));
  OAI22_X1  g0239(.A1(new_n438), .A2(new_n416), .B1(new_n282), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n248), .B1(new_n397), .B2(new_n400), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n395), .A2(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n287), .B1(new_n442), .B2(KEYINPUT16), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n440), .B1(new_n443), .B2(new_n402), .ZN(new_n444));
  OAI21_X1  g0244(.A(G169), .B1(new_n430), .B2(new_n422), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n445), .A2(new_n429), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT18), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT77), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n419), .A2(new_n420), .A3(new_n432), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n423), .A2(G190), .A3(new_n428), .ZN(new_n451));
  OAI21_X1  g0251(.A(G200), .B1(new_n430), .B2(new_n422), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n412), .A2(new_n418), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT17), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n452), .A2(new_n451), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n456), .A2(KEYINPUT17), .A3(new_n412), .A4(new_n418), .ZN(new_n457));
  AND2_X1   g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n435), .A2(new_n450), .A3(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n391), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g0260(.A(KEYINPUT5), .B(G41), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n270), .A2(new_n461), .A3(G45), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n462), .A2(new_n347), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(G264), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n254), .A2(G257), .A3(G1698), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n254), .A2(G250), .A3(new_n255), .ZN(new_n466));
  INV_X1    g0266(.A(G294), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n465), .B(new_n466), .C1(new_n294), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n262), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n267), .A2(new_n270), .A3(new_n461), .A4(G45), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n464), .A2(new_n469), .A3(G179), .A4(new_n470), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n471), .A2(KEYINPUT90), .ZN(new_n472));
  AOI22_X1  g0272(.A1(G264), .A2(new_n463), .B1(new_n468), .B2(new_n262), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n364), .B1(new_n473), .B2(new_n470), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n471), .A2(KEYINPUT90), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT91), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n471), .A2(KEYINPUT90), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n471), .A2(KEYINPUT90), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n473), .A2(new_n470), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G169), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n479), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT91), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n331), .A2(new_n372), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT25), .ZN(new_n486));
  XNOR2_X1  g0286(.A(new_n485), .B(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n272), .A2(new_n274), .A3(G33), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n287), .A2(new_n282), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(KEYINPUT78), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT78), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n287), .A2(new_n491), .A3(new_n282), .A4(new_n488), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n490), .A2(G107), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n335), .A2(new_n337), .A3(new_n210), .A4(G87), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT22), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT22), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n254), .A2(new_n498), .A3(new_n210), .A4(G87), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT87), .ZN(new_n501));
  NAND2_X1  g0301(.A1(G33), .A2(G116), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(G20), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n210), .A2(KEYINPUT87), .A3(G33), .A4(G116), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT23), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n210), .B2(G107), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n372), .A2(KEYINPUT23), .A3(G20), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n503), .A2(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n500), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT88), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n500), .A2(KEYINPUT88), .A3(new_n508), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(KEYINPUT24), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT88), .B1(new_n500), .B2(new_n508), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT24), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n287), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n513), .A2(KEYINPUT89), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT89), .B1(new_n513), .B2(new_n516), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n495), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n478), .A2(new_n484), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(G200), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n473), .B2(new_n470), .ZN(new_n522));
  AND4_X1   g0322(.A1(G190), .A2(new_n464), .A3(new_n469), .A4(new_n470), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n495), .B(new_n524), .C1(new_n517), .C2(new_n518), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT79), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G283), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n335), .A2(new_n337), .A3(G250), .A4(G1698), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n335), .A2(new_n337), .A3(G244), .A4(new_n255), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT4), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n529), .B(new_n530), .C1(new_n531), .C2(new_n532), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n531), .A2(new_n532), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n262), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  AND2_X1   g0335(.A1(KEYINPUT5), .A2(G41), .ZN(new_n536));
  NOR2_X1   g0336(.A1(KEYINPUT5), .A2(G41), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(G257), .B(new_n347), .C1(new_n346), .C2(new_n538), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n539), .A2(new_n470), .ZN(new_n540));
  AND4_X1   g0340(.A1(new_n528), .A2(new_n535), .A3(G190), .A4(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT6), .ZN(new_n542));
  AND2_X1   g0342(.A1(G97), .A2(G107), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n542), .B1(new_n543), .B2(new_n204), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n372), .A2(KEYINPUT6), .A3(G97), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(G20), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n409), .A2(G77), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n372), .B1(new_n397), .B2(new_n400), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n291), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n490), .A2(G97), .A3(new_n492), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n282), .A2(G97), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n541), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n521), .B1(new_n535), .B2(new_n540), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n535), .A2(new_n540), .ZN(new_n558));
  OAI22_X1  g0358(.A1(new_n557), .A2(KEYINPUT79), .B1(new_n558), .B2(new_n279), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(G169), .B1(new_n535), .B2(new_n540), .ZN(new_n561));
  OAI21_X1  g0361(.A(G107), .B1(new_n404), .B2(new_n405), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n546), .A2(G20), .B1(G77), .B2(new_n409), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n553), .B1(new_n564), .B2(new_n291), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n561), .B1(new_n565), .B2(new_n552), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n558), .A2(G179), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT80), .ZN(new_n570));
  OAI21_X1  g0370(.A(G274), .B1(new_n261), .B2(new_n283), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n570), .B1(new_n346), .B2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n267), .A2(KEYINPUT80), .A3(new_n270), .A4(G45), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n335), .A2(new_n337), .A3(G238), .A4(new_n255), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n335), .A2(new_n337), .A3(G244), .A4(G1698), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n575), .A2(new_n576), .A3(new_n502), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(new_n262), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n271), .A2(G250), .ZN(new_n579));
  AND4_X1   g0379(.A1(G179), .A2(new_n574), .A3(new_n578), .A4(new_n579), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n572), .A2(new_n573), .B1(new_n271), .B2(G250), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n364), .B1(new_n581), .B2(new_n578), .ZN(new_n582));
  OAI21_X1  g0382(.A(KEYINPUT81), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n574), .A2(new_n578), .A3(new_n579), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(G169), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT81), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n581), .A2(G179), .A3(new_n578), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n379), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n490), .A2(new_n492), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n254), .A2(new_n210), .A3(G68), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT19), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n210), .B1(new_n342), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(G87), .B2(new_n205), .ZN(new_n594));
  INV_X1    g0394(.A(G97), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n592), .B1(new_n300), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n591), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n597), .A2(new_n291), .B1(new_n331), .B2(new_n379), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n590), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n583), .A2(new_n588), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n598), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n490), .A2(G87), .A3(new_n492), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(KEYINPUT82), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT82), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n490), .A2(new_n604), .A3(new_n492), .A4(G87), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n601), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n521), .B1(new_n581), .B2(new_n578), .ZN(new_n607));
  INV_X1    g0407(.A(new_n584), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n607), .B1(G190), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n560), .A2(new_n569), .A3(new_n600), .A4(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n254), .A2(G264), .A3(G1698), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n254), .A2(G257), .A3(new_n255), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n403), .A2(G303), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT83), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n612), .A2(new_n613), .A3(KEYINPUT83), .A4(new_n614), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n617), .A2(new_n262), .A3(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n470), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n620), .B1(new_n463), .B2(G270), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n489), .ZN(new_n623));
  OR3_X1    g0423(.A1(new_n282), .A2(KEYINPUT84), .A3(G116), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT84), .B1(new_n282), .B2(G116), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n623), .A2(G116), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT85), .ZN(new_n627));
  AOI21_X1  g0427(.A(G20), .B1(G33), .B2(G283), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n294), .A2(G97), .ZN(new_n629));
  INV_X1    g0429(.A(G116), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n628), .A2(new_n629), .B1(G20), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(new_n291), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT20), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n627), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n631), .A2(new_n291), .A3(KEYINPUT85), .A4(KEYINPUT20), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n632), .A2(new_n633), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n626), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n622), .A2(new_n638), .A3(G169), .ZN(new_n639));
  NOR2_X1   g0439(.A1(KEYINPUT86), .A2(KEYINPUT21), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n622), .A2(G200), .ZN(new_n642));
  INV_X1    g0442(.A(new_n638), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n619), .A2(G190), .A3(new_n621), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n619), .A2(G179), .A3(new_n621), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n638), .ZN(new_n647));
  INV_X1    g0447(.A(new_n640), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n622), .A2(new_n638), .A3(G169), .A4(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n641), .A2(new_n645), .A3(new_n647), .A4(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n611), .A2(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n460), .A2(new_n527), .A3(new_n651), .ZN(G372));
  INV_X1    g0452(.A(KEYINPUT89), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n500), .A2(KEYINPUT88), .A3(new_n508), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n654), .A2(new_n514), .A3(new_n515), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n509), .A2(new_n510), .A3(new_n515), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n291), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n653), .B1(new_n655), .B2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n513), .A2(KEYINPUT89), .A3(new_n516), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n494), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT93), .B1(new_n660), .B2(new_n476), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT93), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n519), .A2(new_n662), .A3(new_n483), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n641), .A2(new_n647), .A3(new_n649), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n661), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(KEYINPUT92), .B1(new_n580), .B2(new_n582), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT92), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n585), .A2(new_n667), .A3(new_n587), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n669), .A2(new_n599), .B1(new_n606), .B2(new_n609), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n556), .A2(new_n559), .B1(new_n566), .B2(new_n568), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(new_n525), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n665), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n600), .A2(new_n610), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT26), .B1(new_n675), .B2(new_n569), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n669), .A2(new_n599), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT26), .ZN(new_n678));
  INV_X1    g0478(.A(new_n555), .ZN(new_n679));
  NOR3_X1   g0479(.A1(new_n679), .A2(new_n567), .A3(new_n561), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n677), .A2(new_n678), .A3(new_n680), .A4(new_n610), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n676), .A2(new_n677), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n674), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n460), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT94), .ZN(new_n685));
  INV_X1    g0485(.A(new_n366), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n433), .A2(new_n434), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n386), .A2(KEYINPUT95), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT95), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n377), .A2(new_n384), .A3(new_n689), .A4(new_n385), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(KEYINPUT14), .B1(new_n367), .B2(new_n334), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n367), .A2(G179), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(new_n360), .A3(new_n693), .ZN(new_n694));
  AOI22_X1  g0494(.A1(new_n691), .A2(new_n370), .B1(new_n333), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n458), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n687), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n686), .B1(new_n697), .B2(new_n319), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n685), .A2(new_n698), .ZN(G369));
  AND2_X1   g0499(.A1(new_n210), .A2(G13), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n270), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G213), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(G343), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OR3_X1    g0507(.A1(new_n664), .A2(new_n643), .A3(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n643), .A2(new_n707), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n708), .B1(new_n650), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n660), .A2(new_n707), .ZN(new_n713));
  OAI22_X1  g0513(.A1(new_n526), .A2(new_n713), .B1(new_n520), .B2(new_n707), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n706), .B1(new_n661), .B2(new_n663), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n664), .A2(new_n706), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n527), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n715), .A2(new_n717), .A3(new_n719), .ZN(G399));
  INV_X1    g0520(.A(new_n213), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G41), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n205), .A2(G87), .A3(G116), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(G1), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(new_n231), .B2(new_n723), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT28), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n706), .B1(new_n674), .B2(new_n682), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  XOR2_X1   g0529(.A(KEYINPUT96), .B(KEYINPUT29), .Z(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n672), .B1(new_n520), .B2(new_n664), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n680), .A2(new_n600), .A3(new_n610), .A4(new_n678), .ZN(new_n733));
  INV_X1    g0533(.A(new_n610), .ZN(new_n734));
  AOI22_X1  g0534(.A1(new_n666), .A2(new_n668), .B1(new_n598), .B2(new_n590), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n734), .A2(new_n735), .A3(new_n569), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n677), .B(new_n733), .C1(new_n736), .C2(new_n678), .ZN(new_n737));
  OAI211_X1 g0537(.A(KEYINPUT29), .B(new_n707), .C1(new_n732), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n731), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G330), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n651), .A2(new_n520), .A3(new_n525), .A4(new_n707), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n464), .A2(new_n469), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n742), .A2(new_n558), .A3(new_n584), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n743), .A2(new_n646), .A3(KEYINPUT30), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n608), .A2(new_n473), .A3(new_n535), .A4(new_n540), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n619), .A2(G179), .A3(new_n621), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n608), .A2(G179), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n749), .A2(new_n481), .A3(new_n622), .A4(new_n558), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n744), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  AND3_X1   g0551(.A1(new_n751), .A2(KEYINPUT31), .A3(new_n706), .ZN(new_n752));
  AOI21_X1  g0552(.A(KEYINPUT31), .B1(new_n751), .B2(new_n706), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n740), .B1(new_n741), .B2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n739), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n727), .B1(new_n758), .B2(G1), .ZN(G364));
  AOI21_X1  g0559(.A(new_n209), .B1(new_n700), .B2(G45), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n722), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n228), .B1(G20), .B2(new_n364), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n279), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(new_n357), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G97), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n279), .A2(new_n521), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n210), .A2(G179), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G87), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n521), .A2(G190), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n771), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G107), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n769), .A2(new_n774), .A3(new_n778), .A4(new_n254), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n210), .A2(new_n357), .A3(KEYINPUT99), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT99), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(G20), .B2(G179), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n775), .ZN(new_n785));
  NOR2_X1   g0585(.A1(G190), .A2(G200), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n248), .A2(new_n785), .B1(new_n787), .B2(new_n257), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n784), .A2(new_n770), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n779), .B(new_n788), .C1(G50), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n771), .A2(new_n786), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G159), .ZN(new_n794));
  XNOR2_X1  g0594(.A(new_n794), .B(KEYINPUT101), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT32), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT100), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n784), .B2(new_n766), .ZN(new_n798));
  NOR4_X1   g0598(.A1(new_n783), .A2(KEYINPUT100), .A3(new_n279), .A4(G200), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n791), .B(new_n796), .C1(new_n407), .C2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G311), .ZN(new_n802));
  XOR2_X1   g0602(.A(KEYINPUT33), .B(G317), .Z(new_n803));
  OAI22_X1  g0603(.A1(new_n802), .A2(new_n787), .B1(new_n785), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(G326), .B2(new_n790), .ZN(new_n805));
  AOI22_X1  g0605(.A1(G283), .A2(new_n777), .B1(new_n793), .B2(G329), .ZN(new_n806));
  INV_X1    g0606(.A(G303), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n806), .B(new_n403), .C1(new_n807), .C2(new_n772), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n808), .B1(G294), .B2(new_n768), .ZN(new_n809));
  INV_X1    g0609(.A(G322), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n805), .B(new_n809), .C1(new_n810), .C2(new_n800), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n765), .B1(new_n801), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(G13), .A2(G33), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(G20), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n764), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n721), .A2(new_n403), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G355), .A2(new_n817), .B1(new_n630), .B2(new_n721), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n819), .A2(KEYINPUT97), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n213), .A2(new_n403), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n821), .B(KEYINPUT98), .ZN(new_n822));
  INV_X1    g0622(.A(G45), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n822), .B1(new_n232), .B2(new_n268), .C1(new_n252), .C2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n819), .A2(KEYINPUT97), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n820), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n763), .B(new_n812), .C1(new_n816), .C2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n815), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n827), .B1(new_n710), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n710), .A2(G330), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n711), .A2(new_n763), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(G396));
  NOR2_X1   g0632(.A1(new_n764), .A2(new_n813), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G107), .A2(new_n773), .B1(new_n793), .B2(G311), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n777), .A2(G87), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n835), .A2(new_n403), .A3(new_n769), .A4(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n787), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n838), .A2(G116), .B1(new_n790), .B2(G303), .ZN(new_n839));
  XOR2_X1   g0639(.A(KEYINPUT102), .B(G283), .Z(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n785), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n800), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n837), .B(new_n841), .C1(G294), .C2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(G137), .ZN(new_n844));
  OAI22_X1  g0644(.A1(new_n844), .A2(new_n789), .B1(new_n785), .B2(new_n299), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n845), .B(KEYINPUT103), .Z(new_n846));
  INV_X1    g0646(.A(G143), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n846), .B1(new_n847), .B2(new_n800), .C1(new_n394), .C2(new_n787), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT34), .ZN(new_n849));
  AOI22_X1  g0649(.A1(G50), .A2(new_n773), .B1(new_n793), .B2(G132), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n777), .A2(G68), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n850), .A2(new_n254), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(G58), .B2(new_n768), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n843), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n762), .B1(G77), .B2(new_n834), .C1(new_n854), .C2(new_n765), .ZN(new_n855));
  OR2_X1    g0655(.A1(new_n855), .A2(KEYINPUT104), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(KEYINPUT104), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n384), .A2(new_n706), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n688), .A2(new_n690), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n389), .A2(new_n386), .A3(new_n858), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  OAI211_X1 g0662(.A(new_n856), .B(new_n857), .C1(new_n814), .C2(new_n862), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n860), .A2(new_n861), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n729), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n728), .A2(new_n862), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n755), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT106), .ZN(new_n868));
  OR2_X1    g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n867), .A2(new_n868), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n869), .A2(new_n763), .A3(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n865), .A2(new_n755), .A3(new_n866), .ZN(new_n872));
  XNOR2_X1  g0672(.A(new_n872), .B(KEYINPUT105), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n863), .B1(new_n871), .B2(new_n873), .ZN(G384));
  OAI211_X1 g0674(.A(new_n229), .B(G116), .C1(KEYINPUT35), .C2(new_n546), .ZN(new_n875));
  OR2_X1    g0675(.A1(new_n875), .A2(KEYINPUT107), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n546), .A2(KEYINPUT35), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n875), .A2(KEYINPUT107), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT36), .Z(new_n880));
  INV_X1    g0680(.A(new_n231), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n881), .B(G77), .C1(new_n407), .C2(new_n216), .ZN(new_n882));
  AOI211_X1 g0682(.A(G13), .B(new_n270), .C1(new_n882), .C2(new_n247), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n386), .A2(new_n706), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n866), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n442), .A2(KEYINPUT16), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n411), .A2(new_n291), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n418), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n704), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n459), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n419), .A2(new_n432), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n419), .A2(new_n891), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT37), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n895), .A2(new_n896), .A3(new_n897), .A4(new_n453), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n890), .A2(new_n432), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n899), .A2(new_n892), .A3(new_n453), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n898), .B1(new_n900), .B2(new_n897), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n894), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT38), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n901), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n362), .A2(KEYINPUT108), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT108), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n694), .A2(new_n908), .A3(new_n333), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n333), .A2(new_n706), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n911), .B1(new_n369), .B2(new_n368), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n907), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n370), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n911), .B1(new_n914), .B2(new_n694), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n887), .A2(new_n906), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n895), .A2(new_n896), .A3(new_n453), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT37), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n447), .A2(new_n449), .A3(new_n455), .A4(new_n457), .ZN(new_n920));
  INV_X1    g0720(.A(new_n896), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n898), .A2(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT109), .B1(new_n922), .B2(KEYINPUT38), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT109), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n919), .A2(new_n898), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n896), .B1(new_n458), .B2(new_n687), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n924), .B(new_n903), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n923), .A2(new_n905), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT39), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n706), .B1(new_n907), .B2(new_n909), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n904), .A2(KEYINPUT39), .A3(new_n905), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n704), .B1(new_n433), .B2(new_n434), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n917), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n731), .A2(new_n460), .A3(new_n738), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n698), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n935), .B(new_n937), .Z(new_n938));
  INV_X1    g0738(.A(KEYINPUT40), .ZN(new_n939));
  AND3_X1   g0739(.A1(new_n894), .A2(KEYINPUT38), .A3(new_n901), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT38), .B1(new_n894), .B2(new_n901), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n864), .B1(new_n741), .B2(new_n754), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n916), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n939), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n928), .A2(KEYINPUT40), .A3(new_n916), .A4(new_n943), .ZN(new_n946));
  AND2_X1   g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI211_X1 g0747(.A(new_n459), .B(new_n391), .C1(new_n741), .C2(new_n754), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n949), .A2(new_n950), .A3(new_n740), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n938), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n270), .B2(new_n700), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT110), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n953), .A2(new_n954), .B1(new_n938), .B2(new_n951), .ZN(new_n955));
  AND2_X1   g0755(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n884), .B1(new_n955), .B2(new_n956), .ZN(G367));
  OAI21_X1  g0757(.A(new_n671), .B1(new_n679), .B2(new_n707), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n680), .A2(new_n706), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NOR3_X1   g0761(.A1(new_n526), .A2(new_n664), .A3(new_n706), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n961), .B1(new_n962), .B2(new_n716), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT44), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g0765(.A(KEYINPUT44), .B(new_n961), .C1(new_n962), .C2(new_n716), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n719), .A2(new_n717), .A3(new_n960), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT45), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n719), .A2(KEYINPUT45), .A3(new_n717), .A4(new_n960), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AND3_X1   g0772(.A1(new_n967), .A2(new_n972), .A3(new_n715), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n715), .B1(new_n967), .B2(new_n972), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n719), .B1(new_n714), .B2(new_n718), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(new_n711), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n757), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n757), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n722), .B(KEYINPUT41), .Z(new_n980));
  OAI21_X1  g0780(.A(new_n760), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  OR3_X1    g0781(.A1(new_n719), .A2(KEYINPUT42), .A3(new_n961), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n569), .B1(new_n520), .B2(new_n958), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n983), .A2(new_n707), .ZN(new_n984));
  OAI21_X1  g0784(.A(KEYINPUT42), .B1(new_n719), .B2(new_n961), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n982), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n677), .B(new_n610), .C1(new_n606), .C2(new_n707), .ZN(new_n987));
  INV_X1    g0787(.A(new_n606), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n735), .A2(new_n988), .A3(new_n706), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n987), .A2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n986), .A2(new_n992), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT111), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n715), .A2(new_n961), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n986), .A2(new_n995), .A3(new_n992), .ZN(new_n999));
  AND3_X1   g0799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n998), .B1(new_n997), .B2(new_n999), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n990), .A2(new_n815), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n822), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n816), .B1(new_n213), .B2(new_n379), .C1(new_n1004), .C2(new_n241), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(new_n762), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n467), .A2(new_n785), .B1(new_n787), .B2(new_n840), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n789), .A2(new_n802), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n773), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT46), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n772), .B2(new_n630), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n768), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1009), .B(new_n1011), .C1(new_n372), .C2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(G317), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n403), .B1(new_n792), .B2(new_n1014), .C1(new_n595), .C2(new_n776), .ZN(new_n1015));
  NOR4_X1   g0815(.A1(new_n1007), .A2(new_n1008), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n807), .B2(new_n800), .ZN(new_n1017));
  XNOR2_X1  g0817(.A(new_n1017), .B(KEYINPUT112), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n246), .A2(new_n787), .B1(new_n789), .B2(new_n847), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n785), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1019), .B1(G159), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n254), .B1(new_n776), .B2(new_n257), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n772), .A2(new_n407), .B1(new_n792), .B2(new_n844), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1022), .B(new_n1023), .C1(G68), .C2(new_n768), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1021), .B(new_n1024), .C1(new_n299), .C2(new_n800), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1018), .A2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT47), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1006), .B1(new_n1027), .B2(new_n764), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n981), .A2(new_n1002), .B1(new_n1003), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(G387));
  INV_X1    g0830(.A(new_n268), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n822), .B1(new_n238), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n817), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1032), .B1(new_n724), .B2(new_n1033), .ZN(new_n1034));
  OR3_X1    g0834(.A1(new_n301), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1035));
  OAI21_X1  g0835(.A(KEYINPUT50), .B1(new_n301), .B2(G50), .ZN(new_n1036));
  AOI21_X1  g0836(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1035), .A2(new_n724), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n1034), .A2(new_n1038), .B1(new_n372), .B2(new_n721), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n816), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n762), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n248), .A2(new_n787), .B1(new_n789), .B2(new_n394), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n439), .B2(new_n1020), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n773), .A2(G77), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n299), .B2(new_n792), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1012), .A2(new_n379), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n254), .B1(new_n776), .B2(new_n595), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1043), .B(new_n1048), .C1(new_n246), .C2(new_n800), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n793), .A2(G326), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n254), .B1(new_n777), .B2(G116), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1012), .A2(new_n840), .B1(new_n772), .B2(new_n467), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G311), .A2(new_n1020), .B1(new_n790), .B2(G322), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n807), .B2(new_n787), .C1(new_n1014), .C2(new_n800), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT48), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1052), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n1055), .B2(new_n1054), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT49), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n1050), .B(new_n1051), .C1(new_n1057), .C2(new_n1058), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1049), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1041), .B1(new_n1061), .B2(new_n764), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n714), .B2(new_n828), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n722), .B1(new_n757), .B2(new_n977), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n757), .A2(new_n977), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1063), .B1(new_n760), .B2(new_n977), .C1(new_n1064), .C2(new_n1065), .ZN(G393));
  NAND2_X1  g0866(.A1(new_n961), .A2(new_n815), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n816), .B1(new_n595), .B2(new_n213), .C1(new_n1004), .C2(new_n245), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(new_n762), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n800), .A2(new_n802), .B1(new_n1014), .B2(new_n789), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT52), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n840), .A2(new_n772), .B1(new_n792), .B2(new_n810), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n778), .A2(new_n403), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1072), .B(new_n1073), .C1(G116), .C2(new_n768), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n838), .A2(G294), .B1(new_n1020), .B2(G303), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1071), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n800), .A2(new_n394), .B1(new_n299), .B2(new_n789), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT51), .Z(new_n1078));
  AOI22_X1  g0878(.A1(new_n838), .A2(new_n439), .B1(new_n1020), .B2(G50), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n324), .A2(new_n773), .B1(new_n793), .B2(G143), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n1080), .A2(new_n254), .A3(new_n836), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1079), .B(new_n1081), .C1(new_n257), .C2(new_n1012), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1076), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1069), .B1(new_n1083), .B2(new_n764), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n975), .A2(new_n761), .B1(new_n1067), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n974), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n967), .A2(new_n972), .A3(new_n715), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1086), .A2(new_n978), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n722), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n975), .A2(new_n978), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1085), .B1(new_n1089), .B2(new_n1090), .ZN(G390));
  NAND2_X1  g0891(.A1(new_n755), .A2(new_n862), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n916), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT114), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n755), .A2(new_n916), .A3(new_n862), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1092), .A2(KEYINPUT114), .A3(new_n1093), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1097), .A2(new_n887), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1096), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n707), .B(new_n862), .C1(new_n732), .C2(new_n737), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(new_n886), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n755), .A2(KEYINPUT115), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n862), .B1(new_n755), .B2(KEYINPUT115), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1093), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1099), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n460), .A2(new_n755), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n936), .A2(new_n698), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1102), .A2(new_n916), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n931), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1113), .A2(new_n1114), .A3(new_n1115), .A4(new_n928), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n928), .A2(new_n1115), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1101), .A2(new_n886), .B1(new_n913), .B2(new_n915), .ZN(new_n1118));
  OAI21_X1  g0918(.A(KEYINPUT113), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n885), .B1(new_n728), .B2(new_n862), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1115), .B1(new_n1121), .B2(new_n1093), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n930), .A2(new_n932), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1120), .A2(new_n1124), .A3(new_n1096), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1096), .B1(new_n1120), .B2(new_n1124), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1112), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n928), .A2(new_n1115), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1114), .B1(new_n1128), .B2(new_n1113), .ZN(new_n1129));
  NOR3_X1   g0929(.A1(new_n1117), .A2(new_n1118), .A3(KEYINPUT113), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1124), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n1100), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1120), .A2(new_n1124), .A3(new_n1096), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1110), .B1(new_n1099), .B2(new_n1107), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1132), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1127), .A2(new_n1135), .A3(new_n722), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n793), .A2(G294), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n774), .A2(new_n851), .A3(new_n1137), .A4(new_n403), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n838), .A2(G97), .B1(new_n1020), .B2(G107), .ZN(new_n1139));
  INV_X1    g0939(.A(G283), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1139), .B1(new_n1140), .B2(new_n789), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1138), .B(new_n1141), .C1(G77), .C2(new_n768), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n842), .A2(G116), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n842), .A2(G132), .ZN(new_n1144));
  INV_X1    g0944(.A(G128), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT54), .B(G143), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n1145), .A2(new_n789), .B1(new_n787), .B2(new_n1146), .ZN(new_n1147));
  OR3_X1    g0947(.A1(new_n772), .A2(KEYINPUT53), .A3(new_n299), .ZN(new_n1148));
  OAI21_X1  g0948(.A(KEYINPUT53), .B1(new_n772), .B2(new_n299), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1148), .B(new_n1149), .C1(new_n394), .C2(new_n1012), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n785), .A2(new_n844), .ZN(new_n1151));
  INV_X1    g0951(.A(G125), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n254), .B1(new_n792), .B2(new_n1152), .C1(new_n246), .C2(new_n776), .ZN(new_n1153));
  NOR4_X1   g0953(.A1(new_n1147), .A2(new_n1150), .A3(new_n1151), .A4(new_n1153), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1142), .A2(new_n1143), .B1(new_n1144), .B2(new_n1154), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n762), .B1(new_n439), .B2(new_n834), .C1(new_n1155), .C2(new_n765), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n1123), .B2(new_n813), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n761), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n1136), .A2(new_n1159), .A3(KEYINPUT116), .ZN(new_n1160));
  AOI21_X1  g0960(.A(KEYINPUT116), .B1(new_n1136), .B2(new_n1159), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(G378));
  NAND2_X1  g0962(.A1(new_n319), .A2(new_n366), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n308), .A2(new_n704), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1164), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n319), .A2(new_n366), .A3(new_n1166), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1165), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1168), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1166), .B1(new_n319), .B2(new_n366), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n686), .B(new_n1164), .C1(new_n314), .C2(new_n318), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n1169), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(new_n813), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n762), .B1(new_n834), .B2(G50), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G58), .A2(new_n777), .B1(new_n793), .B2(G283), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n254), .A2(G41), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1177), .A2(new_n1044), .A3(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n838), .A2(new_n589), .B1(new_n790), .B2(G116), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n595), .B2(new_n785), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1179), .B(new_n1181), .C1(G68), .C2(new_n768), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT117), .B1(new_n842), .B2(G107), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n842), .A2(KEYINPUT117), .A3(G107), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1182), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT58), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n838), .A2(G137), .B1(new_n790), .B2(G125), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1020), .A2(G132), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1146), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G150), .A2(new_n768), .B1(new_n773), .B2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1188), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G128), .B2(new_n842), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n777), .A2(G159), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT118), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1198), .A2(G124), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(G124), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n793), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(G33), .A2(G41), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1196), .A2(new_n1197), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n246), .B1(G33), .B2(G41), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1187), .B1(new_n1195), .B2(new_n1203), .C1(new_n1178), .C2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1176), .B1(new_n1205), .B2(new_n764), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1175), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n935), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n945), .A2(G330), .A3(new_n946), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n1174), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1169), .A2(new_n1173), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1212), .A2(new_n945), .A3(G330), .A4(new_n946), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1209), .B1(new_n1214), .B2(KEYINPUT119), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1211), .A2(new_n1213), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT119), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1216), .A2(new_n1217), .A3(new_n935), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1215), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1208), .B1(new_n1219), .B2(new_n761), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT57), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n935), .A2(KEYINPUT120), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT120), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n917), .A2(new_n933), .A3(new_n1224), .A4(new_n934), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1214), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1216), .A2(new_n1225), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1222), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1135), .A2(new_n1111), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n723), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1219), .A2(new_n1230), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1231), .A2(KEYINPUT121), .B1(new_n1232), .B2(new_n1222), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1230), .A2(new_n1234), .A3(KEYINPUT57), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1235), .A2(new_n722), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT121), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1221), .B1(new_n1233), .B2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(G375));
  OAI21_X1  g1040(.A(new_n762), .B1(new_n834), .B2(G68), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n299), .A2(new_n787), .B1(new_n785), .B2(new_n1146), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G132), .B2(new_n790), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n254), .B1(new_n776), .B2(new_n407), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n772), .A2(new_n394), .B1(new_n792), .B2(new_n1145), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1244), .B(new_n1245), .C1(G50), .C2(new_n768), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1243), .B(new_n1246), .C1(new_n844), .C2(new_n800), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n838), .A2(G107), .B1(new_n1020), .B2(G116), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT123), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1046), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n790), .A2(G294), .ZN(new_n1252));
  OAI22_X1  g1052(.A1(new_n772), .A2(new_n595), .B1(new_n792), .B2(new_n807), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n254), .B(new_n1253), .C1(G77), .C2(new_n777), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1250), .A2(new_n1251), .A3(new_n1252), .A4(new_n1254), .ZN(new_n1255));
  OAI22_X1  g1055(.A1(new_n1248), .A2(new_n1249), .B1(new_n1140), .B2(new_n800), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1247), .B1(new_n1255), .B2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1241), .B1(new_n1257), .B2(new_n764), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n916), .B2(new_n814), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1108), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n760), .B(KEYINPUT122), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1259), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1134), .A2(new_n980), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1260), .A2(new_n1110), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1262), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(G381));
  NOR2_X1   g1066(.A1(G393), .A2(G396), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(G390), .A2(G384), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1029), .A2(new_n1265), .A3(new_n1267), .A4(new_n1268), .ZN(new_n1269));
  XOR2_X1   g1069(.A(new_n1269), .B(KEYINPUT124), .Z(new_n1270));
  NAND2_X1  g1070(.A1(new_n1136), .A2(new_n1159), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1270), .A2(new_n1272), .A3(new_n1239), .ZN(G407));
  INV_X1    g1073(.A(G213), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1274), .A2(G343), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1239), .A2(new_n1272), .A3(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(G407), .A2(G213), .A3(new_n1276), .ZN(G409));
  INV_X1    g1077(.A(KEYINPUT60), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1264), .B1(new_n1278), .B2(new_n1134), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1108), .A2(new_n1111), .A3(new_n1278), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1280), .A2(new_n723), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1262), .B1(new_n1279), .B2(new_n1281), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1282), .A2(G384), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1282), .A2(G384), .ZN(new_n1284));
  AND2_X1   g1084(.A1(new_n1275), .A2(G2897), .ZN(new_n1285));
  AND3_X1   g1085(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1285), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1216), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1216), .A2(new_n1225), .ZN(new_n1290));
  OAI21_X1  g1090(.A(KEYINPUT57), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1110), .B1(new_n1158), .B2(new_n1108), .ZN(new_n1292));
  OAI211_X1 g1092(.A(KEYINPUT121), .B(new_n722), .C1(new_n1291), .C2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1218), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n935), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1222), .B1(new_n1296), .B2(new_n1292), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1293), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT121), .B1(new_n1235), .B2(new_n722), .ZN(new_n1299));
  OAI211_X1 g1099(.A(G378), .B(new_n1220), .C1(new_n1298), .C2(new_n1299), .ZN(new_n1300));
  OR3_X1    g1100(.A1(new_n1296), .A2(new_n1292), .A3(new_n980), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1261), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1208), .B1(new_n1234), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1301), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1272), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1275), .B1(new_n1300), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT125), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1288), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1271), .B1(new_n1301), .B2(new_n1303), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1309), .B1(new_n1239), .B2(G378), .ZN(new_n1310));
  OAI21_X1  g1110(.A(KEYINPUT125), .B1(new_n1310), .B2(new_n1275), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1308), .A2(new_n1311), .ZN(new_n1312));
  AND2_X1   g1112(.A1(G393), .A2(G396), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1313), .A2(new_n1267), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n980), .B1(new_n1088), .B2(new_n758), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1002), .B1(new_n1315), .B2(new_n761), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1028), .A2(new_n1003), .ZN(new_n1317));
  AND3_X1   g1117(.A1(new_n1316), .A2(new_n1317), .A3(G390), .ZN(new_n1318));
  AOI21_X1  g1118(.A(G390), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1314), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT126), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(KEYINPUT127), .B1(new_n1029), .B2(G390), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT127), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1319), .A2(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1314), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1029), .A2(G390), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1323), .A2(new_n1325), .A3(new_n1326), .A4(new_n1327), .ZN(new_n1328));
  OAI211_X1 g1128(.A(KEYINPUT126), .B(new_n1314), .C1(new_n1318), .C2(new_n1319), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1322), .A2(new_n1328), .A3(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT61), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1330), .A2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1300), .A2(new_n1305), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1275), .ZN(new_n1334));
  AND2_X1   g1134(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1333), .A2(new_n1334), .A3(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT63), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1332), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1306), .A2(KEYINPUT63), .A3(new_n1335), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1312), .A2(new_n1338), .A3(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT62), .ZN(new_n1341));
  AND3_X1   g1141(.A1(new_n1306), .A2(new_n1341), .A3(new_n1335), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1331), .B1(new_n1306), .B2(new_n1288), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1341), .B1(new_n1306), .B2(new_n1335), .ZN(new_n1344));
  NOR3_X1   g1144(.A1(new_n1342), .A2(new_n1343), .A3(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1340), .B1(new_n1345), .B2(new_n1330), .ZN(G405));
  OAI21_X1  g1146(.A(new_n1300), .B1(new_n1239), .B2(new_n1271), .ZN(new_n1347));
  OR2_X1    g1147(.A1(new_n1347), .A2(new_n1335), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1330), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1347), .A2(new_n1335), .ZN(new_n1350));
  AND3_X1   g1150(.A1(new_n1348), .A2(new_n1349), .A3(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1349), .B1(new_n1348), .B2(new_n1350), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(new_n1351), .A2(new_n1352), .ZN(G402));
endmodule


