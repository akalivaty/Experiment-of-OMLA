//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G128), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G119), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G128), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n191), .A2(KEYINPUT23), .A3(G119), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G110), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(new_n192), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT24), .B(G110), .ZN(new_n201));
  OR2_X1    g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G140), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G125), .ZN(new_n204));
  INV_X1    g018(.A(G125), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G140), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT16), .ZN(new_n207));
  OR3_X1    g021(.A1(new_n205), .A2(KEYINPUT16), .A3(G140), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n208), .A3(G146), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(G146), .B1(new_n207), .B2(new_n208), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n199), .B(new_n202), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(new_n212), .B(KEYINPUT77), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT79), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n209), .B(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n204), .A2(new_n206), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n216), .A2(G146), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n200), .A2(new_n201), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n218), .B1(new_n198), .B2(G110), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT78), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n217), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n215), .B(new_n221), .C1(new_n220), .C2(new_n219), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n213), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G953), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G953), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(G221), .A3(G234), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT22), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n229), .B(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G137), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n231), .B(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n223), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n213), .A2(new_n233), .A3(new_n222), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n188), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT25), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n235), .A2(KEYINPUT25), .A3(new_n188), .A4(new_n236), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n190), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n235), .A2(new_n236), .ZN(new_n242));
  NOR3_X1   g056(.A1(new_n242), .A2(G902), .A3(new_n189), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT80), .ZN(new_n245));
  XNOR2_X1  g059(.A(new_n244), .B(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G143), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(G146), .ZN(new_n248));
  INV_X1    g062(.A(G146), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT64), .B1(new_n249), .B2(G143), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT64), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(new_n247), .A3(G146), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n248), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n249), .A2(G143), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n247), .A2(G146), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n253), .A2(new_n255), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n232), .A2(KEYINPUT11), .A3(G134), .ZN(new_n262));
  INV_X1    g076(.A(G134), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G137), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT11), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n266), .B1(new_n263), .B2(G137), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT65), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n232), .A2(G134), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT65), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n270), .A3(new_n266), .ZN(new_n271));
  AOI211_X1 g085(.A(G131), .B(new_n265), .C1(new_n268), .C2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G131), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n268), .A2(new_n271), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n262), .A2(new_n264), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n261), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n195), .A2(G116), .ZN(new_n278));
  INV_X1    g092(.A(G116), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G119), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(KEYINPUT2), .B(G113), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n281), .B(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n191), .B1(new_n258), .B2(KEYINPUT1), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n253), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT1), .ZN(new_n287));
  OAI21_X1  g101(.A(G128), .B1(new_n248), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n260), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n274), .A2(new_n273), .A3(new_n275), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n269), .A2(new_n264), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G131), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n290), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n277), .A2(new_n284), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(G237), .B1(new_n225), .B2(new_n227), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G210), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT26), .B(G101), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n296), .A2(G210), .A3(new_n298), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n301), .B1(new_n300), .B2(new_n302), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n295), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT68), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT30), .ZN(new_n308));
  AND3_X1   g122(.A1(new_n290), .A2(new_n291), .A3(new_n293), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n257), .A2(new_n260), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n250), .A2(new_n252), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n258), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n310), .B1(new_n312), .B2(new_n254), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n270), .B1(new_n269), .B2(new_n266), .ZN(new_n314));
  AOI211_X1 g128(.A(KEYINPUT65), .B(KEYINPUT11), .C1(new_n232), .C2(G134), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n275), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G131), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n313), .B1(new_n317), .B2(new_n291), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n308), .B1(new_n309), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n277), .A2(KEYINPUT30), .A3(new_n294), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n283), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT31), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT68), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n295), .A2(new_n323), .A3(new_n305), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n307), .A2(new_n321), .A3(new_n322), .A4(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT69), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n307), .A2(new_n321), .A3(new_n324), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT31), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n326), .A3(KEYINPUT31), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n283), .B1(new_n309), .B2(new_n318), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT71), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(new_n333), .A3(new_n295), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT28), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n284), .B1(new_n277), .B2(new_n294), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n335), .B1(new_n336), .B2(KEYINPUT71), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n334), .A2(new_n337), .B1(new_n335), .B2(new_n295), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n305), .B(KEYINPUT70), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT72), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n295), .A2(new_n335), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n277), .A2(new_n284), .A3(new_n294), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n342), .A2(new_n336), .A3(KEYINPUT71), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT28), .B1(new_n332), .B2(new_n333), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n341), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT72), .ZN(new_n346));
  INV_X1    g160(.A(new_n339), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n330), .A2(new_n331), .A3(new_n340), .A4(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(G472), .A2(G902), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  XOR2_X1   g165(.A(KEYINPUT73), .B(KEYINPUT32), .Z(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT74), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT74), .ZN(new_n355));
  AOI211_X1 g169(.A(new_n355), .B(new_n352), .C1(new_n349), .C2(new_n350), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n350), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n328), .A2(new_n326), .A3(KEYINPUT31), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n359), .B1(new_n329), .B2(new_n327), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n348), .A2(new_n340), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n358), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n341), .B(new_n339), .C1(new_n343), .C2(new_n344), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT29), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n321), .A2(new_n295), .ZN(new_n365));
  INV_X1    g179(.A(new_n305), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n363), .A2(new_n364), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT75), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT28), .B1(new_n342), .B2(new_n336), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n371), .A2(KEYINPUT29), .A3(new_n305), .A4(new_n341), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT76), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n372), .B(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n363), .A2(new_n367), .A3(KEYINPUT75), .A4(new_n364), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n370), .A2(new_n374), .A3(new_n188), .A4(new_n375), .ZN(new_n376));
  AOI22_X1  g190(.A1(new_n362), .A2(KEYINPUT32), .B1(new_n376), .B2(G472), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n246), .B1(new_n357), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n317), .A2(new_n291), .ZN(new_n379));
  INV_X1    g193(.A(G104), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G107), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n380), .A2(G107), .ZN(new_n383));
  OAI21_X1  g197(.A(G101), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT3), .B1(new_n380), .B2(G107), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT3), .ZN(new_n386));
  INV_X1    g200(.A(G107), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n387), .A3(G104), .ZN(new_n388));
  INV_X1    g202(.A(G101), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n385), .A2(new_n388), .A3(new_n389), .A4(new_n381), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n384), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n290), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n312), .A2(new_n288), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n391), .B1(new_n394), .B2(new_n286), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n379), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT12), .ZN(new_n397));
  INV_X1    g211(.A(new_n286), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n253), .A2(new_n285), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n392), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n379), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n290), .A2(new_n392), .A3(KEYINPUT10), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n385), .A2(new_n388), .A3(new_n381), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G101), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT4), .A3(new_n390), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT4), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n406), .A2(new_n409), .A3(G101), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n261), .A3(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n403), .A2(new_n404), .A3(new_n405), .A4(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT12), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n379), .B(new_n413), .C1(new_n393), .C2(new_n395), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n397), .A2(new_n412), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT83), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT81), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n228), .A2(new_n417), .A3(G227), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n417), .B1(new_n228), .B2(G227), .ZN(new_n420));
  OAI21_X1  g234(.A(G110), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n420), .ZN(new_n422));
  INV_X1    g236(.A(G110), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(new_n418), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n421), .A2(new_n424), .A3(G140), .ZN(new_n425));
  AOI21_X1  g239(.A(G140), .B1(new_n421), .B2(new_n424), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n397), .A2(new_n412), .A3(new_n429), .A4(new_n414), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n416), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n405), .B(new_n411), .C1(new_n395), .C2(new_n401), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n379), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n427), .A3(new_n412), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G469), .ZN(new_n436));
  INV_X1    g250(.A(G469), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n415), .A2(new_n428), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n427), .B1(new_n433), .B2(new_n412), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n437), .B(new_n188), .C1(new_n438), .C2(new_n439), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n437), .A2(new_n188), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n436), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n408), .A2(new_n283), .A3(new_n410), .ZN(new_n445));
  OR2_X1    g259(.A1(new_n281), .A2(new_n282), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n278), .A2(new_n280), .A3(KEYINPUT5), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n447), .B(G113), .C1(KEYINPUT5), .C2(new_n278), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n392), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(G110), .B(G122), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT85), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n451), .B(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n445), .A2(new_n449), .A3(new_n453), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n455), .A2(KEYINPUT6), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n450), .A2(new_n458), .A3(new_n454), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n286), .A2(new_n205), .A3(new_n289), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n462), .B1(new_n205), .B2(new_n261), .ZN(new_n463));
  INV_X1    g277(.A(G224), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(G953), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n463), .B(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(G902), .B1(new_n461), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n463), .A2(new_n465), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT7), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n448), .A2(new_n446), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n391), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n449), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n453), .B(KEYINPUT8), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT86), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT7), .B1(new_n464), .B2(G953), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n463), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n475), .B1(new_n463), .B2(new_n476), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n469), .B(new_n474), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT87), .ZN(new_n481));
  INV_X1    g295(.A(new_n479), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n477), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT87), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n483), .A2(new_n484), .A3(new_n469), .A4(new_n474), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n481), .A2(new_n485), .A3(new_n456), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n467), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G210), .B1(G237), .B2(G902), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n467), .A2(new_n486), .A3(new_n488), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n224), .A2(G952), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n493), .B1(G234), .B2(G237), .ZN(new_n494));
  INV_X1    g308(.A(new_n228), .ZN(new_n495));
  NAND2_X1  g309(.A1(G234), .A2(G237), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(G902), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  XOR2_X1   g312(.A(KEYINPUT21), .B(G898), .Z(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n494), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT9), .B(G234), .Z(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n188), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n504), .A2(G221), .ZN(new_n505));
  OAI21_X1  g319(.A(G214), .B1(G237), .B2(G902), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  OR2_X1    g321(.A1(new_n507), .A2(KEYINPUT84), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(KEYINPUT84), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n502), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n444), .A2(new_n492), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT89), .ZN(new_n514));
  INV_X1    g328(.A(G122), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n514), .B1(new_n515), .B2(G116), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n279), .A2(KEYINPUT89), .A3(G122), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n518), .B1(new_n279), .B2(G122), .ZN(new_n519));
  OR2_X1    g333(.A1(new_n519), .A2(G107), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT90), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n521), .B1(new_n191), .B2(G143), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n247), .A2(KEYINPUT90), .A3(G128), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n191), .A2(G143), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G134), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n524), .A2(new_n263), .A3(new_n525), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT93), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(new_n518), .B2(KEYINPUT14), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT14), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT93), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n532), .B1(new_n516), .B2(new_n517), .ZN(new_n535));
  OAI22_X1  g349(.A1(new_n535), .A2(KEYINPUT92), .B1(new_n279), .B2(G122), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n535), .A2(KEYINPUT92), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n520), .B(new_n529), .C1(new_n538), .C2(new_n387), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT13), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n524), .A2(new_n540), .B1(new_n191), .B2(G143), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n541), .B1(new_n540), .B2(new_n524), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G134), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n519), .B(G107), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n528), .A2(KEYINPUT91), .ZN(new_n545));
  OR2_X1    g359(.A1(new_n528), .A2(KEYINPUT91), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n543), .A2(new_n544), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n539), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n503), .A2(G217), .A3(new_n224), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(KEYINPUT94), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n550), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n539), .A2(new_n552), .A3(new_n547), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(KEYINPUT95), .A3(new_n553), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n539), .A2(new_n547), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT95), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n556), .A3(new_n552), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n554), .A2(new_n188), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(G478), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(KEYINPUT15), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n560), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n554), .A2(new_n188), .A3(new_n557), .A4(new_n562), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n561), .A2(KEYINPUT96), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(KEYINPUT96), .B1(new_n561), .B2(new_n563), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n296), .A2(G143), .A3(G214), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(G143), .B1(new_n296), .B2(G214), .ZN(new_n568));
  OAI21_X1  g382(.A(G131), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT17), .ZN(new_n570));
  INV_X1    g384(.A(G237), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n228), .A2(G214), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n247), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(new_n273), .A3(new_n566), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n569), .A2(new_n570), .A3(new_n574), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n210), .A2(new_n211), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n273), .B1(new_n573), .B2(new_n566), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT17), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n575), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n216), .B(G146), .ZN(new_n581));
  NAND2_X1  g395(.A1(KEYINPUT18), .A2(G131), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n573), .A2(new_n566), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT18), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n581), .B(new_n583), .C1(new_n569), .C2(new_n584), .ZN(new_n585));
  XOR2_X1   g399(.A(G113), .B(G122), .Z(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT88), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(new_n380), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n580), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n588), .B1(new_n580), .B2(new_n585), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n188), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(G475), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT20), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n216), .A2(KEYINPUT19), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT19), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(new_n204), .B2(new_n206), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n249), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n573), .A2(new_n273), .A3(new_n566), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n215), .B(new_n599), .C1(new_n600), .C2(new_n578), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n585), .ZN(new_n602));
  INV_X1    g416(.A(new_n588), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n589), .ZN(new_n605));
  INV_X1    g419(.A(G475), .ZN(new_n606));
  AND4_X1   g420(.A1(new_n594), .A2(new_n605), .A3(new_n606), .A4(new_n188), .ZN(new_n607));
  AOI21_X1  g421(.A(G475), .B1(new_n604), .B2(new_n589), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n594), .B1(new_n608), .B2(new_n188), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n593), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n564), .A2(new_n565), .A3(new_n610), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n513), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n378), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT97), .B(G101), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(G3));
  AOI21_X1  g429(.A(new_n505), .B1(new_n436), .B2(new_n443), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n349), .A2(new_n188), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(G472), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n351), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n246), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n553), .A2(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n552), .B1(new_n539), .B2(new_n547), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n555), .A2(new_n621), .A3(new_n552), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT33), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n554), .A2(new_n627), .A3(new_n557), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n559), .A2(G902), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n626), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n558), .A2(new_n559), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT99), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n632), .A2(new_n633), .A3(new_n610), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n633), .B1(new_n632), .B2(new_n610), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n467), .A2(new_n486), .A3(new_n488), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n488), .B1(new_n467), .B2(new_n486), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n639), .A2(new_n501), .A3(new_n507), .ZN(new_n640));
  AOI21_X1  g454(.A(KEYINPUT100), .B1(new_n636), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n632), .A2(new_n610), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT99), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n632), .A2(new_n633), .A3(new_n610), .ZN(new_n644));
  AND4_X1   g458(.A1(KEYINPUT100), .A2(new_n643), .A3(new_n640), .A4(new_n644), .ZN(new_n645));
  OAI211_X1 g459(.A(new_n616), .B(new_n620), .C1(new_n641), .C2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  AOI211_X1 g462(.A(KEYINPUT101), .B(new_n594), .C1(new_n608), .C2(new_n188), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n607), .A2(new_n609), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n649), .B1(new_n650), .B2(KEYINPUT101), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n651), .B(new_n593), .C1(new_n564), .C2(new_n565), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n507), .B1(new_n490), .B2(new_n491), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n502), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n620), .A2(new_n616), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(KEYINPUT35), .B(G107), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G9));
  NAND2_X1  g472(.A1(new_n239), .A2(new_n240), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n189), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT36), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n233), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n223), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n189), .A2(G902), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n213), .A2(new_n233), .A3(new_n661), .A4(new_n222), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n660), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n612), .A2(new_n351), .A3(new_n618), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT37), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(new_n423), .ZN(G12));
  OAI21_X1  g486(.A(new_n355), .B1(new_n362), .B2(new_n352), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n351), .A2(KEYINPUT74), .A3(new_n353), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n377), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(new_n494), .B(KEYINPUT103), .Z(new_n676));
  INV_X1    g490(.A(G900), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n676), .B1(new_n498), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n652), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n666), .B(KEYINPUT102), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n241), .ZN(new_n681));
  NOR3_X1   g495(.A1(new_n639), .A2(new_n681), .A3(new_n507), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n675), .A2(new_n616), .A3(new_n679), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G128), .ZN(G30));
  XNOR2_X1  g498(.A(new_n492), .B(KEYINPUT38), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n678), .B(KEYINPUT39), .Z(new_n686));
  NAND2_X1  g500(.A1(new_n616), .A2(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n685), .B1(KEYINPUT40), .B2(new_n687), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n689));
  NOR4_X1   g503(.A1(new_n688), .A2(new_n689), .A3(new_n507), .A4(new_n669), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n610), .B1(new_n564), .B2(new_n565), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n362), .A2(KEYINPUT32), .ZN(new_n693));
  INV_X1    g507(.A(G472), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n342), .A2(new_n336), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n328), .B1(new_n695), .B2(new_n339), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n694), .B1(new_n696), .B2(new_n188), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n673), .A2(new_n693), .A3(new_n674), .A4(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n690), .A2(new_n692), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G143), .ZN(G45));
  INV_X1    g515(.A(new_n678), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n632), .A2(new_n610), .A3(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n675), .A2(new_n616), .A3(new_n682), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  OR2_X1    g520(.A1(new_n438), .A2(new_n439), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n188), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(G469), .ZN(new_n709));
  INV_X1    g523(.A(new_n505), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n709), .A2(new_n440), .A3(new_n710), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n378), .B(new_n711), .C1(new_n641), .C2(new_n645), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT41), .B(G113), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G15));
  XNOR2_X1  g528(.A(new_n244), .B(KEYINPUT80), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n675), .A2(new_n715), .A3(new_n655), .A4(new_n711), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  AND4_X1   g531(.A1(new_n502), .A2(new_n711), .A3(new_n653), .A4(new_n669), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n675), .A3(new_n611), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G119), .ZN(G21));
  AND2_X1   g534(.A1(new_n371), .A2(new_n341), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n329), .B(new_n325), .C1(new_n339), .C2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n350), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT104), .B1(new_n617), .B2(G472), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT104), .ZN(new_n725));
  AOI211_X1 g539(.A(new_n725), .B(new_n694), .C1(new_n349), .C2(new_n188), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n244), .B(new_n723), .C1(new_n724), .C2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n709), .A2(new_n440), .A3(new_n710), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n653), .B(new_n610), .C1(new_n564), .C2(new_n565), .ZN(new_n729));
  NOR4_X1   g543(.A1(new_n727), .A2(new_n501), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n515), .ZN(G24));
  INV_X1    g545(.A(new_n724), .ZN(new_n732));
  INV_X1    g546(.A(new_n726), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n711), .A2(new_n653), .A3(new_n669), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n734), .A2(new_n735), .A3(new_n704), .A4(new_n723), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G125), .ZN(G27));
  INV_X1    g551(.A(KEYINPUT105), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n434), .A2(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n433), .A2(new_n412), .A3(new_n427), .A4(KEYINPUT105), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n431), .A2(new_n741), .A3(G469), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n505), .B1(new_n443), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n639), .A3(new_n506), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n703), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n376), .A2(G472), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT32), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n351), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n693), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n745), .A2(new_n749), .A3(new_n244), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT42), .ZN(new_n751));
  INV_X1    g565(.A(new_n744), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n703), .A2(KEYINPUT42), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n675), .A2(new_n715), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G131), .ZN(G33));
  NAND4_X1  g570(.A1(new_n378), .A2(KEYINPUT106), .A3(new_n679), .A4(new_n752), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n675), .A2(new_n715), .A3(new_n679), .A4(new_n752), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT106), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G134), .ZN(G36));
  NOR2_X1   g576(.A1(new_n435), .A2(KEYINPUT45), .ZN(new_n763));
  AND2_X1   g577(.A1(new_n431), .A2(new_n741), .ZN(new_n764));
  AOI211_X1 g578(.A(new_n437), .B(new_n763), .C1(KEYINPUT45), .C2(new_n764), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n765), .A2(new_n441), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT46), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n440), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n769), .B1(new_n766), .B2(new_n767), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n505), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  AND2_X1   g585(.A1(new_n771), .A2(new_n686), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n639), .A2(new_n506), .ZN(new_n773));
  INV_X1    g587(.A(new_n610), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n632), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g589(.A(new_n775), .B(KEYINPUT43), .Z(new_n776));
  AND3_X1   g590(.A1(new_n776), .A2(new_n619), .A3(new_n669), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n773), .B1(new_n777), .B2(KEYINPUT44), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n772), .B(new_n778), .C1(KEYINPUT44), .C2(new_n777), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G137), .ZN(G39));
  NAND2_X1  g594(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n781));
  OR2_X1    g595(.A1(new_n771), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n781), .B1(new_n771), .B2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n773), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n675), .A2(new_n715), .A3(new_n703), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n782), .A2(new_n784), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  AND2_X1   g602(.A1(new_n709), .A2(new_n440), .ZN(new_n789));
  XOR2_X1   g603(.A(new_n789), .B(KEYINPUT49), .Z(new_n790));
  NOR3_X1   g604(.A1(new_n790), .A2(new_n699), .A3(new_n775), .ZN(new_n791));
  INV_X1    g605(.A(new_n685), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n791), .A2(new_n244), .A3(new_n510), .A4(new_n792), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n776), .A2(new_n676), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n794), .A2(new_n785), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n795), .A2(new_n711), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n734), .A2(new_n723), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n796), .A2(new_n669), .A3(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n727), .A2(new_n728), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n794), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n507), .A3(new_n792), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT50), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n785), .A2(new_n494), .A3(new_n711), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n699), .A2(new_n803), .A3(new_n246), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n632), .A2(new_n610), .ZN(new_n805));
  AOI211_X1 g619(.A(new_n798), .B(new_n802), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT51), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n782), .A2(new_n784), .ZN(new_n809));
  XOR2_X1   g623(.A(new_n789), .B(KEYINPUT111), .Z(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n710), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n795), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n806), .B1(new_n727), .B2(new_n812), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n808), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n808), .A2(new_n813), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n804), .A2(new_n636), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n749), .A2(new_n244), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n796), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT48), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n819), .A2(KEYINPUT114), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT113), .Z(new_n821));
  XNOR2_X1  g635(.A(new_n818), .B(new_n821), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n819), .A2(KEYINPUT114), .ZN(new_n823));
  AOI211_X1 g637(.A(new_n493), .B(new_n816), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n814), .A2(new_n815), .A3(new_n824), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n800), .A2(new_n653), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n716), .A2(new_n719), .ZN(new_n827));
  INV_X1    g641(.A(new_n729), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n799), .A2(new_n502), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n561), .A2(new_n563), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n642), .B1(new_n831), .B2(new_n610), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n513), .A2(new_n832), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n833), .A2(new_n246), .A3(new_n619), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n827), .A2(new_n712), .A3(new_n829), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n613), .A2(new_n670), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT108), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n743), .A2(new_n839), .A3(new_n681), .A4(new_n702), .ZN(new_n840));
  INV_X1    g654(.A(new_n742), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n440), .A2(new_n442), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n710), .B(new_n702), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(KEYINPUT108), .B1(new_n843), .B2(new_n669), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n699), .A3(new_n828), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n683), .A2(new_n705), .A3(new_n846), .A4(new_n736), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT52), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n616), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n850), .B1(new_n357), .B2(new_n377), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n851), .B(new_n682), .C1(new_n679), .C2(new_n704), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(KEYINPUT52), .A3(new_n736), .A4(new_n846), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n797), .A2(new_n669), .A3(new_n745), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n761), .A2(new_n755), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n593), .ZN(new_n857));
  NOR4_X1   g671(.A1(new_n681), .A2(new_n830), .A3(new_n857), .A4(new_n678), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n851), .A2(new_n651), .A3(new_n785), .A4(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n838), .A2(new_n854), .A3(new_n856), .A4(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(KEYINPUT110), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT109), .B1(new_n847), .B2(new_n848), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n847), .A2(new_n848), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n847), .A2(KEYINPUT109), .A3(new_n848), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n675), .A2(new_n715), .A3(new_n711), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n636), .A2(new_n640), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT100), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n636), .A2(KEYINPUT100), .A3(new_n640), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n716), .A2(new_n719), .ZN(new_n875));
  NOR4_X1   g689(.A1(new_n874), .A2(new_n875), .A3(new_n730), .A4(new_n834), .ZN(new_n876));
  INV_X1    g690(.A(new_n837), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n856), .A2(new_n876), .A3(new_n877), .A4(new_n859), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n868), .A2(new_n878), .A3(new_n861), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT110), .B1(new_n860), .B2(new_n861), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n863), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n868), .ZN(new_n884));
  INV_X1    g698(.A(new_n878), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n884), .A2(new_n885), .A3(new_n861), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n860), .A2(KEYINPUT53), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n883), .B1(new_n882), .B2(new_n888), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n825), .A2(new_n826), .A3(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(G952), .A2(G953), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n793), .B1(new_n890), .B2(new_n891), .ZN(G75));
  NOR2_X1   g706(.A1(new_n881), .A2(new_n188), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(G210), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n460), .B(new_n466), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT55), .ZN(new_n896));
  NOR2_X1   g710(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n897));
  AND2_X1   g711(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n894), .B(new_n896), .C1(new_n897), .C2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n228), .A2(G952), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT56), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n896), .B1(new_n894), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n903), .A2(KEYINPUT115), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT115), .ZN(new_n905));
  AOI211_X1 g719(.A(new_n905), .B(new_n896), .C1(new_n894), .C2(new_n902), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n899), .B(new_n901), .C1(new_n904), .C2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(G51));
  INV_X1    g722(.A(new_n707), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT118), .B1(new_n881), .B2(new_n882), .ZN(new_n910));
  INV_X1    g724(.A(new_n880), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT53), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n911), .A2(new_n912), .A3(new_n862), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT54), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n910), .A2(new_n883), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g730(.A(KEYINPUT117), .B(KEYINPUT57), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(new_n441), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n909), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n893), .A2(new_n765), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n901), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT119), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  OAI211_X1 g737(.A(KEYINPUT119), .B(new_n901), .C1(new_n919), .C2(new_n920), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(G54));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT58), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n926), .B1(new_n927), .B2(new_n606), .ZN(new_n928));
  NAND3_X1  g742(.A1(KEYINPUT120), .A2(KEYINPUT58), .A3(G475), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n893), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(new_n605), .Z(new_n931));
  NOR2_X1   g745(.A1(new_n931), .A2(new_n900), .ZN(G60));
  NAND2_X1  g746(.A1(new_n626), .A2(new_n628), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT121), .Z(new_n934));
  NAND2_X1  g748(.A1(G478), .A2(G902), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT59), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n934), .B1(new_n889), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n916), .A2(new_n936), .A3(new_n934), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(KEYINPUT122), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n916), .A2(new_n940), .A3(new_n936), .A4(new_n934), .ZN(new_n941));
  AOI211_X1 g755(.A(new_n900), .B(new_n937), .C1(new_n939), .C2(new_n941), .ZN(G63));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT60), .Z(new_n944));
  NAND2_X1  g758(.A1(new_n913), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n900), .B1(new_n945), .B2(new_n242), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n663), .A2(new_n665), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(new_n945), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n948), .B(KEYINPUT61), .Z(G66));
  INV_X1    g763(.A(new_n838), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n224), .B1(new_n499), .B2(G224), .ZN(new_n952));
  AOI22_X1  g766(.A1(new_n950), .A2(new_n228), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n951), .B2(new_n952), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n460), .B1(G898), .B2(new_n228), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n954), .B(new_n955), .ZN(G69));
  AND2_X1   g770(.A1(new_n779), .A2(new_n787), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n378), .A2(new_n832), .ZN(new_n958));
  OR3_X1    g772(.A1(new_n958), .A2(new_n687), .A3(new_n773), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n852), .A2(new_n736), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n700), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT62), .Z(new_n962));
  NAND3_X1  g776(.A1(new_n957), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n228), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n319), .A2(new_n320), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(new_n598), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n495), .A2(new_n677), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n772), .A2(new_n828), .A3(new_n817), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n761), .A2(new_n755), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT124), .Z(new_n971));
  NAND4_X1  g785(.A1(new_n957), .A2(new_n960), .A3(new_n969), .A4(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n966), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n972), .A2(new_n228), .A3(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n967), .A2(new_n968), .A3(new_n974), .ZN(new_n975));
  OR2_X1    g789(.A1(new_n975), .A2(KEYINPUT126), .ZN(new_n976));
  AND2_X1   g790(.A1(G227), .A2(G900), .ZN(new_n977));
  AOI211_X1 g791(.A(new_n228), .B(new_n977), .C1(new_n973), .C2(KEYINPUT125), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n975), .A2(KEYINPUT126), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n978), .B1(new_n976), .B2(new_n979), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n980), .A2(new_n981), .ZN(G72));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT63), .Z(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n963), .B2(new_n950), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n985), .A2(new_n305), .A3(new_n365), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT127), .Z(new_n987));
  OR2_X1    g801(.A1(new_n972), .A2(new_n950), .ZN(new_n988));
  AOI211_X1 g802(.A(new_n305), .B(new_n365), .C1(new_n988), .C2(new_n984), .ZN(new_n989));
  INV_X1    g803(.A(new_n984), .ZN(new_n990));
  AOI211_X1 g804(.A(new_n990), .B(new_n888), .C1(new_n328), .C2(new_n367), .ZN(new_n991));
  NOR4_X1   g805(.A1(new_n987), .A2(new_n900), .A3(new_n989), .A4(new_n991), .ZN(G57));
endmodule


