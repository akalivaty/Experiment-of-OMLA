//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 1 1 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(new_n192), .A3(KEYINPUT77), .ZN(new_n193));
  OR3_X1    g007(.A1(new_n191), .A2(KEYINPUT77), .A3(G140), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n188), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n190), .A2(KEYINPUT16), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n187), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n196), .ZN(new_n198));
  NOR3_X1   g012(.A1(new_n191), .A2(KEYINPUT77), .A3(G140), .ZN(new_n199));
  XNOR2_X1  g013(.A(G125), .B(G140), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(KEYINPUT77), .ZN(new_n201));
  OAI211_X1 g015(.A(G146), .B(new_n198), .C1(new_n201), .C2(new_n188), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(G119), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT68), .B(G128), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G119), .ZN(new_n206));
  XOR2_X1   g020(.A(KEYINPUT24), .B(G110), .Z(new_n207));
  AOI22_X1  g021(.A1(new_n197), .A2(new_n202), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G119), .ZN(new_n209));
  NOR3_X1   g023(.A1(new_n209), .A2(KEYINPUT23), .A3(G128), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n210), .B1(new_n206), .B2(KEYINPUT23), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G110), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n200), .A2(new_n187), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n211), .A2(G110), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n206), .A2(new_n207), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n202), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n213), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G953), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(G221), .A3(G234), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n220), .B(KEYINPUT22), .ZN(new_n221));
  XNOR2_X1  g035(.A(new_n221), .B(G137), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n213), .A2(new_n217), .A3(new_n222), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G217), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT75), .B(G902), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n228), .B1(new_n230), .B2(G234), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(G902), .ZN(new_n232));
  XNOR2_X1  g046(.A(new_n232), .B(KEYINPUT78), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n227), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n226), .A2(new_n230), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT25), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n235), .B(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n234), .B1(new_n237), .B2(new_n231), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G137), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(KEYINPUT11), .A3(G134), .ZN(new_n241));
  INV_X1    g055(.A(G134), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G137), .ZN(new_n243));
  AND2_X1   g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G131), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT67), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT67), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G131), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT11), .ZN(new_n250));
  OAI211_X1 g064(.A(KEYINPUT66), .B(new_n250), .C1(new_n242), .C2(G137), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n240), .A2(G134), .ZN(new_n253));
  AOI21_X1  g067(.A(KEYINPUT66), .B1(new_n253), .B2(new_n250), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n244), .B(new_n249), .C1(new_n252), .C2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n243), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G131), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(G143), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G146), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n187), .A2(G143), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n262), .A2(new_n263), .A3(new_n264), .A4(G128), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT65), .B1(new_n187), .B2(G143), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT65), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(new_n261), .A3(G146), .ZN(new_n268));
  OAI21_X1  g082(.A(KEYINPUT64), .B1(new_n261), .B2(G146), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT64), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(new_n187), .A3(G143), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n266), .A2(new_n268), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n264), .B1(G143), .B2(new_n187), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n205), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n265), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n255), .A2(KEYINPUT70), .A3(new_n257), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n260), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(KEYINPUT69), .B1(new_n209), .B2(G116), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n279));
  INV_X1    g093(.A(G116), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(new_n280), .A3(G119), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n282), .B1(new_n280), .B2(G119), .ZN(new_n283));
  XOR2_X1   g097(.A(KEYINPUT2), .B(G113), .Z(new_n284));
  XNOR2_X1  g098(.A(new_n283), .B(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n241), .A2(new_n243), .ZN(new_n286));
  INV_X1    g100(.A(new_n254), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n286), .B1(new_n287), .B2(new_n251), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n255), .B1(new_n288), .B2(new_n245), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n262), .A2(new_n263), .A3(G128), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT0), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  XOR2_X1   g106(.A(KEYINPUT0), .B(G128), .Z(new_n293));
  NAND2_X1  g107(.A1(new_n266), .A2(new_n268), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n269), .A2(new_n271), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n292), .B1(new_n293), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n289), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n277), .A2(new_n285), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT28), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(G237), .A2(G953), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G210), .ZN(new_n303));
  XOR2_X1   g117(.A(new_n303), .B(KEYINPUT27), .Z(new_n304));
  XNOR2_X1  g118(.A(new_n304), .B(KEYINPUT26), .ZN(new_n305));
  INV_X1    g119(.A(G101), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n305), .B(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n275), .A2(new_n255), .A3(new_n257), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n285), .B1(new_n298), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n299), .A2(KEYINPUT71), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n277), .A2(new_n311), .A3(new_n285), .A4(new_n298), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n309), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n301), .B(new_n307), .C1(new_n313), .C2(new_n300), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT72), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n310), .A2(new_n312), .ZN(new_n317));
  INV_X1    g131(.A(new_n285), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT30), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n319), .B1(new_n277), .B2(new_n298), .ZN(new_n320));
  AND3_X1   g134(.A1(new_n298), .A2(new_n319), .A3(new_n308), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n318), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n305), .B(G101), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT73), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n323), .A2(KEYINPUT73), .A3(new_n324), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n316), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT29), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n330), .B1(new_n314), .B2(new_n315), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n324), .A2(new_n330), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n277), .A2(new_n298), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n310), .A2(new_n312), .B1(new_n318), .B2(new_n334), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n301), .B(new_n333), .C1(new_n335), .C2(new_n300), .ZN(new_n336));
  AND2_X1   g150(.A1(new_n336), .A2(KEYINPUT74), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n336), .A2(KEYINPUT74), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n230), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(G472), .B1(new_n332), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT73), .B1(new_n323), .B2(new_n324), .ZN(new_n343));
  AOI211_X1 g157(.A(new_n326), .B(new_n307), .C1(new_n317), .C2(new_n322), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n310), .A2(new_n312), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT28), .B1(new_n346), .B2(new_n309), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n347), .A2(KEYINPUT72), .A3(new_n301), .A4(new_n307), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n345), .A2(new_n348), .A3(new_n330), .A4(new_n316), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n285), .B1(new_n277), .B2(new_n298), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT28), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT74), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n351), .A2(new_n352), .A3(new_n301), .A4(new_n333), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n336), .A2(KEYINPUT74), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n229), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n349), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(KEYINPUT76), .A3(G472), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n342), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G472), .ZN(new_n359));
  INV_X1    g173(.A(G902), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n317), .A2(new_n322), .A3(new_n307), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT31), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n317), .A2(new_n322), .A3(KEYINPUT31), .A4(new_n307), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n301), .B1(new_n313), .B2(new_n300), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n324), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n361), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT32), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n369), .A2(KEYINPUT32), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n239), .B1(new_n358), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G221), .ZN(new_n375));
  XOR2_X1   g189(.A(KEYINPUT9), .B(G234), .Z(new_n376));
  AOI21_X1  g190(.A(new_n375), .B1(new_n376), .B2(new_n360), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT80), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT3), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G104), .ZN(new_n380));
  NOR2_X1   g194(.A1(KEYINPUT79), .A2(G107), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(KEYINPUT79), .A2(G107), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n380), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G104), .ZN(new_n385));
  AOI21_X1  g199(.A(G107), .B1(new_n385), .B2(KEYINPUT3), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n385), .A2(KEYINPUT3), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n378), .B1(new_n384), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n383), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n387), .B1(new_n390), .B2(new_n381), .ZN(new_n391));
  INV_X1    g205(.A(G107), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n379), .B2(G104), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n380), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(new_n394), .A3(KEYINPUT80), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n389), .A2(new_n395), .A3(G101), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n391), .A2(new_n394), .A3(new_n306), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n397), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n297), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n265), .ZN(new_n402));
  OR2_X1    g216(.A1(new_n205), .A2(new_n273), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n402), .B1(new_n403), .B2(new_n296), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n385), .B1(new_n390), .B2(new_n381), .ZN(new_n405));
  NAND2_X1  g219(.A1(G104), .A2(G107), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(G101), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n399), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT10), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n404), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n203), .B1(new_n263), .B2(KEYINPUT1), .ZN(new_n411));
  XNOR2_X1  g225(.A(G143), .B(G146), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n265), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(new_n399), .A3(new_n407), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT82), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT82), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n414), .A2(new_n418), .A3(new_n415), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n410), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n289), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n401), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT83), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n401), .A2(new_n420), .A3(KEYINPUT83), .A4(new_n421), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n399), .A2(new_n407), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT84), .B1(new_n427), .B2(new_n275), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT84), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n404), .A2(new_n429), .A3(new_n408), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(new_n414), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n289), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT12), .ZN(new_n433));
  OAI21_X1  g247(.A(KEYINPUT85), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n433), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT85), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n431), .A2(new_n436), .A3(KEYINPUT12), .A4(new_n289), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n426), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G140), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n219), .A2(G227), .ZN(new_n441));
  XOR2_X1   g255(.A(new_n440), .B(new_n441), .Z(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(new_n424), .B2(new_n425), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n401), .A2(new_n420), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n289), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n439), .A2(new_n443), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(G469), .B1(new_n447), .B2(G902), .ZN(new_n448));
  INV_X1    g262(.A(G469), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n426), .A2(new_n438), .A3(new_n442), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n442), .B1(new_n426), .B2(new_n446), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n449), .B(new_n230), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  AOI211_X1 g266(.A(KEYINPUT86), .B(new_n377), .C1(new_n448), .C2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT86), .ZN(new_n454));
  NAND2_X1  g268(.A1(G469), .A2(G902), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n439), .A2(new_n443), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n444), .A2(new_n446), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(G469), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n452), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n377), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n454), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OR2_X1    g275(.A1(new_n453), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G475), .ZN(new_n463));
  INV_X1    g277(.A(G237), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(new_n219), .A3(G214), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n261), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n302), .A2(G143), .A3(G214), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n249), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(KEYINPUT17), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n197), .A2(new_n202), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT95), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n466), .A2(new_n249), .A3(new_n467), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT93), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n468), .A2(new_n469), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT17), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT93), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n466), .A2(new_n249), .A3(new_n477), .A4(new_n467), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n474), .A2(new_n475), .A3(new_n476), .A4(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT95), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n197), .A2(new_n202), .A3(new_n480), .A4(new_n470), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n472), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(KEYINPUT18), .A2(G131), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n468), .B(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n193), .A2(new_n194), .A3(G146), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT92), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n485), .A2(new_n486), .A3(new_n214), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n486), .B1(new_n485), .B2(new_n214), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n484), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n482), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(G113), .B(G122), .ZN(new_n491));
  XNOR2_X1  g305(.A(new_n491), .B(new_n385), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n482), .A2(new_n492), .A3(new_n489), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n463), .B1(new_n496), .B2(new_n360), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT94), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n474), .A2(new_n475), .A3(new_n478), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT19), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n200), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n193), .A2(new_n194), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n187), .B(new_n501), .C1(new_n502), .C2(new_n500), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n499), .A2(new_n202), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n489), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n498), .B1(new_n505), .B2(new_n493), .ZN(new_n506));
  AOI211_X1 g320(.A(KEYINPUT94), .B(new_n492), .C1(new_n489), .C2(new_n504), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n495), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT20), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n463), .A2(new_n360), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(KEYINPUT96), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n509), .B1(new_n508), .B2(new_n511), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT97), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND4_X1  g329(.A1(new_n508), .A2(KEYINPUT97), .A3(new_n509), .A4(new_n511), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n497), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT98), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n517), .B(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n297), .A2(new_n191), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(KEYINPUT88), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n404), .A2(new_n191), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(G224), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n524), .A2(G953), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n525), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n521), .A2(new_n522), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n318), .B1(new_n398), .B2(new_n400), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT5), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(new_n209), .A3(G116), .ZN(new_n532));
  OAI211_X1 g346(.A(G113), .B(new_n532), .C1(new_n283), .C2(new_n531), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n284), .B(new_n282), .C1(new_n280), .C2(G119), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n427), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g350(.A(G110), .B(G122), .Z(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n537), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n530), .A2(new_n535), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(KEYINPUT6), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n539), .B1(new_n530), .B2(new_n535), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT87), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT6), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n543), .B1(new_n542), .B2(new_n544), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n529), .B(new_n541), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(new_n521), .B2(KEYINPUT89), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(new_n523), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n521), .B(new_n522), .C1(KEYINPUT89), .C2(new_n548), .ZN(new_n551));
  XOR2_X1   g365(.A(new_n537), .B(KEYINPUT8), .Z(new_n552));
  INV_X1    g366(.A(new_n535), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n427), .B1(new_n533), .B2(new_n534), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n550), .A2(new_n551), .A3(new_n540), .A4(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n547), .A2(new_n360), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(G210), .B1(G237), .B2(G902), .ZN(new_n558));
  XOR2_X1   g372(.A(new_n558), .B(KEYINPUT90), .Z(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT91), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n559), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n547), .A2(new_n360), .A3(new_n562), .A4(new_n556), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(G214), .B1(G237), .B2(G902), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G122), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G116), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(G116), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT14), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  XOR2_X1   g385(.A(new_n571), .B(KEYINPUT100), .Z(new_n572));
  INV_X1    g386(.A(new_n569), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(KEYINPUT14), .ZN(new_n574));
  OAI21_X1  g388(.A(G107), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n573), .A2(new_n568), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n382), .A2(new_n383), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n205), .A2(G143), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n203), .B2(G143), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(G134), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n575), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n576), .B(new_n577), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n203), .A2(G143), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT99), .ZN(new_n585));
  OR3_X1    g399(.A1(new_n584), .A2(new_n585), .A3(KEYINPUT13), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n585), .B1(new_n584), .B2(KEYINPUT13), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n584), .A2(KEYINPUT13), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n586), .A2(new_n587), .A3(new_n588), .A4(new_n579), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G134), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n583), .B(new_n590), .C1(G134), .C2(new_n580), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n582), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n376), .A2(G217), .A3(new_n219), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n592), .A2(new_n593), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n230), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(G478), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(KEYINPUT15), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n596), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(G234), .A2(G237), .ZN(new_n600));
  AND3_X1   g414(.A1(new_n600), .A2(G952), .A3(new_n219), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n229), .A2(G953), .A3(new_n600), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  XOR2_X1   g418(.A(KEYINPUT21), .B(G898), .Z(new_n605));
  OAI21_X1  g419(.A(new_n602), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NOR4_X1   g421(.A1(new_n519), .A2(new_n566), .A3(new_n599), .A4(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n374), .A2(new_n462), .A3(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G101), .ZN(G3));
  AOI22_X1  g424(.A1(new_n364), .A2(new_n365), .B1(new_n367), .B2(new_n324), .ZN(new_n611));
  OAI21_X1  g425(.A(G472), .B1(new_n611), .B2(new_n229), .ZN(new_n612));
  INV_X1    g426(.A(new_n369), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n239), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n615), .B1(new_n453), .B2(new_n461), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT101), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI211_X1 g432(.A(new_n615), .B(KEYINPUT101), .C1(new_n453), .C2(new_n461), .ZN(new_n619));
  INV_X1    g433(.A(new_n565), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n557), .A2(new_n559), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n620), .B1(new_n621), .B2(new_n563), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n515), .A2(new_n516), .ZN(new_n624));
  INV_X1    g438(.A(new_n497), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n518), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI211_X1 g440(.A(KEYINPUT98), .B(new_n497), .C1(new_n515), .C2(new_n516), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OR2_X1    g442(.A1(new_n596), .A2(G478), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n594), .A2(new_n595), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n632), .B1(new_n592), .B2(new_n633), .ZN(new_n634));
  OR2_X1    g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n631), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(new_n230), .A3(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n630), .B1(new_n637), .B2(G478), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NOR4_X1   g453(.A1(new_n623), .A2(new_n628), .A3(new_n607), .A4(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n618), .A2(new_n619), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  NAND2_X1  g457(.A1(new_n508), .A2(new_n511), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(KEYINPUT20), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(KEYINPUT103), .A3(new_n512), .ZN(new_n646));
  OR3_X1    g460(.A1(new_n644), .A2(KEYINPUT103), .A3(KEYINPUT20), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n646), .A2(new_n647), .A3(new_n625), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n599), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n623), .A2(new_n607), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n618), .A2(new_n619), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  INV_X1    g467(.A(new_n614), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n237), .A2(new_n231), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n223), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n218), .B(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n658), .A2(new_n233), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n655), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n608), .A2(new_n462), .A3(new_n654), .A4(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n661), .B(KEYINPUT37), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G110), .ZN(G12));
  INV_X1    g477(.A(new_n660), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n664), .B1(new_n358), .B2(new_n373), .ZN(new_n665));
  INV_X1    g479(.A(G900), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n601), .B1(new_n603), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n649), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n665), .A2(new_n462), .A3(new_n622), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  XNOR2_X1  g484(.A(new_n667), .B(KEYINPUT39), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n462), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT40), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n519), .A2(new_n565), .A3(new_n664), .A4(new_n599), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n677));
  OR2_X1    g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT104), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n564), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT38), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT32), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n613), .A2(new_n682), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n362), .B1(new_n307), .B2(new_n335), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n360), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(G472), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n683), .A2(new_n370), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n676), .B2(new_n677), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n675), .A2(new_n678), .A3(new_n681), .A4(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G143), .ZN(G45));
  INV_X1    g505(.A(new_n667), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n638), .B(new_n692), .C1(new_n626), .C2(new_n627), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n665), .A2(new_n695), .A3(new_n462), .A4(new_n622), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G146), .ZN(G48));
  AOI21_X1  g511(.A(KEYINPUT76), .B1(new_n356), .B2(G472), .ZN(new_n698));
  AOI211_X1 g512(.A(new_n341), .B(new_n359), .C1(new_n349), .C2(new_n355), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n373), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n230), .B1(new_n450), .B2(new_n451), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(G469), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(new_n460), .A3(new_n452), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n640), .A2(new_n700), .A3(new_n238), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT41), .B(G113), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G15));
  NAND4_X1  g521(.A1(new_n700), .A2(new_n650), .A3(new_n238), .A4(new_n704), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G116), .ZN(G18));
  NOR3_X1   g523(.A1(new_n519), .A2(new_n599), .A3(new_n607), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n623), .A2(new_n703), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n700), .A2(new_n710), .A3(new_n660), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  INV_X1    g527(.A(new_n366), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n307), .B1(new_n351), .B2(new_n301), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n359), .B(new_n360), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n612), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n238), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n703), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n599), .B1(new_n626), .B2(new_n627), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI211_X1 g537(.A(KEYINPUT107), .B(new_n599), .C1(new_n626), .C2(new_n627), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n720), .A2(new_n725), .A3(new_n606), .A4(new_n622), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  NAND4_X1  g541(.A1(new_n519), .A2(new_n694), .A3(new_n638), .A4(new_n692), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n693), .A2(KEYINPUT106), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n664), .A2(new_n717), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n728), .A2(new_n729), .A3(new_n711), .A4(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n731), .B(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  AND3_X1   g548(.A1(new_n561), .A2(new_n563), .A3(new_n565), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n377), .B1(new_n448), .B2(new_n452), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n738), .B1(new_n369), .B2(KEYINPUT32), .ZN(new_n739));
  NOR4_X1   g553(.A1(new_n611), .A2(KEYINPUT109), .A3(new_n682), .A4(new_n361), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n739), .A2(new_n740), .A3(new_n372), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n741), .B1(new_n698), .B2(new_n699), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n695), .A2(new_n238), .A3(new_n737), .A4(new_n742), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n700), .A2(new_n238), .A3(new_n737), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n728), .A2(new_n729), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(KEYINPUT42), .ZN(new_n746));
  AOI22_X1  g560(.A1(new_n743), .A2(KEYINPUT42), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G131), .ZN(G33));
  NAND2_X1  g562(.A1(new_n744), .A2(new_n668), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G134), .ZN(G36));
  NOR2_X1   g564(.A1(new_n519), .A2(new_n639), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT43), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n753), .B1(new_n519), .B2(new_n639), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n614), .A2(new_n660), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(KEYINPUT110), .Z(new_n757));
  NAND2_X1  g571(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OR2_X1    g574(.A1(new_n447), .A2(KEYINPUT45), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n447), .A2(KEYINPUT45), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n761), .A2(G469), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n455), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT46), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n763), .A2(KEYINPUT46), .A3(new_n455), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(new_n452), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n460), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(new_n671), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n760), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n735), .B1(new_n758), .B2(new_n759), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G137), .ZN(G39));
  NAND2_X1  g588(.A1(new_n769), .A2(KEYINPUT47), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n358), .A2(new_n239), .A3(new_n373), .A4(new_n735), .ZN(new_n776));
  INV_X1    g590(.A(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT47), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n768), .A2(new_n778), .A3(new_n460), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n775), .A2(new_n695), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G140), .ZN(G42));
  OR2_X1    g595(.A1(G952), .A2(G953), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n566), .A2(new_n607), .ZN(new_n783));
  INV_X1    g597(.A(new_n599), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n519), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n618), .A2(new_n619), .A3(new_n783), .A4(new_n785), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n786), .A2(KEYINPUT112), .A3(new_n661), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT112), .B1(new_n786), .B2(new_n661), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n628), .A2(new_n639), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n618), .A2(new_n619), .A3(new_n789), .A4(new_n783), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n609), .A2(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n787), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n742), .A2(new_n238), .A3(new_n737), .ZN(new_n793));
  OAI21_X1  g607(.A(KEYINPUT42), .B1(new_n793), .B2(new_n745), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT42), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n374), .A2(new_n695), .A3(new_n795), .A4(new_n737), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n728), .A2(new_n729), .A3(new_n730), .A4(new_n737), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n797), .A2(KEYINPUT115), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n797), .A2(KEYINPUT115), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n794), .B(new_n796), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n648), .A2(new_n561), .A3(new_n563), .A4(new_n565), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n599), .A2(new_n667), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(KEYINPUT113), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT113), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n735), .A2(new_n806), .A3(new_n648), .A4(new_n803), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n665), .A2(new_n801), .A3(new_n462), .A4(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n808), .A2(new_n462), .A3(new_n700), .A4(new_n660), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT114), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n749), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n800), .A2(new_n812), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n712), .A2(new_n708), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n814), .A2(KEYINPUT111), .A3(new_n705), .A4(new_n726), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n705), .A2(new_n726), .A3(new_n712), .A4(new_n708), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT111), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n792), .A2(new_n813), .A3(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n731), .A2(new_n732), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n731), .A2(new_n732), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n669), .B(new_n696), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n687), .A2(new_n736), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n660), .A2(new_n667), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n725), .A2(new_n824), .A3(new_n622), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT116), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n623), .B1(new_n723), .B2(new_n724), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n828), .A2(new_n829), .A3(new_n825), .A4(new_n824), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT52), .B1(new_n823), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n827), .A2(new_n830), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT52), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n700), .A2(new_n462), .A3(new_n622), .A4(new_n660), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(new_n668), .B2(new_n695), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n833), .A2(new_n834), .A3(new_n733), .A4(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n820), .A2(new_n838), .A3(KEYINPUT53), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n792), .A2(new_n813), .A3(new_n819), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n832), .A2(new_n837), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n839), .A2(KEYINPUT117), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n845), .B(new_n840), .C1(new_n841), .C2(new_n842), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n844), .A2(KEYINPUT54), .A3(new_n846), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n809), .A2(new_n811), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n797), .B(KEYINPUT115), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n747), .A3(new_n749), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n786), .A2(new_n661), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT112), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n609), .A2(new_n790), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n786), .A2(KEYINPUT112), .A3(new_n661), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n850), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n816), .A2(new_n840), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n837), .A3(new_n832), .A4(new_n858), .ZN(new_n859));
  XOR2_X1   g673(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n860));
  AND3_X1   g674(.A1(new_n843), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n847), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n681), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n602), .B1(new_n752), .B2(new_n754), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n864), .A2(new_n620), .A3(new_n720), .A4(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n868), .A2(KEYINPUT50), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(KEYINPUT50), .ZN(new_n870));
  OR2_X1    g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n775), .A2(new_n779), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n702), .A2(new_n452), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n872), .B1(new_n460), .B2(new_n873), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n865), .A2(new_n735), .ZN(new_n875));
  INV_X1    g689(.A(new_n719), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n687), .A2(new_n602), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n878), .A2(new_n238), .A3(new_n704), .A4(new_n735), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT120), .Z(new_n880));
  NOR2_X1   g694(.A1(new_n519), .A2(new_n638), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n875), .A2(new_n704), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n884), .A2(new_n664), .A3(new_n717), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n871), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT51), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n871), .A2(new_n883), .A3(KEYINPUT51), .A4(new_n886), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n880), .A2(new_n789), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n865), .A2(new_n622), .A3(new_n720), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(G952), .A3(new_n219), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n742), .A2(new_n238), .ZN(new_n894));
  OR3_X1    g708(.A1(new_n884), .A2(KEYINPUT48), .A3(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT48), .B1(new_n884), .B2(new_n894), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n893), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n889), .A2(new_n890), .A3(new_n891), .A4(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n782), .B1(new_n863), .B2(new_n898), .ZN(new_n899));
  NOR4_X1   g713(.A1(new_n681), .A2(new_n239), .A3(new_n377), .A4(new_n620), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n873), .B(KEYINPUT49), .Z(new_n901));
  NAND4_X1  g715(.A1(new_n900), .A2(new_n688), .A3(new_n751), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n899), .A2(new_n902), .ZN(G75));
  OAI21_X1  g717(.A(new_n541), .B1(new_n545), .B2(new_n546), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(new_n529), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT55), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT56), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n843), .A2(new_n859), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(new_n230), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n908), .B1(new_n910), .B2(new_n560), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n843), .A2(new_n859), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n912), .A2(new_n229), .A3(new_n559), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n906), .B1(new_n913), .B2(new_n907), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n219), .A2(G952), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n911), .A2(new_n914), .A3(new_n915), .ZN(G51));
  XOR2_X1   g730(.A(new_n455), .B(KEYINPUT57), .Z(new_n917));
  AOI21_X1  g731(.A(new_n860), .B1(new_n843), .B2(new_n859), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n917), .B1(new_n861), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n451), .B2(new_n450), .ZN(new_n920));
  OR3_X1    g734(.A1(new_n909), .A2(new_n230), .A3(new_n763), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n915), .B1(new_n920), .B2(new_n921), .ZN(G54));
  NAND4_X1  g736(.A1(new_n912), .A2(KEYINPUT58), .A3(G475), .A4(new_n229), .ZN(new_n923));
  INV_X1    g737(.A(new_n508), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n923), .A2(new_n924), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n925), .A2(new_n926), .A3(new_n915), .ZN(G60));
  NAND2_X1  g741(.A1(new_n635), .A2(new_n636), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(G478), .A2(G902), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT59), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n929), .B(new_n931), .C1(new_n861), .C2(new_n918), .ZN(new_n932));
  INV_X1    g746(.A(new_n915), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n863), .A2(new_n931), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n934), .B1(new_n935), .B2(new_n928), .ZN(G63));
  XNOR2_X1  g750(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n228), .A2(new_n360), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n227), .B1(new_n909), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g755(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n940), .B1(new_n843), .B2(new_n859), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n657), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n941), .A2(new_n933), .A3(new_n942), .A4(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n942), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n933), .B1(new_n943), .B2(new_n226), .ZN(new_n947));
  AOI211_X1 g761(.A(new_n658), .B(new_n940), .C1(new_n843), .C2(new_n859), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n945), .A2(new_n949), .ZN(G66));
  AOI21_X1  g764(.A(new_n219), .B1(new_n605), .B2(G224), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n792), .A2(new_n819), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n951), .B1(new_n952), .B2(new_n219), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n904), .B1(G898), .B2(new_n219), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n953), .B(new_n954), .Z(G69));
  AOI21_X1  g769(.A(new_n219), .B1(G227), .B2(G900), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT125), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n320), .A2(new_n321), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n501), .B1(new_n502), .B2(new_n500), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(G900), .A2(G953), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n770), .A2(new_n238), .A3(new_n742), .A4(new_n828), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT126), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n823), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n780), .B(new_n749), .C1(new_n771), .C2(new_n772), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n964), .A2(new_n747), .A3(new_n965), .A4(new_n967), .ZN(new_n968));
  OAI211_X1 g782(.A(new_n960), .B(new_n961), .C1(new_n968), .C2(G953), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT124), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n957), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n785), .A2(new_n789), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT123), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n374), .A2(new_n735), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n973), .A2(new_n673), .A3(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n965), .A2(new_n690), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT62), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n965), .A2(new_n690), .A3(KEYINPUT62), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n975), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n773), .A2(new_n780), .ZN(new_n981));
  AOI21_X1  g795(.A(G953), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n969), .B1(new_n982), .B2(new_n960), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n971), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n971), .A2(new_n983), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(G72));
  NAND4_X1  g800(.A1(new_n980), .A2(new_n819), .A3(new_n792), .A4(new_n981), .ZN(new_n987));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT63), .Z(new_n989));
  AOI21_X1  g803(.A(new_n324), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n323), .B(KEYINPUT127), .Z(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n915), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n989), .B1(new_n968), .B2(new_n952), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n994), .A2(new_n324), .A3(new_n991), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n345), .A2(new_n362), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n844), .A2(new_n846), .A3(new_n989), .A4(new_n996), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n993), .A2(new_n995), .A3(new_n997), .ZN(G57));
endmodule


