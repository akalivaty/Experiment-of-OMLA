//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 0 1 1 0 1 0 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n566, new_n567, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  AND2_X1   g032(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n458));
  NOR2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(G125), .ZN(new_n461));
  INV_X1    g036(.A(G113), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  OAI22_X1  g038(.A1(new_n460), .A2(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(G2105), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n464), .A2(G2105), .B1(G101), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n468), .B1(new_n458), .B2(new_n459), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OR2_X1    g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(KEYINPUT66), .A3(new_n468), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n466), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  INV_X1    g053(.A(G2105), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n479), .B1(new_n472), .B2(new_n473), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  XOR2_X1   g056(.A(new_n481), .B(KEYINPUT68), .Z(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n479), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g060(.A(KEYINPUT67), .B1(new_n460), .B2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT67), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n474), .A2(new_n487), .A3(new_n479), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n485), .B1(G136), .B2(new_n490), .ZN(G162));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n493), .B(new_n495), .C1(new_n459), .C2(new_n458), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n479), .A2(G138), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n497), .B1(new_n472), .B2(new_n473), .ZN(new_n498));
  XNOR2_X1  g073(.A(KEYINPUT71), .B(KEYINPUT4), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n496), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g075(.A(G126), .B(G2105), .C1(new_n458), .C2(new_n459), .ZN(new_n501));
  OR2_X1    g076(.A1(KEYINPUT69), .A2(G114), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT69), .A2(G114), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n479), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n501), .B(KEYINPUT70), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT69), .A2(G114), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT69), .A2(G114), .ZN(new_n509));
  OAI21_X1  g084(.A(G2105), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n505), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(KEYINPUT70), .B1(new_n512), .B2(new_n501), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n500), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(G164));
  NAND2_X1  g090(.A1(G75), .A2(G543), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(G62), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n516), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n520), .A2(new_n521), .ZN(new_n525));
  OR2_X1    g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND2_X1   g103(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n524), .A2(G651), .B1(new_n529), .B2(G88), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n519), .B1(new_n526), .B2(new_n527), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G50), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT72), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n530), .A2(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n525), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n520), .A2(KEYINPUT74), .A3(new_n521), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G63), .ZN(new_n540));
  INV_X1    g115(.A(G651), .ZN(new_n541));
  NOR3_X1   g116(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT7), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n531), .A2(G51), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n525), .A2(new_n528), .ZN(new_n546));
  INV_X1    g121(.A(G89), .ZN(new_n547));
  OAI211_X1 g122(.A(new_n544), .B(new_n545), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n542), .A2(new_n548), .ZN(G168));
  NAND3_X1  g124(.A1(new_n537), .A2(G64), .A3(new_n538), .ZN(new_n550));
  NAND2_X1  g125(.A1(G77), .A2(G543), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n541), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n531), .A2(G52), .ZN(new_n553));
  INV_X1    g128(.A(G90), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n546), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n552), .A2(new_n555), .ZN(G171));
  NAND2_X1  g131(.A1(new_n531), .A2(G43), .ZN(new_n557));
  XNOR2_X1  g132(.A(KEYINPUT75), .B(G81), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n546), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(G68), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G56), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n539), .B2(new_n561), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n559), .B1(new_n562), .B2(G651), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G860), .ZN(G153));
  NAND4_X1  g139(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g140(.A1(G1), .A2(G3), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT8), .ZN(new_n567));
  NAND4_X1  g142(.A1(G319), .A2(G483), .A3(G661), .A4(new_n567), .ZN(G188));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n522), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n571), .A2(G651), .B1(new_n529), .B2(G91), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n531), .A2(G53), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G171), .ZN(G301));
  INV_X1    g151(.A(G168), .ZN(G286));
  INV_X1    g152(.A(KEYINPUT76), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n531), .A2(new_n578), .A3(G49), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n578), .B1(new_n531), .B2(G49), .ZN(new_n581));
  INV_X1    g156(.A(G87), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n580), .A2(new_n581), .B1(new_n582), .B2(new_n546), .ZN(new_n583));
  INV_X1    g158(.A(G74), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n541), .B1(new_n539), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT77), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n528), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G49), .ZN(new_n588));
  OAI21_X1  g163(.A(KEYINPUT76), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(new_n579), .B1(new_n529), .B2(G87), .ZN(new_n590));
  INV_X1    g165(.A(new_n538), .ZN(new_n591));
  AOI21_X1  g166(.A(KEYINPUT74), .B1(new_n520), .B2(new_n521), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n584), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G651), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT77), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n590), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n586), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G288));
  NAND2_X1  g173(.A1(new_n529), .A2(G86), .ZN(new_n599));
  NAND2_X1  g174(.A1(G73), .A2(G543), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT78), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(G61), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n520), .B2(new_n521), .ZN(new_n604));
  OAI21_X1  g179(.A(G651), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n531), .A2(G48), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n599), .A2(new_n605), .A3(new_n606), .ZN(G305));
  NAND3_X1  g182(.A1(new_n537), .A2(G60), .A3(new_n538), .ZN(new_n608));
  NAND2_X1  g183(.A1(G72), .A2(G543), .ZN(new_n609));
  AOI21_X1  g184(.A(new_n541), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n531), .A2(G47), .ZN(new_n611));
  INV_X1    g186(.A(G85), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n546), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n614), .ZN(G290));
  AND3_X1   g190(.A1(new_n525), .A2(G92), .A3(new_n528), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT10), .ZN(new_n617));
  NAND2_X1  g192(.A1(G79), .A2(G543), .ZN(new_n618));
  INV_X1    g193(.A(G66), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n522), .B2(new_n619), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n620), .A2(G651), .B1(G54), .B2(new_n531), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G868), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G171), .B2(new_n623), .ZN(G284));
  OAI21_X1  g200(.A(new_n624), .B1(G171), .B2(new_n623), .ZN(G321));
  NAND2_X1  g201(.A1(G299), .A2(new_n623), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(new_n623), .B2(G168), .ZN(G297));
  OAI21_X1  g203(.A(new_n627), .B1(new_n623), .B2(G168), .ZN(G280));
  INV_X1    g204(.A(new_n622), .ZN(new_n630));
  INV_X1    g205(.A(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(G860), .ZN(G148));
  INV_X1    g207(.A(new_n563), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(new_n623), .ZN(new_n634));
  NOR2_X1   g209(.A1(new_n622), .A2(G559), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n634), .B1(new_n635), .B2(new_n623), .ZN(G323));
  XNOR2_X1  g211(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g212(.A1(new_n490), .A2(G135), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n480), .A2(G123), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT80), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n479), .A2(G111), .ZN(new_n641));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  OAI211_X1 g217(.A(new_n638), .B(new_n640), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT81), .ZN(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n645), .A2(G2096), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(G2096), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n474), .A2(new_n465), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT12), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2100), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT79), .B(KEYINPUT13), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n646), .A2(new_n647), .A3(new_n652), .ZN(G156));
  XOR2_X1   g228(.A(KEYINPUT15), .B(G2435), .Z(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT82), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2427), .B(G2430), .Z(new_n657));
  OAI21_X1  g232(.A(KEYINPUT14), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT83), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2451), .B(G2454), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT16), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n665), .A2(new_n667), .ZN(new_n669));
  AND3_X1   g244(.A1(new_n668), .A2(G14), .A3(new_n669), .ZN(G401));
  XNOR2_X1  g245(.A(G2072), .B(G2078), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT17), .ZN(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n672), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT84), .Z(new_n677));
  NAND2_X1  g252(.A1(new_n672), .A2(new_n673), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n678), .B(new_n675), .C1(new_n671), .C2(new_n673), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n674), .A2(new_n671), .A3(new_n673), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(KEYINPUT18), .Z(new_n681));
  NAND3_X1  g256(.A1(new_n677), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G2096), .B(G2100), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(G227));
  XOR2_X1   g259(.A(G1971), .B(G1976), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT19), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1956), .B(G2474), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  AND2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT20), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n689), .ZN(new_n693));
  NOR3_X1   g268(.A1(new_n686), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n686), .B2(new_n693), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1991), .B(G1996), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT85), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n698), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n701), .B(new_n702), .Z(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(G229));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G23), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n590), .A2(new_n594), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n706), .B1(new_n708), .B2(new_n705), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT33), .B(G1976), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT86), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n705), .A2(G22), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G166), .B2(new_n705), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G1971), .ZN(new_n717));
  NOR2_X1   g292(.A1(G6), .A2(G16), .ZN(new_n718));
  INV_X1    g293(.A(G86), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n606), .B1(new_n546), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n525), .A2(G61), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n541), .B1(new_n721), .B2(new_n601), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n718), .B1(new_n723), .B2(G16), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT32), .B(G1981), .Z(new_n725));
  XOR2_X1   g300(.A(new_n724), .B(new_n725), .Z(new_n726));
  NOR4_X1   g301(.A1(new_n713), .A2(new_n714), .A3(new_n717), .A4(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT34), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  INV_X1    g305(.A(G29), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G25), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n490), .A2(G131), .ZN(new_n733));
  OAI21_X1  g308(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n734));
  INV_X1    g309(.A(G107), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n734), .B1(new_n735), .B2(G2105), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G119), .B2(new_n480), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n732), .B1(new_n739), .B2(new_n731), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT35), .B(G1991), .Z(new_n741));
  XOR2_X1   g316(.A(new_n740), .B(new_n741), .Z(new_n742));
  NAND2_X1  g317(.A1(new_n705), .A2(G24), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n614), .B2(new_n705), .ZN(new_n744));
  NOR2_X1   g319(.A1(new_n744), .A2(G1986), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n744), .A2(G1986), .ZN(new_n746));
  NOR3_X1   g321(.A1(new_n742), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n729), .A2(new_n730), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT36), .ZN(new_n749));
  OAI21_X1  g324(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n750));
  INV_X1    g325(.A(G116), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(G2105), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G128), .B2(new_n480), .ZN(new_n753));
  INV_X1    g328(.A(G140), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n753), .B1(new_n489), .B2(new_n754), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT87), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G29), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT88), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n731), .A2(G26), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT28), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G2067), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n731), .A2(G33), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n765));
  NAND3_X1  g340(.A1(new_n479), .A2(G103), .A3(G2104), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n474), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n479), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G139), .B2(new_n490), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT90), .Z(new_n771));
  AOI21_X1  g346(.A(new_n764), .B1(new_n771), .B2(G29), .ZN(new_n772));
  INV_X1    g347(.A(G2072), .ZN(new_n773));
  NOR2_X1   g348(.A1(G16), .A2(G19), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n563), .B2(G16), .ZN(new_n775));
  OAI22_X1  g350(.A1(new_n772), .A2(new_n773), .B1(G1341), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(G162), .A2(G29), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G29), .B2(G35), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G2090), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n644), .A2(G29), .ZN(new_n782));
  NOR2_X1   g357(.A1(G164), .A2(new_n731), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n783), .B1(G27), .B2(new_n731), .ZN(new_n784));
  INV_X1    g359(.A(G2078), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n781), .A2(new_n782), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT24), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n731), .B1(new_n789), .B2(G34), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n790), .A2(KEYINPUT91), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n789), .A2(G34), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n790), .B2(KEYINPUT91), .ZN(new_n793));
  OAI22_X1  g368(.A1(new_n477), .A2(new_n731), .B1(new_n791), .B2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(G2084), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n705), .A2(G21), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G168), .B2(new_n705), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n796), .B1(new_n798), .B2(G1966), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G1966), .B2(new_n798), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT31), .B(G11), .Z(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT93), .ZN(new_n802));
  INV_X1    g377(.A(G28), .ZN(new_n803));
  AOI21_X1  g378(.A(G29), .B1(new_n803), .B2(KEYINPUT30), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(KEYINPUT30), .B2(new_n803), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n794), .B2(new_n795), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n778), .B2(new_n780), .ZN(new_n808));
  NOR4_X1   g383(.A1(new_n776), .A2(new_n788), .A3(new_n800), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n705), .A2(G4), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n630), .B2(new_n705), .ZN(new_n811));
  INV_X1    g386(.A(G1348), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n772), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(G2072), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n731), .A2(G32), .ZN(new_n816));
  NAND3_X1  g391(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT26), .Z(new_n818));
  NAND2_X1  g393(.A1(new_n480), .A2(G129), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n465), .A2(G105), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n490), .B2(G141), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n816), .B1(new_n822), .B2(new_n731), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT92), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT27), .B(G1996), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n824), .A2(new_n825), .B1(G1341), .B2(new_n775), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n705), .A2(G20), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT23), .Z(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(G299), .B2(G16), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G1956), .ZN(new_n830));
  OAI211_X1 g405(.A(new_n826), .B(new_n830), .C1(new_n824), .C2(new_n825), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n705), .A2(G5), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(G171), .B2(new_n705), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G1961), .ZN(new_n834));
  NOR3_X1   g409(.A1(new_n815), .A2(new_n831), .A3(new_n834), .ZN(new_n835));
  AND4_X1   g410(.A1(new_n749), .A2(new_n763), .A3(new_n809), .A4(new_n835), .ZN(G311));
  NAND4_X1  g411(.A1(new_n749), .A2(new_n763), .A3(new_n809), .A4(new_n835), .ZN(G150));
  NAND2_X1  g412(.A1(new_n630), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT38), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n537), .A2(G67), .A3(new_n538), .ZN(new_n840));
  NAND2_X1  g415(.A1(G80), .A2(G543), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n541), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n531), .A2(G55), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT95), .B(G93), .Z(new_n844));
  OAI21_X1  g419(.A(new_n843), .B1(new_n546), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n563), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n563), .A2(new_n846), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n839), .B(new_n849), .Z(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n851));
  INV_X1    g426(.A(G860), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n846), .A2(new_n852), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT37), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(G145));
  AOI22_X1  g432(.A1(G126), .A2(new_n480), .B1(new_n510), .B2(new_n511), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n858), .A2(KEYINPUT96), .A3(new_n500), .ZN(new_n859));
  AOI21_X1  g434(.A(KEYINPUT96), .B1(new_n858), .B2(new_n500), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n756), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n822), .ZN(new_n863));
  INV_X1    g438(.A(new_n770), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n771), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n480), .A2(G130), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n479), .A2(G118), .ZN(new_n869));
  OAI21_X1  g444(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n871), .B1(new_n490), .B2(G142), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(new_n649), .Z(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n738), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n644), .B(new_n477), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(G162), .ZN(new_n877));
  INV_X1    g452(.A(new_n874), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n865), .A2(new_n878), .A3(new_n866), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n875), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(KEYINPUT97), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT97), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n875), .A2(new_n879), .A3(new_n882), .A4(new_n877), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n877), .B1(new_n875), .B2(new_n879), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n885), .A2(G37), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n884), .A2(KEYINPUT40), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT40), .B1(new_n884), .B2(new_n886), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(G395));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n849), .B(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n635), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n572), .A2(new_n574), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT99), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n895));
  NAND2_X1  g470(.A1(G299), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(new_n630), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT41), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n622), .A2(new_n895), .A3(G299), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n897), .A2(new_n899), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(KEYINPUT41), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n892), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n891), .A2(new_n635), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n891), .A2(new_n635), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(new_n901), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n614), .A2(KEYINPUT100), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n614), .A2(KEYINPUT100), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n909), .A2(new_n708), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(G303), .B(G305), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n708), .B1(new_n909), .B2(new_n910), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n913), .B1(new_n912), .B2(new_n914), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n907), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n919));
  INV_X1    g494(.A(new_n917), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n903), .A2(new_n920), .A3(new_n906), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n919), .B1(new_n918), .B2(new_n921), .ZN(new_n923));
  OAI21_X1  g498(.A(G868), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n924), .B1(G868), .B2(new_n846), .ZN(G295));
  OAI21_X1  g500(.A(new_n924), .B1(G868), .B2(new_n846), .ZN(G331));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n847), .A2(G301), .A3(new_n848), .ZN(new_n930));
  AOI21_X1  g505(.A(G301), .B1(new_n847), .B2(new_n848), .ZN(new_n931));
  OAI21_X1  g506(.A(G286), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n849), .A2(G171), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n847), .A2(G301), .A3(new_n848), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n933), .A2(G168), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n901), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n902), .A2(new_n900), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(new_n932), .A3(new_n935), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n917), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G37), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n917), .B1(new_n938), .B2(new_n940), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n929), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n900), .B(KEYINPUT102), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(new_n901), .B2(KEYINPUT41), .ZN(new_n948));
  AOI211_X1 g523(.A(KEYINPUT103), .B(new_n898), .C1(new_n897), .C2(new_n899), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n936), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n901), .B1(new_n932), .B2(new_n935), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n920), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n953), .A2(KEYINPUT43), .A3(new_n942), .A4(new_n941), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n928), .B1(new_n945), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT43), .B1(new_n943), .B2(new_n944), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n953), .A2(new_n929), .A3(new_n942), .A4(new_n941), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n928), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n927), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(KEYINPUT44), .B1(new_n957), .B2(new_n958), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n955), .A2(new_n962), .A3(KEYINPUT104), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n961), .A2(new_n963), .ZN(G397));
  NAND2_X1  g539(.A1(new_n858), .A2(new_n500), .ZN(new_n965));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT50), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n461), .B1(new_n472), .B2(new_n473), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n462), .A2(new_n463), .ZN(new_n970));
  OAI21_X1  g545(.A(G2105), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n465), .A2(G101), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n476), .A2(G40), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n466), .A2(KEYINPUT105), .A3(G40), .A4(new_n476), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n968), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT70), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n506), .ZN(new_n981));
  AOI21_X1  g556(.A(G1384), .B1(new_n981), .B2(new_n500), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(G1956), .B1(new_n977), .B2(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(new_n975), .B(new_n976), .C1(new_n982), .C2(KEYINPUT45), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n859), .A2(new_n860), .A3(G1384), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n987), .A2(KEYINPUT109), .A3(KEYINPUT45), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT96), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n965), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n858), .A2(new_n500), .A3(KEYINPUT96), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n990), .A2(KEYINPUT45), .A3(new_n966), .A4(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n986), .B1(new_n988), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g570(.A(KEYINPUT56), .B(G2072), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n985), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT57), .B1(new_n574), .B2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n999), .B(G299), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT117), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT45), .B1(new_n514), .B2(new_n966), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n975), .A2(new_n976), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(KEYINPUT109), .B1(new_n987), .B2(KEYINPUT45), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n992), .A2(new_n993), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1004), .B(new_n996), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1956), .ZN(new_n1008));
  INV_X1    g583(.A(new_n984), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n968), .A2(new_n975), .A3(new_n976), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1008), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1000), .B1(new_n1007), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT117), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n982), .A2(new_n983), .ZN(new_n1015));
  AOI21_X1  g590(.A(G1384), .B1(new_n858), .B2(new_n500), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n983), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n975), .A2(new_n1017), .A3(new_n976), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n812), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n975), .A2(new_n976), .A3(new_n1016), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(new_n762), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1001), .B(new_n1014), .C1(new_n622), .C2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1007), .A2(new_n1000), .A3(new_n1011), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1025), .A2(KEYINPUT61), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1001), .A2(new_n1027), .A3(new_n1014), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT118), .ZN(new_n1029));
  XNOR2_X1  g604(.A(KEYINPUT58), .B(G1341), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1021), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G1996), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1031), .B1(new_n995), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT59), .B1(new_n1033), .B2(new_n633), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT59), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1004), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(G1996), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1035), .B(new_n563), .C1(new_n1037), .C2(new_n1031), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT61), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1025), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(new_n1012), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1028), .A2(new_n1029), .A3(new_n1039), .A4(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n1044));
  OAI211_X1 g619(.A(new_n1044), .B(new_n630), .C1(new_n1023), .C2(KEYINPUT60), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1023), .A2(KEYINPUT60), .ZN(new_n1046));
  AOI21_X1  g621(.A(KEYINPUT60), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1047));
  OAI21_X1  g622(.A(KEYINPUT119), .B1(new_n1047), .B2(new_n622), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1045), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1046), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1043), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1000), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1025), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1040), .A2(new_n1056), .B1(new_n1034), .B2(new_n1038), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1029), .B1(new_n1057), .B2(new_n1028), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1026), .B1(new_n1052), .B2(new_n1058), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n785), .B(new_n1004), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n1061));
  INV_X1    g636(.A(G1961), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n975), .A2(new_n976), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1063), .B(new_n1017), .C1(new_n983), .C2(new_n982), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1060), .A2(new_n1061), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT45), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n967), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1067), .A2(new_n1068), .A3(new_n975), .A4(new_n976), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n982), .A2(KEYINPUT45), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1016), .A2(KEYINPUT45), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT115), .B1(new_n1003), .B2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1071), .A2(KEYINPUT53), .A3(new_n785), .A4(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(G301), .B1(new_n1065), .B2(new_n1074), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n987), .A2(KEYINPUT45), .ZN(new_n1076));
  NOR3_X1   g651(.A1(new_n973), .A2(new_n1061), .A3(G2078), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1076), .B(new_n1077), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT122), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n988), .A2(new_n994), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1080), .A2(new_n1081), .A3(new_n1076), .A4(new_n1077), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1083), .A2(G301), .A3(new_n1065), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1075), .B1(new_n1084), .B2(KEYINPUT123), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT123), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1083), .A2(new_n1086), .A3(G301), .A4(new_n1065), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT54), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G1976), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n586), .A2(new_n596), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT52), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1020), .B(G8), .C1(new_n1089), .C2(new_n707), .ZN(new_n1093));
  OR2_X1    g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  XNOR2_X1  g669(.A(KEYINPUT112), .B(G1981), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n599), .A2(new_n605), .A3(new_n606), .A4(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(G1981), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1097), .B(KEYINPUT113), .C1(new_n723), .C2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT113), .ZN(new_n1100));
  NAND3_X1  g675(.A1(G305), .A2(new_n1100), .A3(G1981), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(KEYINPUT49), .ZN(new_n1103));
  INV_X1    g678(.A(G8), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1021), .A2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT49), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1099), .A2(new_n1106), .A3(new_n1101), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1103), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1093), .A2(KEYINPUT111), .A3(KEYINPUT52), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT111), .B1(new_n1093), .B2(KEYINPUT52), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1094), .B(new_n1108), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(G166), .A2(new_n1104), .ZN(new_n1112));
  NAND2_X1  g687(.A1(KEYINPUT110), .A2(KEYINPUT55), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(KEYINPUT110), .A2(KEYINPUT55), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1115), .B1(new_n1112), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  OR2_X1    g695(.A1(new_n1064), .A2(G2090), .ZN(new_n1121));
  INV_X1    g696(.A(G1971), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1036), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1104), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1111), .B1(new_n1120), .B2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1123), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n1009), .A2(new_n1010), .A3(G2090), .ZN(new_n1127));
  OAI21_X1  g702(.A(G8), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(new_n1119), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1065), .A2(G301), .A3(new_n1074), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(KEYINPUT54), .ZN(new_n1131));
  AOI21_X1  g706(.A(G301), .B1(new_n1083), .B2(new_n1065), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1125), .B(new_n1129), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1015), .A2(new_n1018), .A3(G2084), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1073), .A2(new_n1070), .A3(new_n1069), .ZN(new_n1135));
  INV_X1    g710(.A(G1966), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NOR3_X1   g712(.A1(new_n1137), .A2(new_n1104), .A3(G168), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT121), .B1(new_n1137), .B2(new_n1104), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT121), .ZN(new_n1140));
  AOI21_X1  g715(.A(G1966), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1140), .B(G8), .C1(new_n1141), .C2(new_n1134), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1139), .A2(new_n1142), .A3(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1104), .B1(new_n1137), .B2(G168), .ZN(new_n1145));
  XNOR2_X1  g720(.A(KEYINPUT120), .B(KEYINPUT51), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1138), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n1088), .A2(new_n1133), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1059), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n1151));
  OR2_X1    g726(.A1(new_n1148), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1148), .A2(new_n1151), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1125), .A2(new_n1129), .A3(new_n1075), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1152), .A2(KEYINPUT124), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1154), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1153), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1156), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n597), .A2(new_n1089), .ZN(new_n1160));
  XOR2_X1   g735(.A(new_n1160), .B(KEYINPUT114), .Z(new_n1161));
  AND2_X1   g736(.A1(new_n1103), .A2(new_n1107), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1097), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n1105), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1124), .A2(new_n1120), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1164), .B1(new_n1165), .B2(new_n1111), .ZN(new_n1166));
  NOR3_X1   g741(.A1(new_n1137), .A2(new_n1104), .A3(G286), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1125), .A2(new_n1129), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT63), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OR2_X1    g745(.A1(new_n1124), .A2(new_n1120), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1125), .A2(new_n1171), .A3(KEYINPUT63), .A4(new_n1167), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1166), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1150), .A2(new_n1155), .A3(new_n1159), .A4(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n756), .B(new_n762), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n987), .A2(KEYINPUT45), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(new_n1063), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  XOR2_X1   g753(.A(new_n1178), .B(KEYINPUT108), .Z(new_n1179));
  NOR2_X1   g754(.A1(new_n1177), .A2(G1996), .ZN(new_n1180));
  XOR2_X1   g755(.A(new_n1180), .B(KEYINPUT107), .Z(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n822), .ZN(new_n1182));
  OR3_X1    g757(.A1(new_n1177), .A2(new_n1032), .A3(new_n822), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1179), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1177), .ZN(new_n1185));
  XOR2_X1   g760(.A(new_n738), .B(new_n741), .Z(new_n1186));
  AOI21_X1  g761(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  OR2_X1    g762(.A1(G290), .A2(G1986), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT106), .ZN(new_n1189));
  NAND2_X1  g764(.A1(G290), .A2(G1986), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  OAI211_X1 g766(.A(new_n1191), .B(new_n1185), .C1(new_n1189), .C2(new_n1190), .ZN(new_n1192));
  AND2_X1   g767(.A1(new_n1187), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1174), .A2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1188), .A2(new_n1177), .ZN(new_n1195));
  XOR2_X1   g770(.A(new_n1195), .B(KEYINPUT48), .Z(new_n1196));
  NAND2_X1  g771(.A1(new_n739), .A2(new_n741), .ZN(new_n1197));
  OAI22_X1  g772(.A1(new_n1184), .A2(new_n1197), .B1(G2067), .B2(new_n756), .ZN(new_n1198));
  AOI22_X1  g773(.A1(new_n1187), .A2(new_n1196), .B1(new_n1198), .B2(new_n1185), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT125), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1201), .B1(new_n1181), .B2(KEYINPUT46), .ZN(new_n1202));
  XNOR2_X1  g777(.A(new_n1180), .B(KEYINPUT107), .ZN(new_n1203));
  INV_X1    g778(.A(KEYINPUT46), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1203), .A2(KEYINPUT125), .A3(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1202), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1177), .B1(new_n1175), .B2(new_n822), .ZN(new_n1207));
  AOI21_X1  g782(.A(new_n1207), .B1(new_n1181), .B2(KEYINPUT46), .ZN(new_n1208));
  NAND3_X1  g783(.A1(new_n1206), .A2(KEYINPUT47), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g784(.A(new_n1209), .ZN(new_n1210));
  AOI21_X1  g785(.A(KEYINPUT47), .B1(new_n1206), .B2(new_n1208), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1200), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  INV_X1    g787(.A(new_n1211), .ZN(new_n1213));
  NAND3_X1  g788(.A1(new_n1213), .A2(KEYINPUT126), .A3(new_n1209), .ZN(new_n1214));
  AND3_X1   g789(.A1(new_n1199), .A2(new_n1212), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1194), .A2(new_n1215), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g791(.A1(new_n884), .A2(new_n886), .ZN(new_n1218));
  INV_X1    g792(.A(G319), .ZN(new_n1219));
  NOR2_X1   g793(.A1(G227), .A2(new_n1219), .ZN(new_n1220));
  XOR2_X1   g794(.A(new_n1220), .B(KEYINPUT127), .Z(new_n1221));
  NOR3_X1   g795(.A1(G401), .A2(G229), .A3(new_n1221), .ZN(new_n1222));
  NAND3_X1  g796(.A1(new_n1218), .A2(new_n1222), .A3(new_n959), .ZN(G225));
  INV_X1    g797(.A(G225), .ZN(G308));
endmodule


