//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 0 1 0 1 0 1 0 0 1 1 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965;
  INV_X1    g000(.A(G237), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT68), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT68), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G237), .ZN(new_n190));
  AOI21_X1  g004(.A(G953), .B1(new_n188), .B2(new_n190), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G210), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT70), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n194), .B(KEYINPUT69), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT26), .B(G101), .ZN(new_n196));
  XOR2_X1   g010(.A(new_n196), .B(KEYINPUT27), .Z(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT69), .ZN(new_n199));
  XNOR2_X1  g013(.A(new_n194), .B(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(new_n197), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G137), .ZN(new_n206));
  INV_X1    g020(.A(G137), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT11), .A3(G134), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(G137), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G131), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n206), .A2(new_n208), .A3(new_n212), .A4(new_n209), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G143), .ZN(new_n216));
  INV_X1    g030(.A(G143), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G146), .ZN(new_n218));
  AND2_X1   g032(.A1(KEYINPUT0), .A2(G128), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(G143), .B(G146), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT0), .B(G128), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n220), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n214), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT1), .B1(new_n217), .B2(G146), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n217), .A2(G146), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n215), .A2(G143), .ZN(new_n228));
  OAI211_X1 g042(.A(G128), .B(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n205), .A2(G137), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n207), .A2(G134), .ZN(new_n231));
  OAI21_X1  g045(.A(G131), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G128), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n216), .B(new_n218), .C1(KEYINPUT1), .C2(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n229), .A2(new_n213), .A3(new_n232), .A4(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n225), .A2(new_n235), .ZN(new_n236));
  XOR2_X1   g050(.A(KEYINPUT2), .B(G113), .Z(new_n237));
  XNOR2_X1  g051(.A(G116), .B(G119), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G119), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G116), .ZN(new_n241));
  INV_X1    g055(.A(G116), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G119), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n244), .A2(KEYINPUT65), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT65), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n238), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n239), .B1(new_n248), .B2(new_n237), .ZN(new_n249));
  OR3_X1    g063(.A1(new_n236), .A2(KEYINPUT67), .A3(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT67), .B1(new_n236), .B2(new_n249), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n223), .B1(new_n211), .B2(new_n213), .ZN(new_n254));
  INV_X1    g068(.A(new_n235), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT64), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT30), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n236), .A2(KEYINPUT64), .A3(KEYINPUT30), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n253), .B1(new_n260), .B2(new_n249), .ZN(new_n261));
  INV_X1    g075(.A(new_n249), .ZN(new_n262));
  AOI211_X1 g076(.A(KEYINPUT66), .B(new_n262), .C1(new_n258), .C2(new_n259), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n203), .B(new_n252), .C1(new_n261), .C2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT31), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT30), .B1(new_n236), .B2(KEYINPUT64), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT64), .ZN(new_n267));
  AOI211_X1 g081(.A(new_n267), .B(new_n257), .C1(new_n225), .C2(new_n235), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n249), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT66), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n260), .A2(new_n253), .A3(new_n249), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT31), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n272), .A2(new_n273), .A3(new_n203), .A4(new_n252), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n249), .B1(new_n236), .B2(KEYINPUT71), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n275), .B1(KEYINPUT71), .B2(new_n236), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT28), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n250), .A2(new_n251), .B1(new_n249), .B2(new_n236), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n278), .B1(new_n279), .B2(new_n277), .ZN(new_n280));
  INV_X1    g094(.A(new_n203), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n265), .A2(new_n274), .A3(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(G472), .A2(G902), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT32), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n283), .A2(KEYINPUT32), .A3(new_n284), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n287), .A2(KEYINPUT72), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT72), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n283), .A2(new_n290), .A3(KEYINPUT32), .A4(new_n284), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n272), .A2(new_n252), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n281), .ZN(new_n293));
  OR2_X1    g107(.A1(new_n280), .A2(new_n281), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT29), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n296), .B(new_n297), .C1(new_n295), .C2(new_n294), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n289), .A2(new_n291), .B1(G472), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(G217), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n300), .B1(G234), .B2(new_n297), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT25), .ZN(new_n303));
  XNOR2_X1  g117(.A(G125), .B(G140), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT16), .ZN(new_n305));
  INV_X1    g119(.A(G125), .ZN(new_n306));
  OR3_X1    g120(.A1(new_n306), .A2(KEYINPUT16), .A3(G140), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n215), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n305), .A2(G146), .A3(new_n307), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT23), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n312), .B1(G119), .B2(new_n233), .ZN(new_n313));
  NOR3_X1   g127(.A1(new_n240), .A2(KEYINPUT23), .A3(G128), .ZN(new_n314));
  OAI22_X1  g128(.A1(new_n313), .A2(new_n314), .B1(G119), .B2(new_n233), .ZN(new_n315));
  XNOR2_X1  g129(.A(G119), .B(G128), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT24), .B(G110), .Z(new_n317));
  AOI22_X1  g131(.A1(new_n315), .A2(G110), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n311), .A2(new_n318), .ZN(new_n319));
  OAI22_X1  g133(.A1(new_n315), .A2(G110), .B1(new_n316), .B2(new_n317), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n304), .A2(new_n215), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n310), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT22), .B(G137), .ZN(new_n324));
  INV_X1    g138(.A(G953), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(G221), .A3(G234), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n324), .B(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n327), .B(KEYINPUT73), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n323), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n319), .A2(new_n322), .A3(new_n327), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n303), .B1(new_n332), .B2(G902), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n330), .A2(KEYINPUT25), .A3(new_n297), .A4(new_n331), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n302), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n301), .A2(G902), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n299), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n188), .A2(new_n190), .ZN(new_n342));
  AND4_X1   g156(.A1(G143), .A2(new_n342), .A3(G214), .A4(new_n325), .ZN(new_n343));
  AOI21_X1  g157(.A(G143), .B1(new_n191), .B2(G214), .ZN(new_n344));
  OAI211_X1 g158(.A(KEYINPUT18), .B(G131), .C1(new_n343), .C2(new_n344), .ZN(new_n345));
  OR2_X1    g159(.A1(new_n304), .A2(new_n215), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n321), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n189), .A2(G237), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n187), .A2(KEYINPUT68), .ZN(new_n350));
  OAI211_X1 g164(.A(G214), .B(new_n325), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n217), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n191), .A2(G143), .A3(G214), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT18), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n352), .B(new_n353), .C1(new_n354), .C2(new_n212), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n355), .A2(KEYINPUT84), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(KEYINPUT84), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n348), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n352), .A2(new_n353), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n359), .A2(G131), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n212), .B1(new_n352), .B2(new_n353), .ZN(new_n361));
  OR3_X1    g175(.A1(new_n360), .A2(KEYINPUT17), .A3(new_n361), .ZN(new_n362));
  OAI211_X1 g176(.A(KEYINPUT17), .B(G131), .C1(new_n343), .C2(new_n344), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT86), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n359), .A2(KEYINPUT86), .A3(KEYINPUT17), .A4(G131), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n311), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n362), .B1(new_n367), .B2(KEYINPUT87), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT87), .ZN(new_n369));
  AOI211_X1 g183(.A(new_n369), .B(new_n311), .C1(new_n365), .C2(new_n366), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n358), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(G113), .B(G122), .ZN(new_n372));
  INV_X1    g186(.A(G104), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n372), .B(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n374), .B(new_n358), .C1(new_n368), .C2(new_n370), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(G475), .B1(new_n378), .B2(G902), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n345), .A2(new_n347), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n343), .A2(new_n344), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT84), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n381), .B(new_n382), .C1(new_n354), .C2(new_n212), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n355), .A2(KEYINPUT84), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n380), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  XOR2_X1   g199(.A(new_n304), .B(KEYINPUT19), .Z(new_n386));
  OAI21_X1  g200(.A(new_n310), .B1(new_n386), .B2(G146), .ZN(new_n387));
  INV_X1    g201(.A(new_n360), .ZN(new_n388));
  INV_X1    g202(.A(new_n361), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n387), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT85), .B1(new_n385), .B2(new_n390), .ZN(new_n391));
  OAI221_X1 g205(.A(new_n310), .B1(G146), .B2(new_n386), .C1(new_n360), .C2(new_n361), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT85), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n358), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(new_n394), .A3(new_n375), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n377), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT88), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT20), .ZN(new_n398));
  NOR2_X1   g212(.A1(G475), .A2(G902), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n396), .A2(new_n397), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n399), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n401), .B1(new_n377), .B2(new_n395), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n400), .B1(new_n398), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n397), .B1(new_n402), .B2(new_n398), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n379), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT89), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n396), .A2(new_n398), .A3(new_n399), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT88), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n396), .A2(new_n399), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(KEYINPUT20), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n400), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT89), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n411), .A2(new_n412), .A3(new_n379), .ZN(new_n413));
  INV_X1    g227(.A(G478), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(KEYINPUT15), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT9), .B(G234), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n417), .B(KEYINPUT74), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(G217), .A3(new_n325), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n242), .A2(G122), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT90), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n421), .A2(new_n242), .A3(G122), .ZN(new_n422));
  INV_X1    g236(.A(G122), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT90), .B1(new_n423), .B2(G116), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n420), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT91), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n425), .A2(KEYINPUT91), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(G107), .ZN(new_n430));
  INV_X1    g244(.A(G107), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n431), .B1(new_n427), .B2(new_n428), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n217), .A2(G128), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n217), .A2(G128), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AND2_X1   g251(.A1(new_n437), .A2(new_n205), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT13), .ZN(new_n439));
  OR3_X1    g253(.A1(new_n436), .A2(KEYINPUT92), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n434), .B1(new_n439), .B2(new_n436), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT92), .B1(new_n436), .B2(new_n439), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n438), .B1(new_n443), .B2(G134), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n433), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n437), .A2(new_n205), .ZN(new_n447));
  OR2_X1    g261(.A1(new_n438), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n420), .B(KEYINPUT14), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n422), .A2(new_n424), .ZN(new_n450));
  OAI21_X1  g264(.A(G107), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  OR2_X1    g265(.A1(new_n451), .A2(KEYINPUT94), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(KEYINPUT94), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n448), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n432), .A2(KEYINPUT93), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n432), .A2(KEYINPUT93), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n454), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n419), .B1(new_n446), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n419), .ZN(new_n460));
  INV_X1    g274(.A(new_n457), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(new_n455), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n460), .B(new_n445), .C1(new_n462), .C2(new_n454), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n416), .B1(new_n464), .B2(new_n297), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n464), .A2(new_n297), .A3(new_n416), .ZN(new_n467));
  AND2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(G234), .A2(G237), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n469), .A2(G952), .A3(new_n325), .ZN(new_n470));
  XOR2_X1   g284(.A(KEYINPUT21), .B(G898), .Z(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n469), .A2(G902), .A3(G953), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AND4_X1   g289(.A1(new_n406), .A2(new_n413), .A3(new_n468), .A4(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n418), .ZN(new_n477));
  OAI21_X1  g291(.A(G221), .B1(new_n477), .B2(G902), .ZN(new_n478));
  XOR2_X1   g292(.A(new_n478), .B(KEYINPUT75), .Z(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G469), .ZN(new_n481));
  XNOR2_X1  g295(.A(G110), .B(G140), .ZN(new_n482));
  INV_X1    g296(.A(G227), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n483), .A2(G953), .ZN(new_n484));
  XOR2_X1   g298(.A(new_n482), .B(new_n484), .Z(new_n485));
  NAND2_X1  g299(.A1(new_n431), .A2(G104), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n373), .A2(G107), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(G101), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT78), .ZN(new_n490));
  INV_X1    g304(.A(G101), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT3), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n431), .A3(G104), .ZN(new_n493));
  AOI21_X1  g307(.A(KEYINPUT3), .B1(new_n373), .B2(G107), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n373), .A2(G107), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n491), .B(new_n493), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT78), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n488), .A2(new_n497), .A3(G101), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n490), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT79), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n490), .A2(KEYINPUT79), .A3(new_n498), .A4(new_n496), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n229), .A2(new_n234), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT10), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n504), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n508), .A2(new_n496), .A3(new_n490), .A4(new_n498), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n505), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT77), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G101), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(KEYINPUT76), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT76), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n516), .B(new_n493), .C1(new_n494), .C2(new_n495), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n513), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n518), .A2(KEYINPUT4), .ZN(new_n519));
  INV_X1    g333(.A(new_n496), .ZN(new_n520));
  OAI21_X1  g334(.A(KEYINPUT4), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n223), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n214), .B1(new_n511), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT81), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n519), .A2(new_n521), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n224), .ZN(new_n527));
  AOI22_X1  g341(.A1(new_n503), .A2(new_n506), .B1(new_n509), .B2(new_n505), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(KEYINPUT81), .A3(new_n214), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n214), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n527), .A2(new_n528), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n485), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n499), .A2(new_n504), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n499), .A2(new_n504), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n214), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT80), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT12), .B1(new_n214), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n537), .B(new_n539), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n540), .A2(new_n533), .A3(new_n485), .ZN(new_n541));
  OAI211_X1 g355(.A(new_n481), .B(new_n297), .C1(new_n534), .C2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n485), .B1(new_n540), .B2(new_n533), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n533), .A2(new_n485), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n543), .B1(new_n531), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(G469), .B1(new_n545), .B2(G902), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n480), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(G210), .B1(G237), .B2(G902), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n526), .A2(new_n249), .ZN(new_n550));
  OAI21_X1  g364(.A(G113), .B1(new_n241), .B2(KEYINPUT5), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT5), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n245), .A2(new_n247), .A3(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n503), .B(new_n239), .C1(new_n551), .C2(new_n553), .ZN(new_n554));
  XOR2_X1   g368(.A(G110), .B(G122), .Z(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n550), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n262), .B1(new_n519), .B2(new_n521), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n239), .B1(new_n553), .B2(new_n551), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n559), .B1(new_n501), .B2(new_n502), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n555), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n557), .A2(new_n561), .A3(KEYINPUT6), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT6), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n563), .B(new_n555), .C1(new_n558), .C2(new_n560), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n223), .A2(G125), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n565), .B1(new_n508), .B2(G125), .ZN(new_n566));
  INV_X1    g380(.A(G224), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(G953), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n566), .B(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n562), .A2(new_n564), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT7), .ZN(new_n571));
  OAI221_X1 g385(.A(new_n565), .B1(KEYINPUT82), .B2(new_n571), .C1(new_n508), .C2(G125), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n568), .A2(new_n571), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n499), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n244), .A2(new_n552), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n239), .B1(new_n577), .B2(new_n551), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g393(.A(new_n555), .B(KEYINPUT8), .Z(new_n580));
  OAI211_X1 g394(.A(new_n579), .B(new_n580), .C1(new_n559), .C2(new_n576), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n572), .A2(new_n574), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n575), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(G902), .B1(new_n583), .B2(new_n557), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n549), .B1(new_n570), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT83), .ZN(new_n586));
  INV_X1    g400(.A(new_n585), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n570), .A2(new_n549), .A3(new_n584), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n586), .B1(new_n589), .B2(KEYINPUT83), .ZN(new_n590));
  OAI21_X1  g404(.A(G214), .B1(G237), .B2(G902), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n548), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n341), .A2(new_n476), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G101), .ZN(G3));
  NAND3_X1  g409(.A1(new_n547), .A2(new_n339), .A3(new_n475), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n592), .B1(new_n587), .B2(new_n588), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  AOI22_X1  g412(.A1(new_n264), .A2(KEYINPUT31), .B1(new_n280), .B2(new_n281), .ZN(new_n599));
  AOI21_X1  g413(.A(G902), .B1(new_n599), .B2(new_n274), .ZN(new_n600));
  INV_X1    g414(.A(G472), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n285), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OR3_X1    g416(.A1(new_n596), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(G478), .B1(new_n464), .B2(new_n297), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n464), .A2(KEYINPUT95), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT33), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n464), .A2(KEYINPUT95), .A3(KEYINPUT33), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n414), .A2(G902), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n604), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n406), .B2(new_n413), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n603), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT34), .B(G104), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  NAND2_X1  g430(.A1(new_n466), .A2(new_n467), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n410), .A2(new_n407), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n617), .A2(new_n618), .A3(new_n379), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n603), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT35), .B(G107), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G9));
  AND2_X1   g436(.A1(new_n476), .A2(new_n593), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n333), .A2(new_n334), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n301), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT36), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n328), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(new_n323), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n628), .A2(new_n337), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT96), .B1(new_n625), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT96), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n335), .A2(new_n632), .A3(new_n629), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n602), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n623), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT37), .B(G110), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G12));
  NOR2_X1   g451(.A1(new_n631), .A2(new_n633), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n547), .A2(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n299), .A2(new_n598), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(G900), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n473), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n470), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n619), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(new_n233), .ZN(G30));
  XOR2_X1   g462(.A(new_n590), .B(KEYINPUT38), .Z(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n644), .B(KEYINPUT39), .Z(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n547), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(KEYINPUT40), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n468), .B1(new_n406), .B2(new_n413), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n289), .A2(new_n291), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n292), .A2(new_n203), .ZN(new_n658));
  AOI21_X1  g472(.A(G902), .B1(new_n281), .B2(new_n279), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n657), .B1(new_n601), .B2(new_n660), .ZN(new_n661));
  AOI211_X1 g475(.A(new_n592), .B(new_n638), .C1(new_n653), .C2(KEYINPUT40), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n655), .A2(new_n656), .A3(new_n661), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G143), .ZN(G45));
  AOI211_X1 g478(.A(new_n611), .B(new_n645), .C1(new_n406), .C2(new_n413), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n640), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G146), .ZN(G48));
  NAND2_X1  g481(.A1(new_n597), .A2(new_n475), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n613), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(KEYINPUT81), .B1(new_n529), .B2(new_n214), .ZN(new_n670));
  AOI211_X1 g484(.A(new_n524), .B(new_n532), .C1(new_n527), .C2(new_n528), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n533), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n485), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n541), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(G469), .B1(new_n674), .B2(G902), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n675), .A2(new_n478), .A3(new_n542), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n299), .A2(new_n340), .A3(new_n677), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n669), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT41), .B(G113), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G15));
  NOR2_X1   g495(.A1(new_n668), .A2(new_n619), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G116), .ZN(G18));
  INV_X1    g498(.A(new_n299), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n597), .A2(new_n675), .A3(new_n478), .A4(new_n542), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n685), .A2(new_n476), .A3(new_n638), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G119), .ZN(G21));
  NAND2_X1  g503(.A1(new_n283), .A2(new_n297), .ZN(new_n690));
  XOR2_X1   g504(.A(new_n284), .B(KEYINPUT97), .Z(new_n691));
  AOI22_X1  g505(.A1(new_n690), .A2(G472), .B1(new_n283), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n677), .A2(new_n668), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n656), .A2(new_n339), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G122), .ZN(G24));
  INV_X1    g509(.A(KEYINPUT98), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n609), .A2(new_n610), .ZN(new_n697));
  INV_X1    g511(.A(new_n604), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n411), .A2(new_n412), .A3(new_n379), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n412), .B1(new_n411), .B2(new_n379), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n699), .B(new_n644), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n676), .A2(new_n597), .A3(new_n638), .A4(new_n692), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n696), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n283), .A2(new_n691), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n638), .B(new_n705), .C1(new_n601), .C2(new_n600), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n686), .A2(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n612), .A2(new_n707), .A3(KEYINPUT98), .A4(new_n644), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G125), .ZN(G27));
  INV_X1    g524(.A(new_n588), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n711), .A2(new_n585), .A3(KEYINPUT83), .ZN(new_n712));
  INV_X1    g526(.A(new_n586), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n591), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(KEYINPUT99), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT99), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n590), .A2(new_n716), .A3(new_n591), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n542), .A2(new_n546), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n715), .A2(new_n717), .A3(new_n478), .A4(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n702), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT42), .B1(new_n720), .B2(new_n341), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT101), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n287), .B(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n298), .A2(G472), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT100), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n288), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n288), .A2(new_n725), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n724), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI211_X1 g542(.A(KEYINPUT42), .B(new_n339), .C1(new_n723), .C2(new_n728), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n729), .A2(new_n702), .A3(new_n719), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n721), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n212), .ZN(G33));
  NAND2_X1  g546(.A1(new_n341), .A2(new_n646), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n719), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(new_n205), .ZN(G36));
  NAND2_X1  g549(.A1(new_n715), .A2(new_n717), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n406), .A2(new_n413), .A3(new_n699), .ZN(new_n737));
  XOR2_X1   g551(.A(new_n737), .B(KEYINPUT43), .Z(new_n738));
  INV_X1    g552(.A(KEYINPUT103), .ZN(new_n739));
  OR2_X1    g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n739), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n740), .A2(new_n602), .A3(new_n638), .A4(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n736), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g558(.A(new_n744), .B1(new_n743), .B2(new_n742), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT104), .ZN(new_n746));
  OR2_X1    g560(.A1(new_n545), .A2(KEYINPUT45), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n545), .A2(KEYINPUT45), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(G469), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(G469), .A2(G902), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(KEYINPUT46), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n542), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT46), .B1(new_n749), .B2(new_n750), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n478), .A3(new_n652), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT102), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n746), .A2(new_n756), .ZN(new_n757));
  XOR2_X1   g571(.A(KEYINPUT105), .B(G137), .Z(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G39));
  NAND2_X1  g573(.A1(new_n754), .A2(new_n478), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT47), .ZN(new_n761));
  INV_X1    g575(.A(new_n736), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n762), .A2(new_n299), .A3(new_n340), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n761), .A2(new_n702), .A3(new_n763), .ZN(new_n764));
  XOR2_X1   g578(.A(new_n764), .B(KEYINPUT106), .Z(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G140), .ZN(G42));
  NAND3_X1  g580(.A1(new_n650), .A2(new_n591), .A3(new_n479), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n675), .A2(new_n542), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT107), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n767), .B1(KEYINPUT49), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(KEYINPUT49), .ZN(new_n771));
  XOR2_X1   g585(.A(new_n771), .B(KEYINPUT108), .Z(new_n772));
  NOR3_X1   g586(.A1(new_n661), .A2(new_n340), .A3(new_n737), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n770), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n736), .A2(new_n643), .A3(new_n677), .ZN(new_n775));
  INV_X1    g589(.A(new_n661), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n339), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n406), .A2(new_n413), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n777), .A2(new_n778), .A3(new_n699), .ZN(new_n779));
  INV_X1    g593(.A(new_n706), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n738), .A2(new_n775), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AND4_X1   g596(.A1(new_n339), .A2(new_n738), .A3(new_n470), .A4(new_n692), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n783), .A2(new_n592), .A3(new_n650), .A4(new_n676), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT50), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n784), .A2(new_n785), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n782), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n761), .B1(new_n479), .B2(new_n769), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n762), .A3(new_n783), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n788), .A2(new_n789), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n790), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n796), .A2(KEYINPUT115), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(KEYINPUT115), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n639), .B1(new_n657), .B2(new_n724), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n597), .B(new_n800), .C1(new_n665), .C2(new_n646), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n335), .A2(new_n629), .A3(new_n645), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n718), .A2(new_n478), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT110), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n718), .A2(KEYINPUT110), .A3(new_n478), .A4(new_n802), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n661), .A2(new_n807), .A3(new_n597), .A4(new_n656), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n709), .A2(new_n801), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT111), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT111), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n709), .A2(new_n801), .A3(new_n811), .A4(new_n808), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n799), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n594), .A2(new_n688), .A3(new_n694), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n623), .A2(new_n634), .B1(new_n669), .B2(new_n678), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n613), .B1(new_n778), .B2(new_n468), .ZN(new_n817));
  NOR4_X1   g631(.A1(new_n596), .A2(new_n590), .A3(new_n602), .A4(new_n592), .ZN(new_n818));
  AOI22_X1  g632(.A1(new_n817), .A2(new_n818), .B1(new_n678), .B2(new_n682), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT109), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n468), .A2(new_n644), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n618), .A2(new_n379), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n617), .A2(new_n645), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n824), .A2(new_n618), .A3(KEYINPUT109), .A4(new_n379), .ZN(new_n825));
  AND4_X1   g639(.A1(new_n715), .A2(new_n823), .A3(new_n717), .A4(new_n825), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n720), .A2(new_n780), .B1(new_n826), .B2(new_n800), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n815), .A2(new_n816), .A3(new_n819), .A4(new_n827), .ZN(new_n828));
  OAI22_X1  g642(.A1(new_n721), .A2(new_n730), .B1(new_n719), .B2(new_n733), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n810), .A2(new_n799), .A3(new_n812), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n814), .A2(new_n830), .A3(KEYINPUT53), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n830), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n809), .A2(KEYINPUT52), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT112), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n831), .A2(KEYINPUT112), .A3(new_n834), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n833), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n832), .B1(new_n839), .B2(KEYINPUT53), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT54), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n831), .A2(KEYINPUT112), .A3(new_n834), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT112), .B1(new_n831), .B2(new_n834), .ZN(new_n843));
  OAI211_X1 g657(.A(KEYINPUT53), .B(new_n830), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n814), .A2(new_n830), .A3(new_n831), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n844), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT113), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n841), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n840), .A2(new_n850), .A3(KEYINPUT54), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(G952), .B(new_n325), .C1(new_n777), .C2(new_n613), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n783), .B2(new_n687), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n723), .A2(new_n728), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n857), .A2(new_n340), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n781), .A2(new_n858), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(KEYINPUT116), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT48), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n859), .A2(KEYINPUT116), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n856), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n864), .B1(new_n862), .B2(new_n863), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n792), .A2(KEYINPUT51), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n865), .B1(new_n788), .B2(new_n866), .ZN(new_n867));
  NOR4_X1   g681(.A1(new_n797), .A2(new_n798), .A3(new_n854), .A4(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(G952), .A2(G953), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n774), .B1(new_n868), .B2(new_n869), .ZN(G75));
  AOI21_X1  g684(.A(new_n297), .B1(new_n844), .B2(new_n848), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT56), .B1(new_n871), .B2(G210), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n562), .A2(new_n564), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(new_n569), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT55), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n872), .A2(new_n875), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n325), .A2(G952), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(G51));
  NAND2_X1  g693(.A1(new_n844), .A2(new_n848), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT54), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n882), .A3(new_n849), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n880), .A2(KEYINPUT117), .A3(KEYINPUT54), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n750), .B(KEYINPUT57), .ZN(new_n886));
  OAI22_X1  g700(.A1(new_n885), .A2(new_n886), .B1(new_n534), .B2(new_n541), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n871), .A2(G469), .A3(new_n748), .A4(new_n747), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n878), .B1(new_n887), .B2(new_n888), .ZN(G54));
  AND3_X1   g703(.A1(new_n871), .A2(KEYINPUT58), .A3(G475), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n890), .A2(new_n396), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n891), .A2(KEYINPUT118), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n891), .A2(KEYINPUT118), .ZN(new_n893));
  INV_X1    g707(.A(new_n878), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n894), .B1(new_n890), .B2(new_n396), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(G60));
  NAND2_X1  g710(.A1(G478), .A2(G902), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT59), .Z(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n883), .A2(new_n609), .A3(new_n884), .A4(new_n899), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n900), .A2(new_n894), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n898), .B1(new_n852), .B2(new_n853), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n902), .A2(new_n903), .A3(new_n609), .ZN(new_n904));
  AOI22_X1  g718(.A1(KEYINPUT54), .A2(new_n840), .B1(new_n849), .B2(new_n850), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n830), .B1(new_n842), .B2(new_n843), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n847), .ZN(new_n907));
  AOI211_X1 g721(.A(KEYINPUT113), .B(new_n845), .C1(new_n907), .C2(new_n832), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n899), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(new_n609), .ZN(new_n910));
  AOI21_X1  g724(.A(KEYINPUT119), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n901), .B1(new_n904), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT120), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n901), .B(KEYINPUT120), .C1(new_n904), .C2(new_n911), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(G63));
  NAND2_X1  g730(.A1(G217), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT121), .Z(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT60), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n844), .B2(new_n848), .ZN(new_n920));
  INV_X1    g734(.A(new_n628), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n878), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n332), .B(KEYINPUT122), .Z(new_n923));
  OAI21_X1  g737(.A(new_n922), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n924), .B(KEYINPUT61), .Z(G66));
  NAND3_X1  g739(.A1(new_n815), .A2(new_n816), .A3(new_n819), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n325), .ZN(new_n927));
  OAI21_X1  g741(.A(G953), .B1(new_n472), .B2(new_n567), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n873), .B1(G898), .B2(new_n325), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(G69));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n709), .A2(new_n801), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n756), .A2(new_n597), .A3(new_n656), .A4(new_n858), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT125), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n765), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(new_n829), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n757), .A2(new_n937), .A3(new_n325), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n260), .B(new_n386), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(G900), .B2(G953), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n663), .B(new_n933), .C1(KEYINPUT123), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(KEYINPUT123), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n943), .B(new_n944), .Z(new_n945));
  NAND4_X1  g759(.A1(new_n341), .A2(new_n762), .A3(new_n547), .A4(new_n652), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT124), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(new_n817), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n948), .B1(new_n947), .B2(new_n817), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n765), .A2(new_n945), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(new_n746), .B2(new_n756), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n939), .B1(new_n951), .B2(G953), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n932), .B1(new_n941), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n483), .B1(new_n939), .B2(KEYINPUT126), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n325), .B1(new_n954), .B2(G900), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n953), .B(new_n955), .ZN(G72));
  NAND3_X1  g770(.A1(new_n951), .A2(new_n203), .A3(new_n292), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n292), .A2(new_n203), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n757), .A2(new_n937), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n926), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(G472), .A2(G902), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT63), .Z(new_n962));
  NAND2_X1  g776(.A1(new_n293), .A2(new_n264), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n840), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n894), .B1(new_n963), .B2(new_n962), .ZN(new_n965));
  NOR3_X1   g779(.A1(new_n960), .A2(new_n964), .A3(new_n965), .ZN(G57));
endmodule


