//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n822, new_n823, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948;
  OR2_X1    g000(.A1(G57gat), .A2(G64gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G57gat), .A2(G64gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g003(.A1(G71gat), .A2(G78gat), .ZN(new_n205));
  INV_X1    g004(.A(G71gat), .ZN(new_n206));
  INV_X1    g005(.A(G78gat), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n206), .B(new_n207), .C1(KEYINPUT88), .C2(KEYINPUT9), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n204), .B1(new_n205), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT9), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT88), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n206), .A2(new_n207), .A3(KEYINPUT87), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT87), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n215), .B1(G71gat), .B2(G78gat), .ZN(new_n216));
  AND3_X1   g015(.A1(new_n214), .A2(new_n216), .A3(new_n205), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n211), .A2(new_n202), .A3(new_n203), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT21), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G231gat), .A2(G233gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n222), .B(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n224), .B(G127gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(G15gat), .B(G22gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT16), .ZN(new_n227));
  AOI21_X1  g026(.A(G1gat), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(G22gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G15gat), .ZN(new_n230));
  INV_X1    g029(.A(G15gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G22gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT81), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n230), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G8gat), .ZN(new_n235));
  INV_X1    g034(.A(G8gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n226), .A2(new_n233), .A3(new_n236), .ZN(new_n237));
  AND3_X1   g036(.A1(new_n228), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n228), .B1(new_n235), .B2(new_n237), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(new_n220), .B2(new_n221), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n225), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(G155gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(G183gat), .B(G211gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n243), .B(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  AND2_X1   g048(.A1(G232gat), .A2(G233gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n250), .A2(KEYINPUT41), .ZN(new_n251));
  XNOR2_X1  g050(.A(G134gat), .B(G162gat), .ZN(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  XOR2_X1   g053(.A(G190gat), .B(G218gat), .Z(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G29gat), .ZN(new_n257));
  INV_X1    g056(.A(G36gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT14), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT14), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(G29gat), .B2(G36gat), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G43gat), .B(G50gat), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  AND2_X1   g063(.A1(KEYINPUT80), .A2(G29gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(KEYINPUT80), .A2(G29gat), .ZN(new_n266));
  OAI21_X1  g065(.A(G36gat), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n262), .A2(new_n264), .A3(KEYINPUT15), .A4(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT17), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT82), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n267), .A2(KEYINPUT15), .A3(new_n261), .A4(new_n259), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(new_n263), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT15), .B1(new_n262), .B2(new_n267), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n268), .B(new_n270), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n269), .A2(KEYINPUT82), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT15), .ZN(new_n277));
  OR2_X1    g076(.A1(KEYINPUT80), .A2(G29gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(KEYINPUT80), .A2(G29gat), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n258), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n259), .A2(new_n261), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n277), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n282), .A2(new_n271), .A3(new_n263), .ZN(new_n283));
  INV_X1    g082(.A(new_n275), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n283), .A2(new_n268), .A3(new_n270), .A4(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n276), .A2(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(G99gat), .B(G106gat), .Z(new_n287));
  NAND2_X1  g086(.A1(G85gat), .A2(G92gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT89), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT90), .ZN(new_n291));
  NAND3_X1  g090(.A1(KEYINPUT89), .A2(G85gat), .A3(G92gat), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT7), .A4(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G99gat), .ZN(new_n294));
  INV_X1    g093(.A(G106gat), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT8), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G85gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT91), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT91), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(G85gat), .ZN(new_n300));
  INV_X1    g099(.A(G92gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n298), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n293), .A2(new_n296), .A3(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT90), .B1(new_n288), .B2(KEYINPUT7), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT7), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n305), .B1(new_n288), .B2(new_n289), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n304), .B1(new_n292), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n287), .B1(new_n303), .B2(new_n307), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n302), .A2(new_n296), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n290), .A2(KEYINPUT7), .A3(new_n292), .ZN(new_n310));
  INV_X1    g109(.A(new_n304), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n287), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n309), .A2(new_n312), .A3(new_n313), .A4(new_n293), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n308), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT92), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n308), .A2(new_n314), .A3(KEYINPUT92), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(KEYINPUT93), .B1(new_n286), .B2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n286), .A2(new_n319), .A3(KEYINPUT93), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n283), .A2(new_n268), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n317), .A2(new_n324), .A3(new_n318), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n250), .A2(KEYINPUT41), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n256), .B1(new_n323), .B2(new_n328), .ZN(new_n329));
  AOI211_X1 g128(.A(new_n255), .B(new_n327), .C1(new_n321), .C2(new_n322), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n254), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n323), .A2(new_n256), .A3(new_n328), .ZN(new_n332));
  INV_X1    g131(.A(new_n322), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n328), .B1(new_n333), .B2(new_n320), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n255), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n332), .A2(new_n335), .A3(new_n253), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n249), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G230gat), .A2(G233gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n315), .A2(new_n220), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT10), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n209), .A2(new_n212), .B1(new_n217), .B2(new_n218), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n308), .A2(new_n343), .A3(new_n314), .ZN(new_n344));
  AND3_X1   g143(.A1(new_n341), .A2(new_n342), .A3(new_n344), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n308), .A2(new_n314), .A3(KEYINPUT92), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT92), .B1(new_n308), .B2(new_n314), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n343), .A2(KEYINPUT10), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n340), .B1(new_n345), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n341), .A2(new_n344), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n351), .A2(G230gat), .A3(G233gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(G120gat), .B(G148gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(G176gat), .B(G204gat), .ZN(new_n354));
  XOR2_X1   g153(.A(new_n353), .B(new_n354), .Z(new_n355));
  NAND3_X1  g154(.A1(new_n350), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT94), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n342), .A3(new_n344), .ZN(new_n359));
  INV_X1    g158(.A(new_n348), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n317), .A2(new_n318), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n358), .B1(new_n362), .B2(new_n340), .ZN(new_n363));
  INV_X1    g162(.A(new_n340), .ZN(new_n364));
  AOI211_X1 g163(.A(KEYINPUT94), .B(new_n364), .C1(new_n359), .C2(new_n361), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n352), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n355), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n357), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n339), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(KEYINPUT95), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT36), .ZN(new_n371));
  XNOR2_X1  g170(.A(G127gat), .B(G134gat), .ZN(new_n372));
  INV_X1    g171(.A(G113gat), .ZN(new_n373));
  INV_X1    g172(.A(G120gat), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT1), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G113gat), .A2(G120gat), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n372), .A2(KEYINPUT68), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  XOR2_X1   g176(.A(G127gat), .B(G134gat), .Z(new_n378));
  INV_X1    g177(.A(KEYINPUT68), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(new_n377), .B(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT24), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n382), .A2(G183gat), .A3(G190gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(G183gat), .B(G190gat), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n383), .B1(new_n384), .B2(new_n382), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n385), .B(KEYINPUT66), .ZN(new_n386));
  NOR2_X1   g185(.A1(G169gat), .A2(G176gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT65), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT23), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n387), .ZN(new_n391));
  NAND2_X1  g190(.A1(G169gat), .A2(G176gat), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n391), .B1(new_n393), .B2(new_n389), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n386), .A2(KEYINPUT25), .A3(new_n390), .A4(new_n394), .ZN(new_n395));
  XOR2_X1   g194(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n396));
  NAND2_X1  g195(.A1(new_n387), .A2(KEYINPUT23), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n394), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n396), .B1(new_n398), .B2(new_n385), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT27), .B(G183gat), .ZN(new_n401));
  INV_X1    g200(.A(G190gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AND2_X1   g202(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n404));
  NOR2_X1   g203(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n405));
  OR3_X1    g204(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n393), .B1(new_n391), .B2(KEYINPUT26), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n407), .B1(new_n388), .B2(KEYINPUT26), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n403), .A2(new_n404), .B1(G183gat), .B2(G190gat), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n406), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n400), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT69), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n410), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n414), .B1(new_n395), .B2(new_n399), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT69), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n381), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n381), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n411), .B2(new_n412), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(G227gat), .A2(G233gat), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT32), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT33), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n423), .B1(new_n420), .B2(new_n421), .ZN(new_n424));
  XOR2_X1   g223(.A(G15gat), .B(G43gat), .Z(new_n425));
  XNOR2_X1  g224(.A(G71gat), .B(G99gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n422), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n427), .ZN(new_n429));
  OAI221_X1 g228(.A(KEYINPUT32), .B1(new_n423), .B2(new_n429), .C1(new_n420), .C2(new_n421), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n428), .A2(KEYINPUT72), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT72), .B1(new_n428), .B2(new_n430), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n420), .A2(KEYINPUT70), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT70), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n434), .B1(new_n417), .B2(new_n419), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(new_n421), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT34), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT34), .B1(G227gat), .B2(G233gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n420), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT71), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT71), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n420), .A2(new_n441), .A3(new_n438), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n437), .A2(new_n443), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n431), .A2(new_n432), .A3(new_n444), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n436), .A2(KEYINPUT34), .B1(new_n440), .B2(new_n442), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n428), .A2(new_n430), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT72), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n371), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n432), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n428), .A2(KEYINPUT72), .A3(new_n430), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n452), .A3(new_n446), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n431), .B1(new_n432), .B2(new_n444), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(new_n454), .A3(KEYINPUT36), .ZN(new_n455));
  XNOR2_X1  g254(.A(G8gat), .B(G36gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(G64gat), .B(G92gat), .ZN(new_n457));
  XOR2_X1   g256(.A(new_n456), .B(new_n457), .Z(new_n458));
  INV_X1    g257(.A(G226gat), .ZN(new_n459));
  INV_X1    g258(.A(G233gat), .ZN(new_n460));
  OAI22_X1  g259(.A1(new_n415), .A2(KEYINPUT29), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NOR3_X1   g261(.A1(new_n415), .A2(new_n459), .A3(new_n460), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT75), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n459), .A2(new_n460), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n411), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT75), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n462), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(G197gat), .ZN(new_n470));
  INV_X1    g269(.A(G204gat), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(G197gat), .A2(G204gat), .ZN(new_n473));
  AND2_X1   g272(.A1(G211gat), .A2(G218gat), .ZN(new_n474));
  OAI22_X1  g273(.A1(new_n472), .A2(new_n473), .B1(KEYINPUT22), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n475), .A2(KEYINPUT73), .ZN(new_n476));
  XNOR2_X1  g275(.A(G211gat), .B(G218gat), .ZN(new_n477));
  OR2_X1    g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n477), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n461), .A2(new_n466), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(KEYINPUT74), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT74), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n469), .A2(new_n481), .B1(new_n482), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT37), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n458), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI22_X1  g288(.A1(new_n469), .A2(new_n481), .B1(new_n482), .B2(new_n486), .ZN(new_n490));
  AOI21_X1  g289(.A(KEYINPUT38), .B1(new_n490), .B2(KEYINPUT37), .ZN(new_n491));
  AOI22_X1  g290(.A1(new_n489), .A2(new_n491), .B1(new_n487), .B2(new_n458), .ZN(new_n492));
  XNOR2_X1  g291(.A(G1gat), .B(G29gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(KEYINPUT0), .ZN(new_n494));
  XNOR2_X1  g293(.A(G57gat), .B(G85gat), .ZN(new_n495));
  XOR2_X1   g294(.A(new_n494), .B(new_n495), .Z(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT76), .ZN(new_n498));
  XOR2_X1   g297(.A(G141gat), .B(G148gat), .Z(new_n499));
  INV_X1    g298(.A(G155gat), .ZN(new_n500));
  INV_X1    g299(.A(G162gat), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT2), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G155gat), .B(G162gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n381), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT4), .ZN(new_n507));
  XOR2_X1   g306(.A(new_n503), .B(new_n504), .Z(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT3), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT3), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n509), .A2(new_n418), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(G225gat), .A2(G233gat), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n507), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  OR2_X1    g313(.A1(new_n514), .A2(KEYINPUT5), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n381), .B(new_n505), .ZN(new_n516));
  INV_X1    g315(.A(new_n513), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n514), .A2(KEYINPUT5), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n498), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n498), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  OAI211_X1 g321(.A(KEYINPUT6), .B(new_n497), .C1(new_n520), .C2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n458), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n463), .A2(KEYINPUT75), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n466), .A2(new_n467), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n461), .B(new_n481), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n482), .A2(new_n486), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n524), .B1(new_n529), .B2(KEYINPUT37), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n487), .A2(new_n488), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT38), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AND2_X1   g331(.A1(new_n515), .A2(new_n519), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n496), .B(new_n521), .C1(new_n533), .C2(new_n498), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT6), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n497), .B1(new_n520), .B2(new_n522), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n492), .A2(new_n523), .A3(new_n532), .A4(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT29), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n511), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n475), .A2(new_n477), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(new_n539), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n475), .A2(new_n477), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n510), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n508), .A2(new_n544), .ZN(new_n545));
  AOI22_X1  g344(.A1(new_n540), .A2(new_n480), .B1(new_n545), .B2(KEYINPUT78), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n545), .A2(KEYINPUT78), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(G228gat), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n548), .B1(new_n549), .B2(new_n460), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n483), .A2(new_n485), .A3(new_n540), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n510), .B1(new_n480), .B2(KEYINPUT29), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n508), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n551), .A2(G228gat), .A3(new_n553), .A4(G233gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(G22gat), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n550), .A2(new_n554), .A3(new_n229), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT77), .ZN(new_n559));
  OAI21_X1  g358(.A(G78gat), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n559), .B1(new_n556), .B2(new_n557), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n561), .A2(new_n207), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT31), .B(G50gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(new_n295), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n560), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n564), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n561), .A2(new_n207), .ZN(new_n567));
  AOI211_X1 g366(.A(new_n559), .B(G78gat), .C1(new_n556), .C2(new_n557), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n487), .A2(new_n458), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n529), .A2(new_n524), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT30), .ZN(new_n573));
  OR3_X1    g372(.A1(new_n529), .A2(KEYINPUT30), .A3(new_n524), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n513), .B1(new_n507), .B2(new_n512), .ZN(new_n575));
  XNOR2_X1  g374(.A(KEYINPUT79), .B(KEYINPUT39), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n497), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(KEYINPUT39), .B1(new_n516), .B2(new_n517), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n577), .B1(new_n575), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n579), .B(KEYINPUT40), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n573), .A2(new_n574), .A3(new_n536), .A4(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n538), .A2(new_n570), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n537), .A2(new_n523), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n573), .A2(new_n574), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(new_n565), .A3(new_n569), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n450), .A2(new_n455), .A3(new_n582), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n453), .A2(new_n454), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n537), .A2(new_n523), .B1(new_n573), .B2(new_n574), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n588), .A2(KEYINPUT35), .A3(new_n589), .A4(new_n570), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n589), .B(new_n570), .C1(new_n445), .C2(new_n449), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT35), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n587), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT86), .ZN(new_n595));
  AOI211_X1 g394(.A(KEYINPUT82), .B(new_n269), .C1(new_n283), .C2(new_n268), .ZN(new_n596));
  AND4_X1   g395(.A1(new_n283), .A2(new_n268), .A3(new_n270), .A4(new_n284), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n241), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(G229gat), .A2(G233gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n240), .A2(new_n324), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n598), .A2(KEYINPUT18), .A3(new_n599), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT83), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n240), .A2(new_n324), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n603), .B1(new_n286), .B2(new_n241), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT83), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n604), .A2(new_n605), .A3(KEYINPUT18), .A4(new_n599), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n602), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n599), .B(KEYINPUT13), .Z(new_n608));
  OAI21_X1  g407(.A(KEYINPUT84), .B1(new_n240), .B2(new_n324), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(new_n600), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT18), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n608), .A2(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G113gat), .B(G141gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G197gat), .ZN(new_n616));
  XOR2_X1   g415(.A(KEYINPUT11), .B(G169gat), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n614), .A2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n607), .A2(new_n613), .A3(new_n619), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(new_n623), .B(KEYINPUT85), .Z(new_n624));
  AND3_X1   g423(.A1(new_n594), .A2(new_n595), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n595), .B1(new_n594), .B2(new_n624), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n370), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT96), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT96), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n629), .B(new_n370), .C1(new_n625), .C2(new_n626), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n583), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G1gat), .ZN(G1324gat));
  INV_X1    g433(.A(new_n584), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n236), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT16), .B(G8gat), .ZN(new_n637));
  AOI211_X1 g436(.A(new_n584), .B(new_n637), .C1(new_n628), .C2(new_n630), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT42), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n639), .B1(KEYINPUT42), .B2(new_n638), .ZN(G1325gat));
  AOI21_X1  g439(.A(G15gat), .B1(new_n631), .B2(new_n588), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n450), .A2(new_n455), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n231), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT97), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n641), .B1(new_n631), .B2(new_n644), .ZN(G1326gat));
  INV_X1    g444(.A(KEYINPUT98), .ZN(new_n646));
  INV_X1    g445(.A(new_n570), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n646), .B1(new_n631), .B2(new_n647), .ZN(new_n648));
  AOI211_X1 g447(.A(KEYINPUT98), .B(new_n570), .C1(new_n628), .C2(new_n630), .ZN(new_n649));
  XNOR2_X1  g448(.A(KEYINPUT43), .B(G22gat), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NOR3_X1   g450(.A1(new_n648), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n594), .A2(new_n624), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT86), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n594), .A2(new_n595), .A3(new_n624), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n629), .B1(new_n656), .B2(new_n370), .ZN(new_n657));
  INV_X1    g456(.A(new_n630), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n647), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT98), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n631), .A2(new_n646), .A3(new_n647), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n650), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n652), .A2(new_n662), .ZN(G1327gat));
  NAND2_X1  g462(.A1(new_n248), .A2(new_n368), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(new_n337), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n656), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n667), .A2(new_n632), .A3(new_n278), .A4(new_n279), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT45), .ZN(new_n669));
  INV_X1    g468(.A(new_n337), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n594), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(KEYINPUT99), .A2(KEYINPUT44), .ZN(new_n672));
  OR2_X1    g471(.A1(KEYINPUT99), .A2(KEYINPUT44), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n671), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n671), .A2(new_n673), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n623), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n664), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  OAI22_X1  g478(.A1(new_n679), .A2(new_n583), .B1(new_n266), .B2(new_n265), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n669), .A2(new_n680), .ZN(G1328gat));
  NAND3_X1  g480(.A1(new_n667), .A2(new_n258), .A3(new_n635), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(KEYINPUT46), .ZN(new_n683));
  OAI21_X1  g482(.A(G36gat), .B1(new_n679), .B2(new_n584), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n682), .A2(KEYINPUT46), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(G1329gat));
  OAI21_X1  g485(.A(G43gat), .B1(new_n679), .B2(new_n642), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT47), .ZN(new_n688));
  INV_X1    g487(.A(new_n588), .ZN(new_n689));
  OR3_X1    g488(.A1(new_n666), .A2(G43gat), .A3(new_n689), .ZN(new_n690));
  AND3_X1   g489(.A1(new_n687), .A2(new_n688), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n688), .B1(new_n687), .B2(new_n690), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n691), .A2(new_n692), .ZN(G1330gat));
  INV_X1    g492(.A(KEYINPUT100), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n570), .B1(new_n666), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n656), .A2(KEYINPUT100), .A3(new_n665), .ZN(new_n696));
  AOI21_X1  g495(.A(G50gat), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT48), .ZN(new_n699));
  AND2_X1   g498(.A1(new_n647), .A2(G50gat), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n676), .A2(new_n678), .A3(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n698), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n701), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT48), .B1(new_n697), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(G1331gat));
  NOR3_X1   g504(.A1(new_n338), .A2(new_n623), .A3(new_n368), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n594), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n583), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT101), .B(G57gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1332gat));
  NOR2_X1   g509(.A1(new_n707), .A2(new_n584), .ZN(new_n711));
  NOR2_X1   g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  AND2_X1   g511(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(new_n711), .B2(new_n712), .ZN(G1333gat));
  OAI21_X1  g514(.A(G71gat), .B1(new_n707), .B2(new_n642), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n588), .A2(new_n206), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(new_n707), .B2(new_n717), .ZN(new_n718));
  XOR2_X1   g517(.A(new_n718), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g518(.A1(new_n707), .A2(new_n570), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(new_n207), .ZN(G1335gat));
  NAND2_X1  g520(.A1(new_n248), .A2(new_n677), .ZN(new_n722));
  XOR2_X1   g521(.A(new_n722), .B(KEYINPUT102), .Z(new_n723));
  NAND3_X1  g522(.A1(new_n594), .A2(new_n670), .A3(new_n723), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n724), .B(KEYINPUT51), .Z(new_n725));
  INV_X1    g524(.A(new_n368), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n298), .A2(new_n300), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n727), .A2(new_n632), .A3(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n728), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n723), .A2(new_n726), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n676), .A2(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n732), .B2(new_n583), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n729), .A2(new_n733), .ZN(G1336gat));
  INV_X1    g533(.A(KEYINPUT52), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n635), .B(new_n731), .C1(new_n674), .C2(new_n675), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G92gat), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n735), .B1(new_n737), .B2(KEYINPUT104), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n584), .A2(G92gat), .A3(new_n368), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT103), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n725), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n738), .B(new_n742), .ZN(G1337gat));
  NAND3_X1  g542(.A1(new_n727), .A2(new_n294), .A3(new_n588), .ZN(new_n744));
  OAI21_X1  g543(.A(G99gat), .B1(new_n732), .B2(new_n642), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(G1338gat));
  OAI21_X1  g545(.A(G106gat), .B1(new_n732), .B2(new_n570), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n647), .A2(new_n295), .A3(new_n726), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT105), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT106), .B1(new_n725), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT53), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n747), .A2(new_n753), .A3(new_n750), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(G1339gat));
  NAND3_X1  g554(.A1(new_n339), .A2(new_n677), .A3(new_n368), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n610), .A2(new_n608), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n604), .A2(new_n599), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n618), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n331), .A2(new_n336), .A3(new_n622), .A4(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n359), .A2(new_n361), .A3(new_n364), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n359), .A2(new_n361), .A3(KEYINPUT107), .A4(new_n364), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT54), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n766), .B1(new_n362), .B2(new_n340), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n350), .A2(KEYINPUT94), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n362), .A2(new_n358), .A3(new_n340), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n769), .A2(new_n766), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n768), .A2(new_n771), .A3(new_n367), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n768), .A2(new_n771), .A3(KEYINPUT55), .A4(new_n367), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n356), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n760), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n772), .A2(new_n773), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n623), .A2(new_n778), .A3(new_n356), .A4(new_n775), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT108), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n622), .A2(new_n759), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n781), .B2(new_n368), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n726), .A2(KEYINPUT108), .A3(new_n622), .A4(new_n759), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n779), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n777), .B1(new_n784), .B2(new_n337), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT109), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n248), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AOI211_X1 g586(.A(KEYINPUT109), .B(new_n777), .C1(new_n337), .C2(new_n784), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n756), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT110), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT110), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n791), .B(new_n756), .C1(new_n787), .C2(new_n788), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n689), .A2(new_n647), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n793), .A2(new_n632), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n795), .A2(new_n635), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n623), .A2(new_n373), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT114), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n790), .A2(new_n570), .A3(new_n792), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT111), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n790), .A2(KEYINPUT111), .A3(new_n570), .A4(new_n792), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n632), .A2(new_n584), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n689), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT112), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n804), .A2(KEYINPUT112), .A3(new_n806), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(new_n624), .A3(new_n810), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n811), .A2(KEYINPUT113), .A3(G113gat), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT113), .B1(new_n811), .B2(G113gat), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n799), .B1(new_n812), .B2(new_n813), .ZN(G1340gat));
  AOI21_X1  g613(.A(G120gat), .B1(new_n796), .B2(new_n726), .ZN(new_n815));
  AOI21_X1  g614(.A(KEYINPUT112), .B1(new_n804), .B2(new_n806), .ZN(new_n816));
  INV_X1    g615(.A(new_n806), .ZN(new_n817));
  AOI211_X1 g616(.A(new_n808), .B(new_n817), .C1(new_n802), .C2(new_n803), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n368), .A2(new_n374), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n815), .B1(new_n819), .B2(new_n820), .ZN(G1341gat));
  AND3_X1   g620(.A1(new_n796), .A2(KEYINPUT115), .A3(new_n249), .ZN(new_n822));
  AOI21_X1  g621(.A(KEYINPUT115), .B1(new_n796), .B2(new_n249), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n822), .A2(new_n823), .A3(G127gat), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n249), .A2(G127gat), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n824), .B1(new_n819), .B2(new_n825), .ZN(G1342gat));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n827));
  INV_X1    g626(.A(G134gat), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n828), .B1(new_n819), .B2(new_n670), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n584), .A2(new_n670), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n795), .A2(G134gat), .A3(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT56), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n831), .B(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n827), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n831), .B(KEYINPUT56), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n816), .A2(new_n818), .A3(new_n337), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n835), .B(KEYINPUT116), .C1(new_n828), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n834), .A2(new_n837), .ZN(G1343gat));
  INV_X1    g637(.A(G141gat), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n781), .A2(new_n368), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT117), .ZN(new_n841));
  INV_X1    g640(.A(new_n776), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT55), .B1(new_n772), .B2(KEYINPUT118), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n843), .B1(KEYINPUT118), .B2(new_n772), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n844), .A2(KEYINPUT119), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(KEYINPUT119), .ZN(new_n846));
  OAI211_X1 g645(.A(KEYINPUT120), .B(new_n842), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n624), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n844), .B(KEYINPUT119), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT120), .B1(new_n849), .B2(new_n842), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n841), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n777), .B1(new_n851), .B2(new_n337), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n756), .B1(new_n852), .B2(new_n249), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n647), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT57), .ZN(new_n855));
  INV_X1    g654(.A(new_n642), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n805), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n793), .A2(new_n858), .A3(new_n647), .ZN(new_n859));
  AND3_X1   g658(.A1(new_n855), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n839), .B1(new_n860), .B2(new_n624), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n642), .A2(new_n647), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT121), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(new_n632), .A3(new_n793), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n624), .A2(new_n839), .ZN(new_n865));
  XNOR2_X1  g664(.A(new_n865), .B(KEYINPUT122), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n864), .A2(new_n635), .A3(new_n866), .ZN(new_n867));
  XOR2_X1   g666(.A(KEYINPUT123), .B(KEYINPUT58), .Z(new_n868));
  OR2_X1    g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n855), .A2(new_n623), .A3(new_n859), .A4(new_n857), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n867), .B1(new_n870), .B2(G141gat), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  OAI22_X1  g671(.A1(new_n861), .A2(new_n869), .B1(new_n871), .B2(new_n872), .ZN(G1344gat));
  OR4_X1    g672(.A1(G148gat), .A2(new_n864), .A3(new_n635), .A4(new_n368), .ZN(new_n874));
  INV_X1    g673(.A(G148gat), .ZN(new_n875));
  AOI211_X1 g674(.A(KEYINPUT59), .B(new_n875), .C1(new_n860), .C2(new_n726), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n852), .A2(new_n249), .ZN(new_n878));
  INV_X1    g677(.A(new_n624), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n370), .A2(new_n879), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n858), .B(new_n647), .C1(new_n878), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n793), .A2(new_n647), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(KEYINPUT57), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n726), .A3(new_n857), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n877), .B1(new_n886), .B2(G148gat), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n874), .B1(new_n876), .B2(new_n887), .ZN(G1345gat));
  NOR3_X1   g687(.A1(new_n864), .A2(new_n635), .A3(new_n248), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n889), .A2(KEYINPUT124), .ZN(new_n890));
  AOI21_X1  g689(.A(G155gat), .B1(new_n889), .B2(KEYINPUT124), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n248), .A2(new_n500), .ZN(new_n892));
  AOI22_X1  g691(.A1(new_n890), .A2(new_n891), .B1(new_n860), .B2(new_n892), .ZN(G1346gat));
  OR3_X1    g692(.A1(new_n864), .A2(G162gat), .A3(new_n830), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n860), .A2(new_n670), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n895), .B2(new_n501), .ZN(G1347gat));
  NAND2_X1  g695(.A1(new_n793), .A2(new_n583), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n689), .A2(new_n584), .A3(new_n647), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g700(.A(G169gat), .B1(new_n901), .B2(new_n623), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n632), .A2(new_n584), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  AOI211_X1 g703(.A(new_n689), .B(new_n904), .C1(new_n802), .C2(new_n803), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n624), .A2(G169gat), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(G1348gat));
  INV_X1    g706(.A(G176gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n901), .A2(new_n908), .A3(new_n726), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n905), .A2(new_n726), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n908), .ZN(G1349gat));
  NAND2_X1  g710(.A1(new_n905), .A2(new_n249), .ZN(new_n912));
  INV_X1    g711(.A(new_n401), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n248), .A2(new_n913), .ZN(new_n914));
  AOI22_X1  g713(.A1(new_n912), .A2(G183gat), .B1(new_n901), .B2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT60), .ZN(new_n916));
  XNOR2_X1  g715(.A(new_n915), .B(new_n916), .ZN(G1350gat));
  NAND3_X1  g716(.A1(new_n901), .A2(new_n402), .A3(new_n670), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n402), .B1(new_n905), .B2(new_n670), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(G1351gat));
  INV_X1    g722(.A(KEYINPUT125), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n884), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n881), .A2(new_n883), .A3(KEYINPUT125), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n856), .A2(new_n904), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n928), .A2(new_n470), .A3(new_n879), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n897), .A2(new_n584), .A3(new_n862), .ZN(new_n930));
  AOI21_X1  g729(.A(G197gat), .B1(new_n930), .B2(new_n623), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n929), .A2(new_n931), .ZN(G1352gat));
  OAI21_X1  g731(.A(G204gat), .B1(new_n928), .B2(new_n368), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n930), .A2(new_n471), .A3(new_n726), .ZN(new_n934));
  XOR2_X1   g733(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n935));
  XNOR2_X1  g734(.A(new_n934), .B(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n933), .A2(new_n936), .ZN(G1353gat));
  INV_X1    g736(.A(G211gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n930), .A2(new_n938), .A3(new_n249), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n885), .A2(new_n249), .A3(new_n927), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n940), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT63), .B1(new_n940), .B2(G211gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(G1354gat));
  AOI21_X1  g742(.A(G218gat), .B1(new_n930), .B2(new_n670), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n670), .A2(G218gat), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n945), .B1(new_n928), .B2(new_n946), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n925), .A2(KEYINPUT127), .A3(new_n926), .A4(new_n927), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(G1355gat));
endmodule


