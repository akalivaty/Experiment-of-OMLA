//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(G110), .B(G140), .ZN(new_n192));
  INV_X1    g006(.A(G227), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n193), .A2(G953), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n192), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  AND2_X1   g013(.A1(KEYINPUT0), .A2(G128), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n197), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT64), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(G143), .B(G146), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT64), .A3(new_n200), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n197), .A2(new_n199), .ZN(new_n206));
  NOR2_X1   g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n200), .A2(new_n207), .ZN(new_n208));
  AOI22_X1  g022(.A1(new_n203), .A2(new_n205), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(new_n210), .B2(G107), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(G104), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n210), .A2(G107), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n211), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G101), .ZN(new_n217));
  AND2_X1   g031(.A1(KEYINPUT75), .A2(G101), .ZN(new_n218));
  NOR2_X1   g032(.A1(KEYINPUT75), .A2(G101), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n220), .A2(new_n211), .A3(new_n214), .A4(new_n215), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n217), .A2(KEYINPUT4), .A3(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n209), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT76), .B(KEYINPUT4), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n216), .A2(G101), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT77), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT77), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n216), .A2(new_n227), .A3(G101), .A4(new_n224), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G101), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n213), .A2(G104), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(new_n215), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n211), .A2(new_n214), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  OR2_X1    g048(.A1(KEYINPUT75), .A2(G101), .ZN(new_n235));
  NAND2_X1  g049(.A1(KEYINPUT75), .A2(G101), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(new_n215), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n232), .B1(new_n234), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G128), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n241), .B1(G143), .B2(new_n196), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT78), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT1), .B1(new_n198), .B2(G146), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT78), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n204), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  AND4_X1   g061(.A1(new_n241), .A2(new_n197), .A3(new_n199), .A4(G128), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n239), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT10), .ZN(new_n250));
  AOI22_X1  g064(.A1(new_n223), .A2(new_n229), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT11), .ZN(new_n252));
  INV_X1    g066(.A(G134), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(G137), .ZN(new_n254));
  INV_X1    g068(.A(G137), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(KEYINPUT11), .A3(G134), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n253), .A2(G137), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n254), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G131), .ZN(new_n259));
  INV_X1    g073(.A(G131), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n254), .A2(new_n256), .A3(new_n260), .A4(new_n257), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT80), .ZN(new_n263));
  INV_X1    g077(.A(new_n232), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n221), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT79), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n221), .A2(new_n264), .A3(KEYINPUT79), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n245), .A2(G128), .B1(new_n197), .B2(new_n199), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT10), .B1(new_n248), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n263), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  AOI211_X1 g087(.A(KEYINPUT80), .B(new_n271), .C1(new_n267), .C2(new_n268), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n251), .B(new_n262), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n206), .B1(new_n242), .B2(new_n240), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n204), .A2(new_n241), .A3(G128), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n267), .A2(new_n280), .A3(new_n268), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n249), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n259), .A2(new_n261), .ZN(new_n283));
  AOI21_X1  g097(.A(KEYINPUT12), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT12), .ZN(new_n285));
  AOI211_X1 g099(.A(new_n285), .B(new_n262), .C1(new_n281), .C2(new_n249), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n195), .B1(new_n276), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT81), .ZN(new_n289));
  INV_X1    g103(.A(new_n195), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n275), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n251), .B1(new_n273), .B2(new_n274), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n283), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n289), .B1(new_n275), .B2(new_n290), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n288), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT82), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n288), .B(KEYINPUT82), .C1(new_n294), .C2(new_n295), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(G469), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G469), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n275), .B(new_n290), .C1(new_n286), .C2(new_n284), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n290), .B1(new_n293), .B2(new_n275), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n301), .B(new_n190), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(G469), .A2(G902), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n191), .B1(new_n300), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G210), .B1(G237), .B2(G902), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(G110), .B(G122), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT2), .B(G113), .Z(new_n313));
  XNOR2_X1  g127(.A(G116), .B(G119), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT2), .B(G113), .ZN(new_n316));
  INV_X1    g130(.A(G119), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G116), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n317), .A2(G116), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n316), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n315), .A2(new_n321), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n216), .A2(G101), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT4), .B1(new_n233), .B2(new_n237), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(new_n228), .B2(new_n226), .ZN(new_n326));
  INV_X1    g140(.A(G113), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT5), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n327), .B1(new_n319), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n314), .A2(KEYINPUT5), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n315), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n332), .B1(new_n267), .B2(new_n268), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n312), .B1(new_n326), .B2(new_n333), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n329), .A2(new_n330), .B1(new_n314), .B2(new_n313), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n269), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n229), .A2(new_n322), .A3(new_n222), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(new_n311), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n334), .A2(KEYINPUT6), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT6), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n340), .B(new_n312), .C1(new_n326), .C2(new_n333), .ZN(new_n341));
  INV_X1    g155(.A(G125), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n277), .A2(new_n278), .A3(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n343), .B1(new_n209), .B2(new_n342), .ZN(new_n344));
  INV_X1    g158(.A(G224), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(G953), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n344), .B(new_n346), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n339), .A2(new_n341), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(KEYINPUT7), .B1(new_n345), .B2(G953), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT84), .B1(new_n344), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n349), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n343), .B(new_n351), .C1(new_n209), .C2(new_n342), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n311), .B(KEYINPUT8), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT83), .B1(new_n335), .B2(new_n239), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT83), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n332), .A2(new_n357), .A3(new_n265), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n355), .B1(new_n359), .B2(new_n333), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n344), .A2(KEYINPUT84), .A3(new_n349), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n354), .A2(new_n360), .A3(new_n338), .A4(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n190), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n310), .B1(new_n348), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n339), .A2(new_n341), .A3(new_n347), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n365), .A2(new_n190), .A3(new_n362), .A4(new_n309), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(G214), .B1(G237), .B2(G902), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(G475), .A2(G902), .ZN(new_n370));
  XNOR2_X1  g184(.A(G113), .B(G122), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n371), .B(new_n210), .ZN(new_n372));
  INV_X1    g186(.A(G140), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G125), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n342), .A2(G140), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT71), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT19), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT71), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n376), .A2(KEYINPUT19), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n196), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT86), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT86), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n381), .A2(new_n385), .A3(new_n196), .A4(new_n382), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT69), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n374), .A2(new_n375), .A3(new_n387), .A4(KEYINPUT16), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT16), .ZN(new_n389));
  OAI21_X1  g203(.A(KEYINPUT69), .B1(new_n374), .B2(KEYINPUT16), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(G237), .A2(G953), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(G143), .A3(G214), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(G143), .B1(new_n392), .B2(G214), .ZN(new_n395));
  OAI21_X1  g209(.A(G131), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n392), .A2(G214), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n198), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(new_n260), .A3(new_n393), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n391), .A2(G146), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n384), .A2(new_n386), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n378), .A2(new_n196), .A3(new_n380), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n376), .A2(G146), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n394), .A2(new_n395), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n405), .A2(KEYINPUT85), .B1(KEYINPUT18), .B2(G131), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n398), .A2(new_n393), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT85), .ZN(new_n408));
  NAND2_X1  g222(.A1(KEYINPUT18), .A2(G131), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n404), .B1(new_n406), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n372), .B1(new_n401), .B2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT17), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n396), .A2(new_n413), .A3(new_n399), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n391), .A2(G146), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n196), .B(new_n388), .C1(new_n389), .C2(new_n390), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n407), .A2(KEYINPUT17), .A3(G131), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n414), .A2(new_n415), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n418), .A2(new_n411), .A3(new_n372), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n370), .B1(new_n412), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT20), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n422), .B(new_n370), .C1(new_n412), .C2(new_n419), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n372), .B1(new_n418), .B2(new_n411), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n190), .B1(new_n419), .B2(new_n424), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n421), .A2(new_n423), .B1(G475), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n198), .A2(G128), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n240), .A2(G143), .ZN(new_n428));
  AND3_X1   g242(.A1(new_n427), .A2(new_n428), .A3(new_n253), .ZN(new_n429));
  INV_X1    g243(.A(G122), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G116), .ZN(new_n431));
  INV_X1    g245(.A(G116), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G122), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G107), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n431), .A2(new_n433), .A3(new_n213), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n429), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT13), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n427), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n198), .A2(KEYINPUT13), .A3(G128), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n439), .A2(new_n440), .A3(new_n428), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n437), .B1(new_n253), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n432), .A2(KEYINPUT14), .A3(G122), .ZN(new_n443));
  OAI211_X1 g257(.A(G107), .B(new_n443), .C1(new_n434), .C2(KEYINPUT14), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n253), .B1(new_n427), .B2(new_n428), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n444), .B(new_n436), .C1(new_n429), .C2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G217), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n188), .A2(new_n448), .A3(G953), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n442), .A2(new_n446), .A3(new_n449), .ZN(new_n452));
  AOI21_X1  g266(.A(G902), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G478), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n453), .B1(KEYINPUT15), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n452), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n449), .B1(new_n442), .B2(new_n446), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n190), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n454), .A2(KEYINPUT15), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n455), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G952), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(G953), .ZN(new_n464));
  NAND2_X1  g278(.A1(G234), .A2(G237), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(KEYINPUT87), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT21), .B(G898), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n465), .A2(G902), .A3(G953), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n468), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n426), .A2(new_n462), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n369), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n308), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n253), .A2(G137), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n255), .A2(G134), .ZN(new_n478));
  OAI21_X1  g292(.A(G131), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n261), .B(new_n479), .C1(new_n248), .C2(new_n270), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n206), .A2(new_n208), .ZN(new_n481));
  AOI21_X1  g295(.A(KEYINPUT64), .B1(new_n204), .B2(new_n200), .ZN(new_n482));
  AND4_X1   g296(.A1(KEYINPUT64), .A2(new_n197), .A3(new_n199), .A4(new_n200), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n480), .B1(new_n262), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n322), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n261), .A2(new_n479), .ZN(new_n487));
  AOI22_X1  g301(.A1(new_n209), .A2(new_n283), .B1(new_n487), .B2(new_n279), .ZN(new_n488));
  INV_X1    g302(.A(new_n322), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT28), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT29), .ZN(new_n493));
  AOI21_X1  g307(.A(KEYINPUT28), .B1(new_n488), .B2(new_n489), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n392), .A2(G210), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n496), .B(KEYINPUT27), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT26), .B(G101), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n497), .B(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT65), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n499), .B(new_n500), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n492), .A2(new_n493), .A3(new_n495), .A4(new_n501), .ZN(new_n502));
  XOR2_X1   g316(.A(new_n497), .B(new_n498), .Z(new_n503));
  NAND2_X1  g317(.A1(new_n485), .A2(KEYINPUT30), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n209), .A2(new_n283), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT30), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n506), .A3(new_n480), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n489), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n490), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n503), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n502), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT28), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(new_n486), .B2(new_n490), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(new_n494), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n493), .B1(new_n514), .B2(new_n499), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n190), .B1(new_n511), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G472), .ZN(new_n517));
  NOR2_X1   g331(.A1(G472), .A2(G902), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n499), .B(KEYINPUT65), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n513), .B2(new_n494), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n490), .A2(new_n499), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT31), .B1(new_n508), .B2(new_n522), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n505), .A2(new_n506), .A3(new_n480), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n506), .B1(new_n505), .B2(new_n480), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n322), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT31), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n503), .B1(new_n488), .B2(new_n489), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n521), .A2(new_n523), .A3(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT66), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n521), .A2(new_n523), .A3(new_n529), .A4(KEYINPUT66), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n519), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n517), .B1(new_n534), .B2(KEYINPUT32), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT67), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n532), .A2(new_n533), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT32), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n519), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n536), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n539), .ZN(new_n541));
  AOI211_X1 g355(.A(KEYINPUT67), .B(new_n541), .C1(new_n532), .C2(new_n533), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n535), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT22), .B(G137), .ZN(new_n544));
  INV_X1    g358(.A(G953), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n545), .A2(G221), .A3(G234), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n544), .B(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(G110), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n240), .B(G119), .C1(KEYINPUT68), .C2(KEYINPUT23), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT23), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n551), .B1(new_n317), .B2(G128), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT68), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n553), .B1(new_n317), .B2(G128), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n549), .B(new_n550), .C1(new_n552), .C2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n240), .A2(G119), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n317), .A2(G128), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT24), .B(G110), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n555), .A2(KEYINPUT70), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT70), .B1(new_n555), .B2(new_n560), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n415), .B(new_n402), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n558), .A2(new_n559), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n550), .B1(new_n552), .B2(new_n554), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n564), .B1(G110), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n416), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT16), .ZN(new_n568));
  OR3_X1    g382(.A1(new_n342), .A2(KEYINPUT16), .A3(G140), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT69), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n196), .B1(new_n570), .B2(new_n388), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n566), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT72), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n563), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n573), .B1(new_n563), .B2(new_n572), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n548), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n563), .A2(new_n572), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n547), .B1(new_n577), .B2(KEYINPUT72), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n448), .B1(G234), .B2(new_n190), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n579), .A2(G902), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n576), .A2(new_n190), .A3(new_n578), .ZN(new_n582));
  NOR2_X1   g396(.A1(KEYINPUT73), .A2(KEYINPUT25), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n583), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n576), .A2(new_n190), .A3(new_n585), .A4(new_n578), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n581), .B1(new_n587), .B2(new_n580), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n543), .A2(KEYINPUT74), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT74), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n537), .A2(new_n518), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n538), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n537), .A2(new_n539), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT67), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n537), .A2(new_n536), .A3(new_n539), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n593), .A2(new_n595), .A3(new_n517), .A4(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n591), .B1(new_n597), .B2(new_n588), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n476), .B1(new_n590), .B2(new_n598), .ZN(new_n599));
  XOR2_X1   g413(.A(new_n599), .B(new_n220), .Z(G3));
  INV_X1    g414(.A(G472), .ZN(new_n601));
  AOI21_X1  g415(.A(G902), .B1(new_n532), .B2(new_n533), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n592), .B(new_n588), .C1(new_n601), .C2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n368), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n605), .B1(new_n364), .B2(new_n366), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT88), .B1(new_n453), .B2(G478), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT88), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n458), .A2(new_n608), .A3(new_n454), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT33), .B1(new_n456), .B2(new_n457), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n451), .A2(new_n611), .A3(new_n452), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n454), .A2(G902), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n607), .A2(new_n609), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n421), .A2(new_n423), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n425), .A2(G475), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n615), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n606), .A2(new_n473), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n604), .A2(new_n308), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT34), .B(G104), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  NAND2_X1  g437(.A1(new_n426), .A2(new_n461), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n625), .A2(new_n606), .A3(new_n473), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n604), .A2(new_n308), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT35), .B(G107), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT89), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n627), .B(new_n629), .ZN(G9));
  AOI21_X1  g444(.A(new_n601), .B1(new_n537), .B2(new_n190), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n534), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n547), .A2(KEYINPUT36), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n577), .B(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n580), .A2(G902), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT90), .ZN(new_n637));
  INV_X1    g451(.A(new_n580), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n584), .B2(new_n586), .ZN(new_n639));
  OR2_X1    g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n308), .A2(new_n475), .A3(new_n632), .A4(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT37), .B(G110), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G12));
  INV_X1    g457(.A(G900), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n468), .B1(new_n644), .B2(new_n471), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n624), .A2(new_n645), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n640), .A2(new_n606), .A3(new_n646), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n597), .A2(new_n647), .A3(new_n308), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(new_n240), .ZN(G30));
  XOR2_X1   g463(.A(new_n645), .B(KEYINPUT39), .Z(new_n650));
  NAND2_X1  g464(.A1(new_n308), .A2(new_n650), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n651), .A2(KEYINPUT40), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n367), .B(KEYINPUT38), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n637), .A2(new_n639), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n426), .A2(new_n462), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n653), .A2(new_n368), .A3(new_n654), .A4(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n595), .A2(new_n596), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n508), .A2(new_n522), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n658), .B1(new_n491), .B2(new_n520), .ZN(new_n659));
  OAI21_X1  g473(.A(G472), .B1(new_n659), .B2(G902), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n593), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n651), .A2(KEYINPUT40), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n652), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G143), .ZN(G45));
  NAND2_X1  g480(.A1(new_n616), .A2(new_n617), .ZN(new_n667));
  INV_X1    g481(.A(new_n615), .ZN(new_n668));
  INV_X1    g482(.A(new_n645), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n369), .A2(new_n654), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n597), .A2(new_n308), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(KEYINPUT91), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT91), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n597), .A2(new_n671), .A3(new_n674), .A4(new_n308), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  OAI21_X1  g491(.A(new_n190), .B1(new_n303), .B2(new_n304), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(G469), .ZN(new_n679));
  INV_X1    g493(.A(new_n191), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n679), .A2(new_n680), .A3(new_n305), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n619), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n597), .A2(new_n682), .A3(new_n588), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT41), .B(G113), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G15));
  NAND3_X1  g499(.A1(new_n625), .A2(new_n606), .A3(new_n473), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n681), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n597), .A2(new_n687), .A3(new_n588), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT92), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n597), .A2(new_n687), .A3(KEYINPUT92), .A4(new_n588), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G116), .ZN(G18));
  NOR2_X1   g507(.A1(new_n681), .A2(new_n369), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n654), .A2(new_n474), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n597), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  INV_X1    g511(.A(KEYINPUT95), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n698), .B1(new_n602), .B2(new_n601), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n521), .A2(new_n523), .ZN(new_n700));
  AOI22_X1  g514(.A1(new_n700), .A2(KEYINPUT94), .B1(new_n527), .B2(new_n658), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n701), .B1(KEYINPUT94), .B2(new_n700), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n518), .B(KEYINPUT93), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n679), .A2(new_n680), .A3(new_n305), .A4(new_n473), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n606), .A2(new_n655), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n631), .A2(KEYINPUT95), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n705), .A2(new_n708), .A3(new_n588), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  AOI21_X1  g525(.A(KEYINPUT96), .B1(new_n618), .B2(new_n669), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT96), .ZN(new_n713));
  NOR4_X1   g527(.A1(new_n426), .A2(new_n713), .A3(new_n615), .A4(new_n645), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n694), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n709), .A2(new_n640), .A3(new_n699), .A4(new_n704), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT97), .B(G125), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G27));
  AOI21_X1  g534(.A(KEYINPUT99), .B1(new_n537), .B2(new_n539), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT99), .ZN(new_n722));
  AOI211_X1 g536(.A(new_n722), .B(new_n541), .C1(new_n532), .C2(new_n533), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  AOI22_X1  g538(.A1(new_n592), .A2(new_n538), .B1(G472), .B2(new_n516), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n588), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n364), .A2(new_n368), .A3(new_n366), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n288), .B(G469), .C1(new_n294), .C2(new_n295), .ZN(new_n729));
  XOR2_X1   g543(.A(new_n306), .B(KEYINPUT98), .Z(new_n730));
  NAND3_X1  g544(.A1(new_n305), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  AND3_X1   g545(.A1(new_n728), .A2(new_n731), .A3(new_n680), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(KEYINPUT42), .A3(new_n715), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT100), .B1(new_n727), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n670), .A2(new_n713), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n618), .A2(KEYINPUT96), .A3(new_n669), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n728), .A2(new_n731), .A3(new_n680), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT42), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT100), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n589), .B1(new_n724), .B2(new_n725), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n597), .A2(new_n588), .A3(new_n732), .A4(new_n715), .ZN(new_n744));
  AOI22_X1  g558(.A1(new_n734), .A2(new_n743), .B1(new_n739), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n260), .ZN(G33));
  NAND4_X1  g560(.A1(new_n597), .A2(new_n588), .A3(new_n732), .A4(new_n646), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G134), .ZN(G36));
  NAND3_X1  g562(.A1(new_n364), .A2(new_n368), .A3(new_n366), .ZN(new_n749));
  OAI21_X1  g563(.A(KEYINPUT103), .B1(new_n632), .B2(new_n654), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT103), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n640), .B(new_n751), .C1(new_n534), .C2(new_n631), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n426), .A2(new_n668), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT102), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n755), .A2(KEYINPUT43), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(KEYINPUT43), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n754), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n758), .B1(new_n754), .B2(new_n757), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT44), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n749), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n762), .B1(new_n761), .B2(new_n760), .ZN(new_n763));
  INV_X1    g577(.A(new_n730), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n298), .A2(new_n299), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT101), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n296), .A2(new_n766), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n767), .A2(new_n768), .A3(G469), .A4(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(G469), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT45), .B1(new_n298), .B2(new_n299), .ZN(new_n772));
  OAI21_X1  g586(.A(KEYINPUT101), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n764), .B1(new_n770), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n774), .A2(KEYINPUT46), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n305), .B1(new_n774), .B2(KEYINPUT46), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n680), .B(new_n650), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n763), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(new_n255), .ZN(G39));
  OAI21_X1  g593(.A(new_n680), .B1(new_n775), .B2(new_n776), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT47), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(KEYINPUT47), .B(new_n680), .C1(new_n775), .C2(new_n776), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n588), .A2(new_n670), .A3(new_n749), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(new_n543), .A3(new_n785), .ZN(new_n786));
  XOR2_X1   g600(.A(KEYINPUT104), .B(G140), .Z(new_n787));
  XNOR2_X1  g601(.A(new_n786), .B(new_n787), .ZN(G42));
  OR2_X1    g602(.A1(new_n681), .A2(new_n749), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT107), .ZN(new_n790));
  AND2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  NOR3_X1   g606(.A1(new_n791), .A2(new_n792), .A3(new_n467), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n759), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n727), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT48), .ZN(new_n796));
  INV_X1    g610(.A(new_n662), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(new_n589), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n793), .A2(new_n618), .A3(new_n798), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n709), .A2(new_n699), .A3(new_n704), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n588), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n759), .A2(new_n468), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n694), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n799), .A2(new_n464), .A3(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n796), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n679), .A2(new_n305), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n680), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n728), .B(new_n803), .C1(new_n784), .C2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT51), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n793), .A2(new_n426), .A3(new_n615), .A4(new_n798), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n811), .B1(new_n717), .B2(new_n794), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n653), .A2(new_n368), .A3(new_n681), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n803), .A2(new_n813), .ZN(new_n814));
  OR2_X1    g628(.A1(new_n814), .A2(KEYINPUT50), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(KEYINPUT50), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n812), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n809), .A2(new_n810), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n810), .B1(new_n809), .B2(new_n817), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n806), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT108), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT108), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n822), .B(new_n806), .C1(new_n818), .C2(new_n819), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n648), .A2(new_n718), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n707), .A2(new_n640), .A3(new_n645), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n797), .A2(new_n680), .A3(new_n731), .A4(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n676), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(KEYINPUT52), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n676), .A2(new_n824), .A3(new_n829), .A4(new_n826), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n604), .B(new_n308), .C1(new_n620), .C2(new_n626), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n832), .A2(new_n641), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n599), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n745), .A2(new_n834), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n710), .A2(new_n683), .A3(new_n696), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n737), .A2(new_n738), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT105), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n800), .A2(new_n837), .A3(new_n838), .A4(new_n640), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n732), .A2(new_n715), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT105), .B1(new_n840), .B2(new_n717), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n426), .A2(new_n462), .A3(new_n669), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n654), .A2(new_n749), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n597), .A2(new_n308), .A3(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n747), .A2(new_n845), .ZN(new_n846));
  AND4_X1   g660(.A1(new_n692), .A2(new_n836), .A3(new_n842), .A4(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT106), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n835), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n744), .A2(new_n739), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n727), .A2(new_n733), .A3(KEYINPUT100), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n741), .B1(new_n740), .B2(new_n742), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n832), .A2(new_n641), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT74), .B1(new_n543), .B2(new_n589), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n597), .A2(new_n591), .A3(new_n588), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n854), .B1(new_n857), .B2(new_n476), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n853), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n692), .A2(new_n836), .A3(new_n842), .A4(new_n846), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT106), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n831), .B1(new_n849), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n863), .B1(new_n824), .B2(new_n829), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n862), .A2(KEYINPUT53), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT54), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n859), .A2(new_n860), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n824), .A2(new_n829), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n863), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n868), .A2(new_n830), .A3(new_n828), .A4(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n871), .B1(new_n862), .B2(KEYINPUT53), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n872), .A2(KEYINPUT54), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n821), .A2(new_n823), .A3(new_n867), .A4(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n463), .A2(new_n545), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OR4_X1    g690(.A1(new_n589), .A2(new_n754), .A3(new_n191), .A4(new_n605), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n807), .B(KEYINPUT49), .ZN(new_n878));
  OR4_X1    g692(.A1(new_n797), .A2(new_n877), .A3(new_n878), .A4(new_n653), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n876), .A2(new_n879), .ZN(G75));
  NAND3_X1  g694(.A1(new_n872), .A2(G210), .A3(G902), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT56), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n339), .A2(new_n341), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT109), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n347), .B(KEYINPUT55), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n885), .B(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n463), .A2(G953), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT110), .ZN(new_n890));
  INV_X1    g704(.A(new_n887), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n881), .A2(new_n882), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n888), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT111), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n888), .A2(KEYINPUT111), .A3(new_n890), .A4(new_n892), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(G51));
  INV_X1    g711(.A(new_n890), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n872), .B(KEYINPUT54), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n730), .B(KEYINPUT112), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT57), .Z(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n303), .A2(new_n304), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT113), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n872), .A2(G902), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n770), .A3(new_n773), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n898), .B1(new_n905), .B2(new_n907), .ZN(G54));
  NAND3_X1  g722(.A1(new_n906), .A2(KEYINPUT58), .A3(G475), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n412), .A2(new_n419), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n909), .B(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(new_n898), .ZN(G60));
  NAND2_X1  g726(.A1(G478), .A2(G902), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT59), .Z(new_n914));
  AOI21_X1  g728(.A(new_n914), .B1(new_n873), .B2(new_n867), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n890), .B1(new_n915), .B2(new_n613), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT114), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n914), .B1(new_n610), .B2(new_n612), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n899), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n899), .A2(new_n918), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(KEYINPUT114), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n916), .B1(new_n919), .B2(new_n921), .ZN(G63));
  INV_X1    g736(.A(KEYINPUT119), .ZN(new_n923));
  NAND2_X1  g737(.A1(G217), .A2(G902), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT116), .ZN(new_n925));
  XNOR2_X1  g739(.A(KEYINPUT115), .B(KEYINPUT60), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n872), .A2(new_n634), .A3(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n898), .A2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n579), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n931), .B1(new_n872), .B2(new_n927), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n928), .B(new_n930), .C1(new_n932), .C2(KEYINPUT118), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT118), .ZN(new_n934));
  AOI211_X1 g748(.A(new_n934), .B(new_n931), .C1(new_n872), .C2(new_n927), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n923), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n872), .A2(new_n927), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n579), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n934), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n928), .A2(new_n930), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n932), .A2(KEYINPUT118), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n939), .A2(new_n940), .A3(KEYINPUT119), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n936), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT117), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n938), .A2(new_n944), .A3(new_n890), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT117), .B1(new_n932), .B2(new_n898), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n945), .A2(new_n928), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n929), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n943), .A2(new_n948), .ZN(G66));
  INV_X1    g763(.A(new_n469), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n545), .B1(new_n950), .B2(G224), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n858), .A2(new_n692), .A3(new_n836), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n951), .B1(new_n952), .B2(new_n545), .ZN(new_n953));
  INV_X1    g767(.A(G898), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n885), .B1(new_n954), .B2(G953), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n953), .B(new_n955), .ZN(G69));
  NAND2_X1  g770(.A1(new_n504), .A2(new_n507), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n381), .A2(new_n382), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n957), .B(new_n958), .Z(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(G900), .B2(G953), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n853), .A2(new_n676), .A3(new_n747), .A4(new_n824), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n778), .A2(new_n962), .ZN(new_n963));
  OR3_X1    g777(.A1(new_n777), .A2(new_n707), .A3(new_n727), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n786), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n961), .B1(new_n965), .B2(G953), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n665), .A2(new_n676), .A3(new_n824), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n967), .A2(KEYINPUT121), .A3(KEYINPUT62), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(KEYINPUT62), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT121), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT62), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n665), .A2(new_n676), .A3(new_n972), .A4(new_n824), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT120), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n973), .A2(new_n974), .ZN(new_n976));
  AOI22_X1  g790(.A1(new_n968), .A2(new_n971), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT123), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n624), .B1(new_n426), .B2(new_n615), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n749), .B1(new_n979), .B2(KEYINPUT122), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n980), .B1(KEYINPUT122), .B2(new_n979), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n981), .A2(new_n651), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n978), .B1(new_n857), .B2(new_n982), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n857), .A2(new_n978), .A3(new_n982), .ZN(new_n984));
  OAI22_X1  g798(.A1(new_n763), .A2(new_n777), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n977), .A2(new_n786), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n960), .B1(new_n987), .B2(G953), .ZN(new_n988));
  OAI21_X1  g802(.A(G953), .B1(new_n193), .B2(new_n644), .ZN(new_n989));
  OAI211_X1 g803(.A(new_n966), .B(new_n988), .C1(KEYINPUT124), .C2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(KEYINPUT124), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(G72));
  NAND2_X1  g806(.A1(G472), .A2(G902), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT63), .Z(new_n994));
  INV_X1    g808(.A(new_n510), .ZN(new_n995));
  OAI221_X1 g809(.A(new_n994), .B1(new_n658), .B2(new_n995), .C1(new_n865), .C2(new_n866), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n994), .B1(new_n965), .B2(new_n952), .ZN(new_n997));
  NOR3_X1   g811(.A1(new_n508), .A2(new_n509), .A3(new_n499), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n996), .A2(new_n999), .A3(new_n890), .ZN(new_n1000));
  INV_X1    g814(.A(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT125), .ZN(new_n1002));
  INV_X1    g816(.A(new_n952), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n977), .A2(new_n786), .A3(new_n1003), .A4(new_n986), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1002), .B1(new_n1004), .B2(new_n994), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n499), .B1(new_n508), .B2(new_n509), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n1004), .A2(new_n1002), .A3(new_n994), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1001), .A2(new_n1010), .A3(KEYINPUT126), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT126), .ZN(new_n1012));
  NOR3_X1   g826(.A1(new_n1008), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1012), .B1(new_n1013), .B2(new_n1000), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1011), .A2(new_n1014), .ZN(G57));
endmodule


