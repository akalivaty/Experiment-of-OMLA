//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 1 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:31 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n844, new_n845, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965;
  INV_X1    g000(.A(KEYINPUT36), .ZN(new_n202));
  XOR2_X1   g001(.A(G15gat), .B(G43gat), .Z(new_n203));
  XNOR2_X1  g002(.A(G71gat), .B(G99gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G227gat), .A2(G233gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT64), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G169gat), .ZN(new_n209));
  INV_X1    g008(.A(G176gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n214), .A2(KEYINPUT67), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(KEYINPUT67), .ZN(new_n216));
  AND3_X1   g015(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(G183gat), .B(G190gat), .Z(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT24), .ZN(new_n219));
  INV_X1    g018(.A(G183gat), .ZN(new_n220));
  INV_X1    g019(.A(G190gat), .ZN(new_n221));
  OR3_X1    g020(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT24), .ZN(new_n222));
  NOR2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(KEYINPUT23), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n224), .A2(KEYINPUT25), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n217), .A2(new_n219), .A3(new_n222), .A4(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n226), .B(KEYINPUT68), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n224), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n223), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n229), .A2(new_n214), .A3(new_n230), .A4(new_n213), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT66), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n233), .A2(new_n219), .A3(new_n222), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n231), .A2(new_n232), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n227), .B1(new_n236), .B2(KEYINPUT25), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT27), .B(G183gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(KEYINPUT28), .A3(new_n221), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT27), .B1(new_n220), .B2(KEYINPUT69), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n220), .A2(KEYINPUT27), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n221), .B(new_n240), .C1(new_n241), .C2(KEYINPUT69), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n243));
  AND2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT28), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n245), .B1(new_n242), .B2(new_n243), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n239), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n211), .A2(KEYINPUT26), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT26), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n214), .B1(new_n223), .B2(new_n249), .ZN(new_n250));
  OAI221_X1 g049(.A(new_n247), .B1(new_n220), .B2(new_n221), .C1(new_n248), .C2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n237), .A2(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(G127gat), .B(G134gat), .Z(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(KEYINPUT1), .ZN(new_n254));
  INV_X1    g053(.A(G120gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G113gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(KEYINPUT71), .ZN(new_n257));
  INV_X1    g056(.A(G113gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G120gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT72), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n254), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n256), .A2(new_n259), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n253), .B1(new_n262), .B2(KEYINPUT1), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n252), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n237), .A2(new_n264), .A3(new_n251), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n208), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n205), .B1(new_n268), .B2(KEYINPUT33), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT32), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  OR2_X1    g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n269), .A2(new_n271), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n266), .A2(new_n208), .A3(new_n267), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n275), .A2(KEYINPUT73), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n276), .A2(KEYINPUT34), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n275), .A2(KEYINPUT73), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n272), .B(new_n273), .C1(KEYINPUT34), .C2(new_n276), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n279), .B1(new_n278), .B2(new_n280), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n202), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT31), .B(G50gat), .ZN(new_n285));
  INV_X1    g084(.A(G106gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G228gat), .A2(G233gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n289), .B(KEYINPUT82), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT22), .ZN(new_n291));
  INV_X1    g090(.A(G211gat), .ZN(new_n292));
  INV_X1    g091(.A(G218gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT74), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT74), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n296), .B(new_n291), .C1(new_n292), .C2(new_n293), .ZN(new_n297));
  XNOR2_X1  g096(.A(G197gat), .B(G204gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n295), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  XOR2_X1   g098(.A(G211gat), .B(G218gat), .Z(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT29), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT3), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G148gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n304), .A2(G141gat), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n305), .A2(KEYINPUT76), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(KEYINPUT76), .ZN(new_n307));
  INV_X1    g106(.A(G141gat), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT77), .B1(new_n308), .B2(G148gat), .ZN(new_n309));
  OR3_X1    g108(.A1(new_n308), .A2(KEYINPUT77), .A3(G148gat), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n306), .A2(new_n307), .A3(new_n309), .A4(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312));
  INV_X1    g111(.A(G155gat), .ZN(new_n313));
  INV_X1    g112(.A(G162gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n312), .B1(new_n315), .B2(KEYINPUT2), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT2), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n308), .A2(G148gat), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n317), .B1(new_n305), .B2(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n315), .A2(new_n312), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n311), .A2(new_n316), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n303), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT3), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n301), .B1(new_n324), .B2(new_n302), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n290), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT83), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n325), .A2(new_n289), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n321), .B(KEYINPUT78), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n329), .B1(new_n331), .B2(new_n303), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G22gat), .ZN(new_n334));
  INV_X1    g133(.A(G78gat), .ZN(new_n335));
  INV_X1    g134(.A(G22gat), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n328), .A2(new_n336), .A3(new_n332), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n335), .B1(new_n334), .B2(new_n337), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n288), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n340), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(new_n338), .A3(new_n287), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g143(.A1(G226gat), .A2(G233gat), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n252), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n345), .B1(new_n252), .B2(new_n302), .ZN(new_n347));
  INV_X1    g146(.A(new_n301), .ZN(new_n348));
  NOR3_X1   g147(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(G8gat), .B(G36gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(G64gat), .B(G92gat), .ZN(new_n352));
  XOR2_X1   g151(.A(new_n351), .B(new_n352), .Z(new_n353));
  OAI21_X1  g152(.A(new_n348), .B1(new_n346), .B2(new_n347), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n350), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT30), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n353), .B1(new_n350), .B2(new_n354), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n355), .A2(new_n360), .A3(new_n356), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n360), .B1(new_n355), .B2(new_n356), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n359), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G1gat), .B(G29gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n364), .B(KEYINPUT0), .ZN(new_n365));
  XNOR2_X1  g164(.A(G57gat), .B(G85gat), .ZN(new_n366));
  XOR2_X1   g165(.A(new_n365), .B(new_n366), .Z(new_n367));
  NAND2_X1  g166(.A1(G225gat), .A2(G233gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(KEYINPUT80), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n264), .A2(new_n321), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n372), .B1(new_n373), .B2(new_n370), .ZN(new_n374));
  XOR2_X1   g173(.A(new_n264), .B(KEYINPUT79), .Z(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(new_n324), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n331), .A2(new_n323), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n374), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n370), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n381), .B1(new_n375), .B2(new_n330), .ZN(new_n382));
  INV_X1    g181(.A(new_n369), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT5), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OR2_X1    g183(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n381), .A2(KEYINPUT4), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n369), .A2(KEYINPUT5), .ZN(new_n389));
  OAI211_X1 g188(.A(new_n388), .B(new_n389), .C1(new_n376), .C2(new_n378), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n367), .B1(new_n385), .B2(new_n390), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n390), .B(new_n367), .C1(new_n380), .C2(new_n384), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT6), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  AOI211_X1 g194(.A(new_n393), .B(new_n367), .C1(new_n385), .C2(new_n390), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n344), .B1(new_n363), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n278), .A2(new_n280), .ZN(new_n399));
  INV_X1    g198(.A(new_n279), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n401), .A2(KEYINPUT36), .A3(new_n281), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n284), .A2(new_n398), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n341), .A2(new_n343), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT37), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n350), .A2(new_n406), .A3(new_n354), .ZN(new_n407));
  INV_X1    g206(.A(new_n354), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT37), .B1(new_n408), .B2(new_n349), .ZN(new_n409));
  INV_X1    g208(.A(new_n353), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n407), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT38), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT38), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n407), .A2(new_n409), .A3(new_n413), .A4(new_n410), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n397), .A2(new_n412), .A3(new_n355), .A4(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT84), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT39), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n417), .B1(new_n382), .B2(new_n383), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n388), .B1(new_n376), .B2(new_n378), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n418), .B1(new_n420), .B2(new_n383), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n417), .A3(new_n369), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n367), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT40), .ZN(new_n424));
  AND2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n423), .A2(new_n424), .ZN(new_n426));
  NOR3_X1   g225(.A1(new_n425), .A2(new_n426), .A3(new_n391), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n363), .A2(new_n416), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n416), .B1(new_n363), .B2(new_n427), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n405), .B(new_n415), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n401), .A2(new_n281), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n363), .A2(new_n397), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n405), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT35), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n344), .B1(new_n401), .B2(new_n281), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT35), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n437), .A3(new_n433), .ZN(new_n438));
  AOI22_X1  g237(.A1(new_n404), .A2(new_n431), .B1(new_n435), .B2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(G113gat), .B(G141gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n440), .B(G197gat), .ZN(new_n441));
  XOR2_X1   g240(.A(KEYINPUT11), .B(G169gat), .Z(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  XOR2_X1   g242(.A(new_n443), .B(KEYINPUT12), .Z(new_n444));
  INV_X1    g243(.A(KEYINPUT14), .ZN(new_n445));
  INV_X1    g244(.A(G29gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n448));
  AOI21_X1  g247(.A(G36gat), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n446), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT15), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(G36gat), .ZN(new_n453));
  INV_X1    g252(.A(new_n448), .ZN(new_n454));
  NOR2_X1   g253(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n453), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT15), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(new_n450), .ZN(new_n458));
  XNOR2_X1  g257(.A(G43gat), .B(G50gat), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n452), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n459), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n461), .B(KEYINPUT15), .C1(new_n449), .C2(new_n451), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(KEYINPUT17), .A3(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(G15gat), .B(G22gat), .ZN(new_n464));
  INV_X1    g263(.A(G1gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT16), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n464), .A2(G1gat), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n467), .A2(new_n468), .A3(G8gat), .ZN(new_n469));
  INV_X1    g268(.A(G8gat), .ZN(new_n470));
  XOR2_X1   g269(.A(G15gat), .B(G22gat), .Z(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n465), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n464), .A2(new_n466), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n469), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n463), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT86), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n478));
  XOR2_X1   g277(.A(KEYINPUT85), .B(KEYINPUT17), .Z(new_n479));
  INV_X1    g278(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n477), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  AOI211_X1 g280(.A(KEYINPUT86), .B(new_n479), .C1(new_n460), .C2(new_n462), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n476), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G229gat), .A2(G233gat), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT87), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n485), .B1(new_n469), .B2(new_n474), .ZN(new_n486));
  OAI21_X1  g285(.A(G8gat), .B1(new_n467), .B2(new_n468), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n472), .A2(new_n470), .A3(new_n473), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT87), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n486), .A2(new_n478), .A3(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n483), .A2(KEYINPUT18), .A3(new_n484), .A4(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(KEYINPUT88), .ZN(new_n492));
  INV_X1    g291(.A(new_n478), .ZN(new_n493));
  NOR3_X1   g292(.A1(new_n469), .A2(new_n474), .A3(new_n485), .ZN(new_n494));
  AOI21_X1  g293(.A(KEYINPUT87), .B1(new_n487), .B2(new_n488), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n493), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT89), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(new_n490), .A3(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n494), .A2(new_n495), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(KEYINPUT89), .A3(new_n478), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  XOR2_X1   g300(.A(new_n484), .B(KEYINPUT13), .Z(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n483), .A2(new_n484), .A3(new_n490), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT18), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n444), .B1(new_n492), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT88), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n491), .B(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n444), .ZN(new_n511));
  AOI22_X1  g310(.A1(new_n501), .A2(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n439), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g315(.A1(G57gat), .A2(G64gat), .ZN(new_n517));
  AND2_X1   g316(.A1(G57gat), .A2(G64gat), .ZN(new_n518));
  INV_X1    g317(.A(G71gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n519), .A2(new_n335), .A3(KEYINPUT9), .ZN(new_n520));
  NAND2_X1  g319(.A1(G71gat), .A2(G78gat), .ZN(new_n521));
  AOI211_X1 g320(.A(new_n517), .B(new_n518), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  OR2_X1    g321(.A1(G57gat), .A2(G64gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT92), .ZN(new_n524));
  NAND2_X1  g323(.A1(G57gat), .A2(G64gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT92), .B1(new_n518), .B2(new_n517), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT9), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n521), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(KEYINPUT90), .B1(new_n519), .B2(new_n335), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n521), .A2(KEYINPUT91), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT91), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n533), .A2(G71gat), .A3(G78gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n531), .B1(new_n532), .B2(new_n534), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n530), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT93), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT90), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(G71gat), .B2(G78gat), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n533), .B1(G71gat), .B2(G78gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n521), .A2(KEYINPUT91), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n535), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n546), .A2(KEYINPUT93), .A3(new_n530), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n522), .B1(new_n540), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n548), .A2(KEYINPUT21), .ZN(new_n549));
  NAND2_X1  g348(.A1(G231gat), .A2(G233gat), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n549), .B(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(G127gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n499), .B1(KEYINPUT21), .B2(new_n548), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n552), .A2(new_n553), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n552), .A2(new_n553), .ZN(new_n558));
  INV_X1    g357(.A(new_n555), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(new_n313), .ZN(new_n563));
  XNOR2_X1  g362(.A(G183gat), .B(G211gat), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n563), .B(new_n564), .Z(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n561), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n556), .A2(new_n560), .A3(new_n565), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G190gat), .B(G218gat), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(G85gat), .A2(G92gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT7), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT7), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n574), .A2(G85gat), .A3(G92gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(G99gat), .B(G106gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578));
  INV_X1    g377(.A(G85gat), .ZN(new_n579));
  INV_X1    g378(.A(G92gat), .ZN(new_n580));
  AOI22_X1  g379(.A1(KEYINPUT8), .A2(new_n578), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n576), .A2(new_n577), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n577), .B1(new_n576), .B2(new_n581), .ZN(new_n583));
  NOR3_X1   g382(.A1(new_n582), .A2(new_n583), .A3(KEYINPUT95), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n583), .A2(KEYINPUT95), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n463), .B(new_n586), .C1(new_n481), .C2(new_n482), .ZN(new_n587));
  OR2_X1    g386(.A1(new_n584), .A2(new_n585), .ZN(new_n588));
  NAND2_X1  g387(.A1(G232gat), .A2(G233gat), .ZN(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AOI22_X1  g389(.A1(new_n588), .A2(new_n478), .B1(KEYINPUT41), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n571), .B1(new_n587), .B2(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n592), .A2(KEYINPUT97), .ZN(new_n593));
  AND3_X1   g392(.A1(new_n587), .A2(new_n571), .A3(new_n591), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n590), .A2(KEYINPUT41), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT94), .ZN(new_n596));
  XOR2_X1   g395(.A(G134gat), .B(G162gat), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n592), .A2(KEYINPUT97), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n593), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n598), .B1(new_n594), .B2(new_n592), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT96), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g403(.A(KEYINPUT96), .B(new_n598), .C1(new_n594), .C2(new_n592), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n601), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G120gat), .B(G148gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(G176gat), .B(G204gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT99), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT100), .ZN(new_n613));
  INV_X1    g412(.A(new_n522), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n546), .A2(KEYINPUT93), .A3(new_n530), .ZN(new_n615));
  AOI21_X1  g414(.A(KEYINPUT93), .B1(new_n546), .B2(new_n530), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT10), .B1(new_n584), .B2(new_n585), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n582), .A2(new_n583), .ZN(new_n620));
  OAI211_X1 g419(.A(new_n614), .B(new_n620), .C1(new_n615), .C2(new_n616), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n621), .B1(new_n548), .B2(new_n586), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT98), .B(KEYINPUT10), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n619), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G230gat), .A2(G233gat), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n613), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n617), .A2(new_n588), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n623), .B1(new_n629), .B2(new_n621), .ZN(new_n630));
  OAI211_X1 g429(.A(KEYINPUT100), .B(new_n626), .C1(new_n630), .C2(new_n619), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n629), .A2(new_n627), .A3(new_n621), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n612), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n622), .A2(new_n624), .ZN(new_n635));
  INV_X1    g434(.A(new_n619), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n626), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(new_n610), .A3(new_n633), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n634), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n569), .A2(new_n607), .A3(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n516), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n397), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(new_n465), .ZN(G1324gat));
  INV_X1    g446(.A(new_n644), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT101), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G8gat), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n648), .A2(new_n363), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n363), .ZN(new_n652));
  OAI21_X1  g451(.A(G8gat), .B1(new_n644), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  MUX2_X1   g453(.A(new_n651), .B(new_n654), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g454(.A1(new_n284), .A2(new_n402), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(G15gat), .B1(new_n644), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n432), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n659), .A2(G15gat), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n658), .B1(new_n644), .B2(new_n660), .ZN(G1326gat));
  NOR2_X1   g460(.A1(new_n644), .A2(new_n405), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT43), .B(G22gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1327gat));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n665), .B1(new_n439), .B2(new_n607), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n437), .B1(new_n436), .B2(new_n433), .ZN(new_n667));
  AND4_X1   g466(.A1(new_n437), .A2(new_n432), .A3(new_n405), .A4(new_n433), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n405), .A2(new_n415), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n363), .A2(new_n427), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(KEYINPUT84), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n669), .B1(new_n671), .B2(new_n428), .ZN(new_n672));
  OAI22_X1  g471(.A1(new_n667), .A2(new_n668), .B1(new_n672), .B2(new_n403), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n673), .A2(KEYINPUT44), .A3(new_n606), .ZN(new_n674));
  AND2_X1   g473(.A1(new_n666), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n641), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n569), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n514), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(KEYINPUT102), .Z(new_n679));
  NAND2_X1  g478(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(G29gat), .B1(new_n680), .B2(new_n645), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n439), .A2(new_n607), .A3(new_n678), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n446), .A3(new_n397), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT45), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n684), .ZN(G1328gat));
  NAND3_X1  g484(.A1(new_n682), .A2(new_n453), .A3(new_n363), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n686), .B(KEYINPUT46), .Z(new_n687));
  OAI21_X1  g486(.A(G36gat), .B1(new_n680), .B2(new_n652), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(G1329gat));
  NAND4_X1  g488(.A1(new_n666), .A2(new_n656), .A3(new_n674), .A4(new_n679), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n659), .A2(G43gat), .ZN(new_n691));
  AOI22_X1  g490(.A1(new_n690), .A2(G43gat), .B1(new_n682), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(KEYINPUT103), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT47), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1330gat));
  NOR2_X1   g494(.A1(new_n607), .A2(G50gat), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n516), .A2(new_n344), .A3(new_n677), .A4(new_n696), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n666), .A2(new_n344), .A3(new_n674), .A4(new_n679), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT104), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(G50gat), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n698), .A2(KEYINPUT104), .ZN(new_n701));
  OAI211_X1 g500(.A(KEYINPUT48), .B(new_n697), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n698), .A2(G50gat), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n703), .A2(new_n697), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(KEYINPUT48), .B2(new_n704), .ZN(G1331gat));
  INV_X1    g504(.A(new_n568), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n565), .B1(new_n556), .B2(new_n560), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(new_n606), .ZN(new_n709));
  AND4_X1   g508(.A1(new_n515), .A2(new_n673), .A3(new_n709), .A4(new_n676), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n397), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g511(.A(new_n652), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(KEYINPUT105), .ZN(new_n715));
  NOR2_X1   g514(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n715), .B(new_n716), .ZN(G1333gat));
  AOI21_X1  g516(.A(new_n519), .B1(new_n710), .B2(new_n656), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n659), .A2(G71gat), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n718), .B1(new_n710), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g520(.A1(new_n710), .A2(new_n344), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n515), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT106), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n725), .A2(new_n676), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n675), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(G85gat), .B1(new_n727), .B2(new_n645), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n673), .A2(new_n606), .A3(new_n725), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT51), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n673), .A2(KEYINPUT51), .A3(new_n606), .A4(new_n725), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n729), .A2(KEYINPUT107), .A3(new_n730), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n734), .A2(new_n735), .A3(new_n676), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n397), .A2(new_n579), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n728), .B1(new_n736), .B2(new_n737), .ZN(G1336gat));
  NAND3_X1  g537(.A1(new_n363), .A2(new_n580), .A3(new_n676), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(KEYINPUT108), .Z(new_n740));
  NAND3_X1  g539(.A1(new_n734), .A2(new_n735), .A3(new_n740), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n666), .A2(new_n363), .A3(new_n674), .A4(new_n726), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT52), .B1(new_n742), .B2(G92gat), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n741), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n731), .A2(new_n733), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n740), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n742), .A2(G92gat), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n745), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(KEYINPUT109), .B1(new_n744), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n741), .A2(new_n743), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n747), .A2(new_n748), .ZN(new_n753));
  OAI211_X1 g552(.A(new_n751), .B(new_n752), .C1(new_n753), .C2(new_n745), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n750), .A2(new_n754), .ZN(G1337gat));
  OAI21_X1  g554(.A(G99gat), .B1(new_n727), .B2(new_n657), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n659), .A2(G99gat), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n736), .B2(new_n757), .ZN(G1338gat));
  NAND4_X1  g557(.A1(new_n666), .A2(new_n344), .A3(new_n674), .A4(new_n726), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G106gat), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n405), .A2(G106gat), .A3(new_n641), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n762), .B1(new_n731), .B2(new_n733), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n760), .B1(new_n763), .B2(KEYINPUT110), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n763), .A2(KEYINPUT110), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT53), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n734), .A2(new_n735), .A3(new_n761), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n759), .A2(KEYINPUT111), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G106gat), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n759), .A2(KEYINPUT111), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n767), .B(new_n768), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n766), .A2(new_n772), .ZN(G1339gat));
  INV_X1    g572(.A(KEYINPUT118), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n363), .A2(new_n645), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n432), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT116), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n628), .A2(new_n780), .A3(new_n631), .ZN(new_n781));
  INV_X1    g580(.A(new_n610), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(KEYINPUT54), .B1(new_n625), .B2(new_n627), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n637), .B2(new_n626), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n625), .A2(KEYINPUT113), .A3(new_n627), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n784), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n779), .B1(new_n783), .B2(new_n788), .ZN(new_n789));
  NOR4_X1   g588(.A1(new_n630), .A2(new_n785), .A3(new_n626), .A4(new_n619), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT113), .B1(new_n625), .B2(new_n627), .ZN(new_n791));
  OAI211_X1 g590(.A(KEYINPUT54), .B(new_n638), .C1(new_n790), .C2(new_n791), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n792), .A2(KEYINPUT55), .A3(new_n782), .A4(new_n781), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n514), .A2(new_n789), .A3(new_n639), .A4(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n501), .A2(new_n502), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n484), .B1(new_n483), .B2(new_n490), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n443), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n513), .B(new_n797), .C1(new_n634), .C2(new_n640), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n607), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n789), .A2(new_n793), .A3(new_n639), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n606), .A2(new_n513), .A3(new_n797), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n800), .A2(new_n801), .A3(new_n805), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n606), .B1(new_n794), .B2(new_n798), .ZN(new_n807));
  OAI21_X1  g606(.A(KEYINPUT114), .B1(new_n807), .B2(new_n804), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n806), .A2(new_n708), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n709), .A2(new_n810), .A3(new_n515), .A4(new_n641), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT112), .B1(new_n642), .B2(new_n514), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n809), .A2(KEYINPUT115), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT115), .B1(new_n809), .B2(new_n813), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n778), .B1(new_n816), .B2(new_n405), .ZN(new_n817));
  NOR4_X1   g616(.A1(new_n814), .A2(new_n815), .A3(KEYINPUT116), .A4(new_n344), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n777), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI211_X1 g620(.A(KEYINPUT117), .B(new_n777), .C1(new_n817), .C2(new_n818), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(new_n514), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G113gat), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n813), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n809), .A2(new_n813), .A3(KEYINPUT115), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(new_n645), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n436), .ZN(new_n831));
  NOR4_X1   g630(.A1(new_n831), .A2(G113gat), .A3(new_n515), .A4(new_n363), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n774), .B1(new_n824), .B2(new_n833), .ZN(new_n834));
  AOI211_X1 g633(.A(KEYINPUT118), .B(new_n832), .C1(new_n823), .C2(G113gat), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(G1340gat));
  NOR2_X1   g635(.A1(new_n831), .A2(new_n363), .ZN(new_n837));
  AOI21_X1  g636(.A(G120gat), .B1(new_n837), .B2(new_n676), .ZN(new_n838));
  INV_X1    g637(.A(new_n821), .ZN(new_n839));
  INV_X1    g638(.A(new_n822), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n641), .A2(new_n255), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n838), .B1(new_n841), .B2(new_n842), .ZN(G1341gat));
  NAND3_X1  g642(.A1(new_n837), .A2(new_n553), .A3(new_n569), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n839), .A2(new_n708), .A3(new_n840), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n844), .B1(new_n845), .B2(new_n553), .ZN(G1342gat));
  INV_X1    g645(.A(G134gat), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n363), .A2(new_n607), .ZN(new_n848));
  NAND4_X1  g647(.A1(new_n830), .A2(new_n847), .A3(new_n436), .A4(new_n848), .ZN(new_n849));
  XOR2_X1   g648(.A(new_n849), .B(KEYINPUT56), .Z(new_n850));
  NOR3_X1   g649(.A1(new_n839), .A2(new_n607), .A3(new_n840), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n850), .B1(new_n851), .B2(new_n847), .ZN(G1343gat));
  AOI21_X1  g651(.A(KEYINPUT57), .B1(new_n816), .B2(new_n344), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT57), .ZN(new_n854));
  INV_X1    g653(.A(new_n798), .ZN(new_n855));
  XOR2_X1   g654(.A(new_n789), .B(KEYINPUT119), .Z(new_n856));
  NAND3_X1  g655(.A1(new_n514), .A2(new_n639), .A3(new_n793), .ZN(new_n857));
  INV_X1    g656(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n855), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n805), .B1(new_n859), .B2(new_n606), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n708), .ZN(new_n861));
  AOI211_X1 g660(.A(new_n854), .B(new_n405), .C1(new_n861), .C2(new_n813), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n853), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n657), .A2(new_n775), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n514), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT58), .B1(new_n866), .B2(G141gat), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n656), .A2(new_n405), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n830), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT120), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n830), .A2(new_n871), .A3(new_n868), .ZN(new_n872));
  AND2_X1   g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n873), .A2(new_n308), .A3(new_n514), .A4(new_n652), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n867), .A2(new_n874), .ZN(new_n875));
  NOR4_X1   g674(.A1(new_n869), .A2(G141gat), .A3(new_n515), .A4(new_n363), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n876), .B1(new_n866), .B2(G141gat), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(G1344gat));
  NAND3_X1  g678(.A1(new_n873), .A2(new_n652), .A3(new_n676), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT59), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n304), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n816), .A2(KEYINPUT57), .A3(new_n344), .ZN(new_n883));
  AOI22_X1  g682(.A1(new_n860), .A2(new_n708), .B1(new_n515), .B2(new_n643), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n854), .B1(new_n884), .B2(new_n405), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n886), .A2(new_n657), .A3(new_n676), .A4(new_n775), .ZN(new_n887));
  AND2_X1   g686(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n888));
  INV_X1    g687(.A(new_n863), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n864), .A2(KEYINPUT59), .A3(new_n641), .ZN(new_n890));
  AOI22_X1  g689(.A1(new_n887), .A2(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n882), .A2(new_n891), .ZN(G1345gat));
  AOI21_X1  g691(.A(new_n313), .B1(new_n865), .B2(new_n569), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n708), .A2(G155gat), .ZN(new_n894));
  AND4_X1   g693(.A1(new_n652), .A2(new_n870), .A3(new_n872), .A4(new_n894), .ZN(new_n895));
  OR3_X1    g694(.A1(new_n893), .A2(new_n895), .A3(KEYINPUT121), .ZN(new_n896));
  OAI21_X1  g695(.A(KEYINPUT121), .B1(new_n893), .B2(new_n895), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1346gat));
  NAND3_X1  g697(.A1(new_n873), .A2(new_n314), .A3(new_n848), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n863), .A2(new_n607), .A3(new_n864), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(new_n314), .ZN(G1347gat));
  NAND2_X1  g700(.A1(new_n436), .A2(new_n363), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT122), .B1(new_n829), .B2(new_n397), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n816), .A2(new_n904), .A3(new_n645), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n902), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(G169gat), .B1(new_n906), .B2(new_n514), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n652), .A2(new_n397), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(new_n432), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT123), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT116), .B1(new_n829), .B2(new_n344), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n816), .A2(new_n778), .A3(new_n405), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n515), .A2(new_n209), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n907), .B1(new_n913), .B2(new_n914), .ZN(G1348gat));
  NAND3_X1  g714(.A1(new_n906), .A2(new_n210), .A3(new_n676), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n913), .A2(new_n676), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(new_n210), .ZN(G1349gat));
  NAND3_X1  g717(.A1(new_n906), .A2(new_n238), .A3(new_n569), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n913), .A2(new_n569), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n919), .B1(new_n920), .B2(new_n220), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g721(.A1(new_n906), .A2(new_n221), .A3(new_n606), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT61), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n913), .A2(new_n606), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n925), .B2(G190gat), .ZN(new_n926));
  AOI211_X1 g725(.A(KEYINPUT61), .B(new_n221), .C1(new_n913), .C2(new_n606), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(G1351gat));
  NAND2_X1  g727(.A1(new_n903), .A2(new_n905), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n868), .A2(new_n363), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT124), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n929), .A2(KEYINPUT124), .A3(new_n931), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n515), .A2(G197gat), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n657), .A2(new_n908), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n937), .B1(new_n883), .B2(new_n885), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(G197gat), .B1(new_n939), .B2(new_n515), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n936), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT125), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n936), .A2(new_n943), .A3(new_n940), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(G1352gat));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n947));
  INV_X1    g746(.A(G204gat), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n676), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n946), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n948), .B1(new_n938), .B2(new_n676), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n953), .B1(new_n950), .B2(new_n951), .ZN(new_n954));
  OAI211_X1 g753(.A(KEYINPUT126), .B(KEYINPUT62), .C1(new_n947), .C2(new_n949), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n952), .A2(new_n954), .A3(new_n955), .ZN(G1353gat));
  AOI21_X1  g755(.A(new_n292), .B1(new_n938), .B2(new_n569), .ZN(new_n957));
  OR3_X1    g756(.A1(new_n957), .A2(KEYINPUT127), .A3(KEYINPUT63), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n957), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n959));
  NAND2_X1  g758(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n933), .A2(new_n292), .A3(new_n569), .A4(new_n934), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(G1354gat));
  NAND4_X1  g762(.A1(new_n933), .A2(new_n293), .A3(new_n606), .A4(new_n934), .ZN(new_n964));
  OAI21_X1  g763(.A(G218gat), .B1(new_n939), .B2(new_n607), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1355gat));
endmodule


