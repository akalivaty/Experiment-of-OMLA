//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1228, new_n1229, new_n1230, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n202), .A2(G77), .A3(new_n204), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n204), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n210), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(KEYINPUT65), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n223), .A2(new_n224), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n212), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n215), .B(new_n220), .C1(new_n230), .C2(KEYINPUT1), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G238), .B(G244), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XOR2_X1   g0041(.A(G50), .B(G58), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G351));
  INV_X1    g0047(.A(G41), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(KEYINPUT66), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT66), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G41), .ZN(new_n251));
  INV_X1    g0051(.A(G45), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT67), .ZN(new_n254));
  AND3_X1   g0054(.A1(new_n253), .A2(new_n254), .A3(new_n209), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n254), .B1(new_n253), .B2(new_n209), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT68), .ZN(new_n257));
  AND2_X1   g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n257), .B1(new_n258), .B2(new_n218), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n260), .A2(KEYINPUT68), .A3(G1), .A4(G13), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n259), .A2(G274), .A3(new_n261), .ZN(new_n262));
  NOR3_X1   g0062(.A1(new_n255), .A2(new_n256), .A3(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n264));
  AND3_X1   g0064(.A1(new_n259), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n263), .B1(G226), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n258), .A2(new_n218), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G1698), .ZN(new_n274));
  INV_X1    g0074(.A(G223), .ZN(new_n275));
  INV_X1    g0075(.A(G77), .ZN(new_n276));
  OAI22_X1  g0076(.A1(new_n274), .A2(new_n275), .B1(new_n276), .B2(new_n273), .ZN(new_n277));
  AOI21_X1  g0077(.A(G1698), .B1(new_n271), .B2(new_n272), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n277), .B1(G222), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n266), .B1(new_n268), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G200), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n218), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT8), .B(G58), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n210), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(G150), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n284), .A2(new_n285), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n210), .B1(new_n201), .B2(new_n203), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n283), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(new_n283), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n209), .A2(G20), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n294), .A2(G50), .A3(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n291), .B(new_n296), .C1(G50), .C2(new_n292), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT9), .ZN(new_n298));
  INV_X1    g0098(.A(G190), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n281), .B(new_n298), .C1(new_n299), .C2(new_n280), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT10), .ZN(new_n301));
  XOR2_X1   g0101(.A(KEYINPUT69), .B(G179), .Z(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n280), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n280), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n304), .A2(new_n297), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n301), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n256), .A2(new_n262), .ZN(new_n309));
  INV_X1    g0109(.A(new_n255), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G226), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G1698), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n313), .B1(G223), .B2(G1698), .ZN(new_n314));
  AND2_X1   g0114(.A1(KEYINPUT3), .A2(G33), .ZN(new_n315));
  NOR2_X1   g0115(.A1(KEYINPUT3), .A2(G33), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G87), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n314), .A2(new_n317), .B1(new_n270), .B2(new_n318), .ZN(new_n319));
  AOI22_X1  g0119(.A1(G232), .A2(new_n265), .B1(new_n319), .B2(new_n267), .ZN(new_n320));
  AOI21_X1  g0120(.A(G169), .B1(new_n311), .B2(new_n320), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n259), .A2(G232), .A3(new_n261), .A4(new_n264), .ZN(new_n322));
  NOR2_X1   g0122(.A1(G223), .A2(G1698), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n323), .B1(new_n312), .B2(G1698), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n324), .A2(new_n273), .B1(G33), .B2(G87), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n322), .B1(new_n325), .B2(new_n268), .ZN(new_n326));
  NOR3_X1   g0126(.A1(new_n263), .A2(new_n326), .A3(new_n303), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n321), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT16), .ZN(new_n329));
  INV_X1    g0129(.A(G68), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT7), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n331), .B1(new_n273), .B2(G20), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n317), .A2(KEYINPUT7), .A3(new_n210), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n330), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G58), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n335), .A2(new_n330), .ZN(new_n336));
  OAI21_X1  g0136(.A(G20), .B1(new_n336), .B2(new_n203), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n287), .A2(G159), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n329), .B1(new_n334), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT7), .B1(new_n317), .B2(new_n210), .ZN(new_n341));
  NOR4_X1   g0141(.A1(new_n315), .A2(new_n316), .A3(new_n331), .A4(G20), .ZN(new_n342));
  OAI21_X1  g0142(.A(G68), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n339), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n343), .A2(KEYINPUT16), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n340), .A2(new_n283), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n284), .B1(new_n209), .B2(G20), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n347), .A2(new_n294), .B1(new_n293), .B2(new_n284), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n328), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT18), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT18), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n328), .A2(new_n349), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n348), .ZN(new_n355));
  INV_X1    g0155(.A(new_n283), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n343), .A2(new_n344), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n356), .B1(new_n357), .B2(new_n329), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n355), .B1(new_n358), .B2(new_n345), .ZN(new_n359));
  INV_X1    g0159(.A(G200), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n263), .B2(new_n326), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n311), .A2(new_n320), .A3(new_n299), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n359), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT77), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT17), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n359), .A2(new_n363), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n365), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n265), .A2(G244), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n311), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT70), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n311), .A2(KEYINPUT70), .A3(new_n370), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n278), .A2(G232), .ZN(new_n375));
  INV_X1    g0175(.A(G107), .ZN(new_n376));
  INV_X1    g0176(.A(G238), .ZN(new_n377));
  OAI221_X1 g0177(.A(new_n375), .B1(new_n376), .B2(new_n273), .C1(new_n377), .C2(new_n274), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n267), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n373), .A2(new_n374), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n305), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n356), .A2(KEYINPUT71), .A3(new_n292), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT71), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n293), .B2(new_n283), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n382), .A2(new_n384), .A3(new_n295), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G77), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n293), .A2(new_n276), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n284), .A2(new_n288), .B1(new_n210), .B2(new_n276), .ZN(new_n388));
  XNOR2_X1  g0188(.A(KEYINPUT15), .B(G87), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n389), .A2(new_n285), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n283), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n386), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  NAND4_X1  g0192(.A1(new_n373), .A2(new_n302), .A3(new_n374), .A4(new_n379), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n381), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n380), .A2(G200), .ZN(new_n395));
  INV_X1    g0195(.A(new_n392), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n380), .B2(new_n299), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n394), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  NOR4_X1   g0198(.A1(new_n308), .A2(new_n354), .A3(new_n369), .A4(new_n398), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n309), .A2(new_n310), .B1(G238), .B2(new_n265), .ZN(new_n400));
  INV_X1    g0200(.A(G1698), .ZN(new_n401));
  OAI211_X1 g0201(.A(G226), .B(new_n401), .C1(new_n315), .C2(new_n316), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G97), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI211_X1 g0204(.A(G232), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT72), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n273), .A2(KEYINPUT72), .A3(G232), .A4(G1698), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n404), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n267), .B1(new_n409), .B2(KEYINPUT73), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT73), .ZN(new_n411));
  AOI211_X1 g0211(.A(new_n411), .B(new_n404), .C1(new_n407), .C2(new_n408), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n400), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT13), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT13), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n400), .B(new_n415), .C1(new_n410), .C2(new_n412), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(G190), .A3(new_n416), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n417), .B(KEYINPUT75), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT74), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n414), .A2(new_n419), .A3(new_n416), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n413), .A2(KEYINPUT74), .A3(KEYINPUT13), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(G200), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(G50), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n288), .A2(new_n423), .B1(new_n210), .B2(G68), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n285), .A2(new_n276), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n283), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n426), .B(KEYINPUT11), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n385), .A2(G68), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT76), .ZN(new_n429));
  AOI211_X1 g0229(.A(G68), .B(new_n292), .C1(new_n429), .C2(KEYINPUT12), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n429), .A2(KEYINPUT12), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n430), .B(new_n431), .ZN(new_n432));
  AND3_X1   g0232(.A1(new_n427), .A2(new_n428), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n422), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n418), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n433), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n420), .A2(G169), .A3(new_n421), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT14), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n414), .A2(G179), .A3(new_n416), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT14), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n420), .A2(new_n440), .A3(G169), .A4(new_n421), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n438), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n435), .B1(new_n436), .B2(new_n442), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n399), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT83), .ZN(new_n445));
  OAI211_X1 g0245(.A(G244), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(KEYINPUT80), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT80), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n273), .A2(new_n448), .A3(G244), .A4(G1698), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G116), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n273), .A2(G238), .A3(new_n401), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n447), .A2(new_n449), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n267), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n209), .A2(G45), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n454), .A2(G274), .ZN(new_n455));
  INV_X1    g0255(.A(G250), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  AND4_X1   g0257(.A1(new_n259), .A2(new_n455), .A3(new_n261), .A4(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n360), .B1(new_n453), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n273), .A2(new_n210), .A3(G68), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT19), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n210), .B1(new_n403), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(G87), .B2(new_n207), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n210), .A2(G33), .A3(G97), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT82), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n465), .A2(new_n466), .A3(new_n462), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n466), .B1(new_n465), .B2(new_n462), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n461), .B(new_n464), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n283), .ZN(new_n470));
  INV_X1    g0270(.A(new_n389), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(new_n292), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n209), .A2(G33), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n292), .A2(new_n474), .A3(new_n218), .A4(new_n282), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(new_n318), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n470), .A2(new_n473), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n445), .B1(new_n460), .B2(new_n478), .ZN(new_n479));
  AOI211_X1 g0279(.A(new_n472), .B(new_n476), .C1(new_n469), .C2(new_n283), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n458), .B1(new_n452), .B2(new_n267), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n480), .B(KEYINPUT83), .C1(new_n360), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(G190), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n479), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n481), .A2(new_n302), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT81), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n481), .A2(KEYINPUT81), .A3(new_n302), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n453), .A2(new_n459), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n305), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n470), .B(new_n473), .C1(new_n389), .C2(new_n475), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n487), .A2(new_n488), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n484), .A2(KEYINPUT84), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT84), .B1(new_n484), .B2(new_n492), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g0295(.A(KEYINPUT85), .B(KEYINPUT22), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n210), .B(G87), .C1(new_n315), .C2(new_n316), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n273), .A2(new_n496), .A3(new_n210), .A4(G87), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n450), .A2(G20), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT23), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n210), .B2(G107), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n376), .A2(KEYINPUT23), .A3(G20), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n501), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n499), .A2(new_n500), .A3(new_n505), .ZN(new_n506));
  XNOR2_X1  g0306(.A(KEYINPUT86), .B(KEYINPUT24), .ZN(new_n507));
  INV_X1    g0307(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n499), .A2(new_n500), .A3(new_n507), .A4(new_n505), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n283), .ZN(new_n512));
  AND2_X1   g0312(.A1(new_n259), .A2(new_n261), .ZN(new_n513));
  INV_X1    g0313(.A(new_n454), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n248), .A2(KEYINPUT5), .ZN(new_n515));
  XNOR2_X1  g0315(.A(KEYINPUT66), .B(G41), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n514), .B(new_n515), .C1(new_n516), .C2(KEYINPUT5), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n513), .A2(new_n517), .A3(G264), .ZN(new_n518));
  OAI211_X1 g0318(.A(G257), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n519));
  OAI211_X1 g0319(.A(G250), .B(new_n401), .C1(new_n315), .C2(new_n316), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G294), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n267), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT79), .ZN(new_n524));
  AOI21_X1  g0324(.A(KEYINPUT5), .B1(new_n249), .B2(new_n251), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(new_n454), .ZN(new_n526));
  OAI211_X1 g0326(.A(KEYINPUT79), .B(new_n514), .C1(new_n516), .C2(KEYINPUT5), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n259), .A2(G274), .A3(new_n261), .A4(new_n515), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n518), .B(new_n523), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G200), .ZN(new_n531));
  INV_X1    g0331(.A(new_n475), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n293), .A2(KEYINPUT25), .A3(new_n376), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT25), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n292), .B2(G107), .ZN(new_n535));
  AOI22_X1  g0335(.A1(G107), .A2(new_n532), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  AND3_X1   g0336(.A1(new_n259), .A2(G274), .A3(new_n261), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n537), .A2(new_n526), .A3(new_n515), .A4(new_n527), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n538), .A2(G190), .A3(new_n518), .A4(new_n523), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n512), .A2(new_n531), .A3(new_n536), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n530), .A2(new_n305), .ZN(new_n541));
  INV_X1    g0341(.A(G179), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n538), .A2(new_n542), .A3(new_n518), .A4(new_n523), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n356), .B1(new_n509), .B2(new_n510), .ZN(new_n544));
  INV_X1    g0344(.A(new_n536), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n541), .B(new_n543), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G283), .ZN(new_n547));
  OAI211_X1 g0347(.A(G250), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n548));
  OAI211_X1 g0348(.A(G244), .B(new_n401), .C1(new_n315), .C2(new_n316), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT4), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n547), .B(new_n548), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(KEYINPUT4), .B1(new_n278), .B2(G244), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n267), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n513), .A2(new_n517), .A3(G257), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n538), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n305), .ZN(new_n556));
  AND2_X1   g0356(.A1(G97), .A2(G107), .ZN(new_n557));
  OAI22_X1  g0357(.A1(new_n557), .A2(new_n206), .B1(KEYINPUT78), .B2(KEYINPUT6), .ZN(new_n558));
  NOR2_X1   g0358(.A1(KEYINPUT78), .A2(KEYINPUT6), .ZN(new_n559));
  INV_X1    g0359(.A(G97), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n559), .B1(KEYINPUT6), .B2(new_n560), .ZN(new_n561));
  XNOR2_X1  g0361(.A(G97), .B(G107), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n558), .B(G20), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n287), .A2(G77), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n376), .B1(new_n332), .B2(new_n333), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n283), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n293), .A2(new_n560), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n532), .A2(G97), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n553), .A2(new_n538), .A3(new_n302), .A4(new_n554), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n556), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n555), .A2(G200), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n569), .A2(new_n568), .ZN(new_n574));
  OAI21_X1  g0374(.A(G107), .B1(new_n341), .B2(new_n342), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n575), .A2(new_n563), .A3(new_n564), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n574), .B1(new_n576), .B2(new_n283), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n553), .A2(new_n538), .A3(G190), .A4(new_n554), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n573), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n540), .A2(new_n546), .A3(new_n572), .A4(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(G264), .B(G1698), .C1(new_n315), .C2(new_n316), .ZN(new_n581));
  OAI211_X1 g0381(.A(G257), .B(new_n401), .C1(new_n315), .C2(new_n316), .ZN(new_n582));
  INV_X1    g0382(.A(G303), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n581), .B(new_n582), .C1(new_n583), .C2(new_n273), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n267), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n513), .A2(new_n517), .A3(G270), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n538), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n382), .A2(new_n384), .A3(G116), .A4(new_n474), .ZN(new_n588));
  INV_X1    g0388(.A(G13), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n589), .A2(G1), .ZN(new_n590));
  INV_X1    g0390(.A(G116), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n590), .A2(G20), .A3(new_n591), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n547), .B(new_n210), .C1(G33), .C2(new_n560), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n593), .B(new_n283), .C1(new_n210), .C2(G116), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT20), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n594), .A2(new_n595), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n588), .B(new_n592), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n587), .A2(new_n598), .A3(G169), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT21), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n587), .A2(G200), .ZN(new_n602));
  INV_X1    g0402(.A(new_n598), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n538), .A2(G190), .A3(new_n585), .A4(new_n586), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  AND4_X1   g0405(.A1(G179), .A2(new_n538), .A3(new_n585), .A4(new_n586), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n598), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n587), .A2(new_n598), .A3(KEYINPUT21), .A4(G169), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n601), .A2(new_n605), .A3(new_n607), .A4(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n580), .A2(new_n609), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n444), .A2(new_n495), .A3(new_n610), .ZN(G372));
  INV_X1    g0411(.A(KEYINPUT87), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n489), .A2(new_n612), .A3(new_n305), .ZN(new_n613));
  OAI21_X1  g0413(.A(KEYINPUT87), .B1(new_n481), .B2(G169), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n485), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT88), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT88), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n613), .A2(new_n614), .A3(new_n617), .A4(new_n485), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n491), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT26), .ZN(new_n621));
  INV_X1    g0421(.A(new_n572), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n483), .B(new_n480), .C1(new_n360), .C2(new_n481), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n620), .A2(new_n621), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  AND2_X1   g0424(.A1(new_n607), .A2(new_n608), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n625), .A2(new_n601), .A3(new_n546), .ZN(new_n626));
  AND4_X1   g0426(.A1(new_n540), .A2(new_n572), .A3(new_n579), .A4(new_n623), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n626), .A2(new_n627), .B1(new_n619), .B2(new_n491), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n493), .A2(new_n494), .A3(new_n572), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n624), .B(new_n628), .C1(new_n629), .C2(new_n621), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n444), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n307), .ZN(new_n632));
  INV_X1    g0432(.A(new_n353), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n352), .B1(new_n328), .B2(new_n349), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n435), .A2(new_n369), .ZN(new_n636));
  INV_X1    g0436(.A(new_n394), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n637), .B1(new_n442), .B2(new_n436), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n635), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n632), .B1(new_n639), .B2(new_n301), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n631), .A2(new_n640), .ZN(G369));
  NAND2_X1  g0441(.A1(new_n625), .A2(new_n601), .ZN(new_n642));
  INV_X1    g0442(.A(new_n590), .ZN(new_n643));
  OR3_X1    g0443(.A1(new_n643), .A2(KEYINPUT27), .A3(G20), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT27), .B1(new_n643), .B2(G20), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n644), .A2(G213), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(G343), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n603), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n642), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n649), .B1(new_n609), .B2(new_n648), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(G330), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n546), .ZN(new_n653));
  INV_X1    g0453(.A(new_n647), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(KEYINPUT89), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n654), .B1(new_n544), .B2(new_n545), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n540), .A2(new_n546), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT89), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n658), .B1(new_n546), .B2(new_n647), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n655), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n652), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n654), .B1(new_n625), .B2(new_n601), .ZN(new_n662));
  AOI22_X1  g0462(.A1(new_n660), .A2(new_n662), .B1(new_n653), .B2(new_n647), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(G399));
  NAND2_X1  g0464(.A1(new_n213), .A2(new_n516), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n665), .A2(G1), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n216), .B2(new_n665), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT28), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n530), .A2(new_n302), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n670), .A2(new_n489), .A3(new_n587), .A4(new_n555), .ZN(new_n671));
  AND4_X1   g0471(.A1(new_n453), .A2(new_n459), .A3(new_n518), .A4(new_n523), .ZN(new_n672));
  INV_X1    g0472(.A(new_n555), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT30), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT90), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n672), .A2(new_n606), .A3(new_n673), .A4(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n481), .A2(new_n518), .A3(new_n523), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(new_n555), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n675), .B1(new_n679), .B2(new_n606), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n654), .B1(new_n677), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT31), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OAI211_X1 g0483(.A(KEYINPUT31), .B(new_n654), .C1(new_n677), .C2(new_n680), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n685), .A2(KEYINPUT91), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n495), .A2(new_n610), .A3(new_n647), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(KEYINPUT91), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n689), .A2(G330), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n484), .A2(new_n492), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT84), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n484), .A2(KEYINPUT84), .A3(new_n492), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n693), .A2(new_n621), .A3(new_n694), .A4(new_n622), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(new_n628), .ZN(new_n696));
  INV_X1    g0496(.A(new_n623), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n619), .B2(new_n491), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n621), .B1(new_n698), .B2(new_n622), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n647), .B1(new_n696), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(KEYINPUT92), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI211_X1 g0502(.A(KEYINPUT92), .B(new_n647), .C1(new_n696), .C2(new_n699), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT29), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n630), .A2(new_n647), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT29), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n690), .B1(new_n705), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n669), .B1(new_n709), .B2(G1), .ZN(G364));
  INV_X1    g0510(.A(new_n665), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n589), .A2(G20), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n209), .B1(new_n712), .B2(G45), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g0515(.A(new_n715), .B(KEYINPUT93), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n213), .A2(new_n273), .ZN(new_n717));
  INV_X1    g0517(.A(G355), .ZN(new_n718));
  OAI22_X1  g0518(.A1(new_n717), .A2(new_n718), .B1(G116), .B2(new_n213), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n243), .A2(G45), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n213), .A2(new_n317), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n721), .B1(new_n252), .B2(new_n217), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n719), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(G13), .A2(G33), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G20), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n218), .B1(G20), .B2(new_n305), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n716), .B1(new_n723), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(G283), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n210), .A2(G179), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(new_n299), .A3(G200), .ZN(new_n733));
  NOR4_X1   g0533(.A1(new_n302), .A2(new_n210), .A3(new_n299), .A4(G200), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G322), .ZN(new_n736));
  OAI221_X1 g0536(.A(new_n317), .B1(new_n731), .B2(new_n733), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n210), .A2(G190), .A3(G200), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n303), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n542), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n739), .A2(G311), .B1(new_n741), .B2(G329), .ZN(new_n742));
  INV_X1    g0542(.A(G294), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n299), .A2(G179), .A3(G200), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n210), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n742), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n732), .A2(G190), .A3(G200), .ZN(new_n747));
  OR2_X1    g0547(.A1(new_n747), .A2(KEYINPUT95), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(KEYINPUT95), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI211_X1 g0551(.A(new_n737), .B(new_n746), .C1(G303), .C2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G326), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n303), .A2(G20), .A3(G200), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT94), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n756), .A2(G190), .A3(new_n757), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n752), .B1(new_n753), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n756), .A2(new_n299), .A3(new_n757), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(KEYINPUT33), .B(G317), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n763), .A2(KEYINPUT96), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(KEYINPUT96), .ZN(new_n765));
  INV_X1    g0565(.A(new_n745), .ZN(new_n766));
  INV_X1    g0566(.A(new_n733), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n766), .A2(G97), .B1(new_n767), .B2(G107), .ZN(new_n768));
  INV_X1    g0568(.A(new_n739), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n273), .B(new_n768), .C1(new_n769), .C2(new_n276), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n770), .B1(G87), .B2(new_n751), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n741), .A2(G159), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n735), .A2(new_n335), .B1(KEYINPUT32), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n773), .B1(KEYINPUT32), .B2(new_n772), .ZN(new_n774));
  AND2_X1   g0574(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n775), .B1(new_n423), .B2(new_n758), .C1(new_n330), .C2(new_n760), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n764), .A2(new_n765), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n730), .B1(new_n777), .B2(new_n727), .ZN(new_n778));
  INV_X1    g0578(.A(new_n726), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n778), .B1(new_n650), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT97), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n652), .A2(new_n715), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(G330), .B2(new_n650), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n781), .A2(new_n783), .ZN(G396));
  INV_X1    g0584(.A(new_n715), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n394), .A2(new_n654), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n395), .A2(new_n397), .B1(new_n396), .B2(new_n647), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n786), .B1(new_n394), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n630), .A2(new_n647), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(KEYINPUT99), .ZN(new_n790));
  INV_X1    g0590(.A(new_n788), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n790), .A2(new_n706), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n706), .A2(new_n791), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n793), .A2(KEYINPUT99), .A3(new_n789), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n690), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT100), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(KEYINPUT100), .B1(new_n795), .B2(new_n690), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n785), .B1(new_n690), .B2(new_n795), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n733), .A2(new_n330), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n317), .ZN(new_n802));
  INV_X1    g0602(.A(G132), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n802), .B1(new_n335), .B2(new_n745), .C1(new_n803), .C2(new_n740), .ZN(new_n804));
  INV_X1    g0604(.A(G137), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n805), .A2(new_n758), .B1(new_n760), .B2(new_n286), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT98), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G159), .A2(new_n739), .B1(new_n734), .B2(G143), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT34), .Z(new_n810));
  AOI211_X1 g0610(.A(new_n804), .B(new_n810), .C1(G50), .C2(new_n751), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n767), .A2(G87), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n769), .B2(new_n591), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n317), .B1(new_n745), .B2(new_n560), .C1(new_n735), .C2(new_n743), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n813), .B(new_n814), .C1(G311), .C2(new_n741), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n815), .B1(new_n376), .B2(new_n750), .C1(new_n731), .C2(new_n760), .ZN(new_n816));
  INV_X1    g0616(.A(new_n758), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n816), .B1(G303), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n727), .B1(new_n811), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n716), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n727), .A2(new_n724), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n820), .B1(new_n276), .B2(new_n821), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n819), .B(new_n822), .C1(new_n725), .C2(new_n788), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n800), .A2(new_n823), .ZN(G384));
  INV_X1    g0624(.A(KEYINPUT40), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n349), .A2(new_n646), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n363), .A2(new_n346), .A3(new_n348), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n350), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT37), .ZN(new_n829));
  INV_X1    g0629(.A(new_n826), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n830), .B1(new_n369), .B2(new_n354), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n829), .A2(new_n831), .A3(KEYINPUT38), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(KEYINPUT38), .B1(new_n829), .B2(new_n831), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  AND4_X1   g0636(.A1(new_n693), .A2(new_n610), .A3(new_n694), .A4(new_n647), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n788), .B1(new_n837), .B2(new_n685), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n442), .A2(new_n436), .ZN(new_n839));
  OR2_X1    g0639(.A1(new_n418), .A2(new_n434), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n436), .A2(new_n654), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n436), .B(new_n654), .C1(new_n435), .C2(new_n442), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n838), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n836), .B1(new_n844), .B2(KEYINPUT103), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT103), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n846), .B(new_n838), .C1(new_n842), .C2(new_n843), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n825), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(KEYINPUT101), .B1(new_n365), .B2(new_n368), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n366), .A2(new_n367), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n827), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT101), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n359), .A2(new_n363), .A3(new_n364), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n849), .A2(new_n635), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n830), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT38), .B1(new_n856), .B2(new_n829), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT102), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n833), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT38), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n852), .B1(new_n851), .B2(new_n853), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n861), .A2(new_n354), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n826), .B1(new_n862), .B2(new_n854), .ZN(new_n863));
  INV_X1    g0663(.A(new_n829), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n860), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT102), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n825), .B1(new_n859), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n844), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n848), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n399), .A2(new_n443), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n683), .A2(new_n684), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n870), .B1(new_n871), .B2(new_n687), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n869), .A2(new_n872), .ZN(new_n874));
  INV_X1    g0674(.A(G330), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT39), .B1(new_n859), .B2(new_n866), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n839), .A2(new_n654), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NOR3_X1   g0681(.A1(new_n877), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n786), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n789), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n842), .A2(new_n843), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n886), .A2(new_n835), .B1(new_n635), .B2(new_n646), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n705), .A2(new_n444), .A3(new_n708), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n640), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n888), .B(new_n890), .ZN(new_n891));
  OAI22_X1  g0691(.A1(new_n876), .A2(new_n891), .B1(new_n209), .B2(new_n712), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n891), .B2(new_n876), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT35), .ZN(new_n895));
  OAI211_X1 g0695(.A(G116), .B(new_n219), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n895), .B2(new_n894), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT36), .ZN(new_n898));
  OR3_X1    g0698(.A1(new_n216), .A2(new_n276), .A3(new_n336), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n201), .A2(G68), .ZN(new_n900));
  AOI211_X1 g0700(.A(new_n209), .B(G13), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  OR3_X1    g0701(.A1(new_n893), .A2(new_n898), .A3(new_n901), .ZN(G367));
  OAI221_X1 g0702(.A(new_n728), .B1(new_n213), .B2(new_n389), .C1(new_n239), .C2(new_n721), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n716), .A2(new_n903), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n739), .A2(new_n202), .B1(new_n741), .B2(G137), .ZN(new_n905));
  OAI221_X1 g0705(.A(new_n905), .B1(new_n330), .B2(new_n745), .C1(new_n286), .C2(new_n735), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(G58), .B2(new_n751), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n273), .B1(new_n733), .B2(new_n276), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT109), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n817), .A2(G143), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n761), .A2(G159), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n907), .A2(new_n909), .A3(new_n910), .A4(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n751), .A2(KEYINPUT46), .A3(G116), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT46), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n750), .B2(new_n591), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n745), .A2(new_n376), .B1(new_n733), .B2(new_n560), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n739), .B2(G283), .ZN(new_n917));
  INV_X1    g0717(.A(G317), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n317), .B1(new_n740), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n734), .B2(G303), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n913), .A2(new_n915), .A3(new_n917), .A4(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(G311), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n743), .A2(new_n760), .B1(new_n758), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n912), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  XOR2_X1   g0724(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n925));
  XNOR2_X1  g0725(.A(new_n924), .B(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n904), .B1(new_n926), .B2(new_n727), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n480), .A2(new_n647), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n697), .B(new_n928), .C1(new_n619), .C2(new_n491), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n929), .A2(KEYINPUT104), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(KEYINPUT104), .ZN(new_n931));
  INV_X1    g0731(.A(new_n928), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n930), .B(new_n931), .C1(new_n620), .C2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n927), .B1(new_n933), .B2(new_n779), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT105), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n935), .B(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n622), .A2(new_n654), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n572), .B(new_n579), .C1(new_n577), .C2(new_n647), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n660), .A2(new_n662), .A3(new_n940), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n941), .A2(KEYINPUT42), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n572), .B1(new_n939), .B2(new_n546), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n647), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n941), .A2(KEYINPUT42), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n942), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n946), .A2(KEYINPUT106), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(KEYINPUT106), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n947), .A2(new_n948), .B1(KEYINPUT43), .B2(new_n933), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n937), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n937), .A2(new_n949), .ZN(new_n952));
  INV_X1    g0752(.A(new_n940), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n951), .A2(new_n952), .B1(new_n661), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n952), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n661), .A2(new_n953), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n955), .A2(new_n956), .A3(new_n950), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT44), .ZN(new_n959));
  OR3_X1    g0759(.A1(new_n663), .A2(new_n959), .A3(new_n940), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n959), .B1(new_n663), .B2(new_n940), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n663), .A2(new_n940), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT45), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n663), .A2(KEYINPUT45), .A3(new_n940), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n962), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n661), .ZN(new_n969));
  OAI21_X1  g0769(.A(KEYINPUT108), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(KEYINPUT108), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n962), .A2(new_n967), .A3(new_n971), .A4(new_n661), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n652), .A2(KEYINPUT107), .ZN(new_n974));
  XOR2_X1   g0774(.A(new_n660), .B(new_n662), .Z(new_n975));
  XNOR2_X1  g0775(.A(new_n974), .B(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n968), .A2(new_n969), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n973), .A2(new_n709), .A3(new_n976), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n709), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n665), .B(KEYINPUT41), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n714), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n934), .B1(new_n958), .B2(new_n982), .ZN(G387));
  OAI22_X1  g0783(.A1(new_n717), .A2(new_n666), .B1(G107), .B2(new_n213), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n236), .A2(new_n252), .ZN(new_n985));
  INV_X1    g0785(.A(new_n666), .ZN(new_n986));
  AOI211_X1 g0786(.A(G45), .B(new_n986), .C1(G68), .C2(G77), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n284), .A2(G50), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT50), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n721), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n984), .B1(new_n985), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n766), .A2(new_n471), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n769), .B2(new_n330), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n273), .B1(new_n560), .B2(new_n733), .C1(new_n735), .C2(new_n423), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n993), .B(new_n994), .C1(G150), .C2(new_n741), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n276), .B2(new_n750), .C1(new_n284), .C2(new_n760), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(G159), .B2(new_n817), .ZN(new_n997));
  AOI22_X1  g0797(.A1(G303), .A2(new_n739), .B1(new_n734), .B2(G317), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n760), .B2(new_n922), .C1(new_n736), .C2(new_n758), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT48), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n999), .A2(new_n1000), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n750), .A2(new_n743), .B1(new_n731), .B2(new_n745), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT111), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT49), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n317), .B1(new_n733), .B2(new_n591), .C1(new_n753), .C2(new_n740), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n997), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n727), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n716), .B1(new_n729), .B2(new_n991), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1013), .A2(KEYINPUT112), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n660), .A2(new_n779), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1013), .A2(KEYINPUT112), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n1016), .A2(new_n1017), .B1(new_n714), .B2(new_n976), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n709), .A2(new_n976), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n711), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n709), .A2(new_n976), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1018), .B1(new_n1020), .B2(new_n1021), .ZN(G393));
  INV_X1    g0822(.A(G159), .ZN(new_n1023));
  OAI22_X1  g0823(.A1(new_n758), .A2(new_n286), .B1(new_n1023), .B2(new_n735), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT51), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n284), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n761), .A2(new_n202), .B1(new_n1026), .B2(new_n739), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1027), .A2(KEYINPUT115), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(KEYINPUT115), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n766), .A2(G77), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n741), .A2(G143), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1030), .A2(new_n1031), .A3(new_n273), .A4(new_n812), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G68), .B2(new_n751), .ZN(new_n1033));
  NAND4_X1  g0833(.A1(new_n1025), .A2(new_n1028), .A3(new_n1029), .A4(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(KEYINPUT116), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n758), .A2(new_n918), .B1(new_n922), .B2(new_n735), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT52), .Z(new_n1037));
  NAND2_X1  g0837(.A1(new_n739), .A2(G294), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n273), .B1(new_n767), .B2(G107), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G116), .A2(new_n766), .B1(new_n741), .B2(G322), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1038), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(G283), .B2(new_n751), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n583), .B2(new_n760), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1035), .B1(new_n1037), .B2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1034), .A2(KEYINPUT116), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n727), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n953), .A2(new_n726), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n728), .B1(new_n560), .B2(new_n213), .C1(new_n246), .C2(new_n721), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1046), .A2(new_n716), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n977), .A2(KEYINPUT113), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT113), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n968), .A2(new_n1052), .A3(new_n969), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n973), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1055), .A2(KEYINPUT114), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n713), .B1(new_n1055), .B2(KEYINPUT114), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1050), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1055), .A2(new_n1019), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1059), .A2(new_n711), .A3(new_n978), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT117), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1058), .A2(KEYINPUT117), .A3(new_n1060), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1063), .A2(new_n1064), .ZN(G390));
  OAI21_X1  g0865(.A(G330), .B1(new_n837), .B2(new_n685), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n791), .B1(new_n1066), .B2(KEYINPUT119), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n875), .B1(new_n871), .B2(new_n687), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT119), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n885), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n689), .A2(G330), .A3(new_n788), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n1073), .A2(KEYINPUT120), .B1(new_n1074), .B2(new_n885), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n885), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT120), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n702), .A2(new_n703), .A3(new_n883), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n787), .A2(new_n394), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1076), .A2(new_n1077), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1075), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n844), .A2(G330), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n1074), .B2(new_n885), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(new_n884), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n444), .A2(KEYINPUT118), .A3(new_n1068), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT118), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n870), .B2(new_n1066), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1089), .A2(new_n640), .A3(new_n889), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1085), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1078), .A2(new_n1079), .A3(new_n885), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n880), .B1(new_n859), .B2(new_n866), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1074), .A2(new_n885), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n789), .A2(new_n883), .B1(new_n842), .B2(new_n843), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n877), .A2(new_n879), .B1(new_n1097), .B2(new_n880), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1095), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT39), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n832), .B1(new_n865), .B2(KEYINPUT102), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n857), .A2(new_n858), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1100), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n878), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n886), .A2(new_n881), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n1104), .A2(new_n1105), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1099), .B1(new_n1106), .B2(new_n1082), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n665), .B1(new_n1092), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1108), .B1(new_n1092), .B2(new_n1107), .ZN(new_n1109));
  OR2_X1    g0909(.A1(new_n1107), .A2(new_n713), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT121), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n821), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n716), .B1(new_n1026), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1030), .B1(new_n743), .B2(new_n740), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n317), .B1(new_n330), .B2(new_n733), .C1(new_n735), .C2(new_n591), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n1114), .B(new_n1115), .C1(G97), .C2(new_n739), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n1116), .B1(new_n318), .B2(new_n750), .C1(new_n731), .C2(new_n758), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n760), .A2(new_n376), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n735), .A2(new_n803), .ZN(new_n1119));
  XOR2_X1   g0919(.A(KEYINPUT54), .B(G143), .Z(new_n1120));
  AOI211_X1 g0920(.A(new_n317), .B(new_n1119), .C1(new_n739), .C2(new_n1120), .ZN(new_n1121));
  OR3_X1    g0921(.A1(new_n750), .A2(KEYINPUT53), .A3(new_n286), .ZN(new_n1122));
  OAI21_X1  g0922(.A(KEYINPUT53), .B1(new_n750), .B2(new_n286), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n745), .A2(new_n1023), .B1(new_n733), .B2(new_n201), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(G125), .B2(new_n741), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(G128), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n1127), .A2(new_n758), .B1(new_n760), .B2(new_n805), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n1117), .A2(new_n1118), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1113), .B1(new_n1129), .B2(new_n727), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1104), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1130), .B1(new_n1131), .B2(new_n725), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1110), .A2(new_n1111), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1111), .B1(new_n1110), .B2(new_n1132), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1109), .B1(new_n1133), .B2(new_n1134), .ZN(G378));
  INV_X1    g0935(.A(new_n888), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n875), .B1(new_n867), .B2(new_n844), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n308), .A2(new_n297), .A3(new_n646), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n297), .A2(new_n646), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n301), .A2(new_n307), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1141), .B(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n848), .A2(new_n1137), .A3(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1144), .B1(new_n848), .B2(new_n1137), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1136), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n838), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n885), .A2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n835), .B1(new_n1149), .B2(new_n846), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n844), .A2(KEYINPUT103), .ZN(new_n1151));
  AOI21_X1  g0951(.A(KEYINPUT40), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n868), .A2(G330), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1143), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n848), .A2(new_n1144), .A3(new_n1137), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1154), .A2(new_n888), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n713), .B1(new_n1147), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT122), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1143), .A2(new_n724), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n715), .B1(new_n202), .B2(new_n1112), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n317), .A2(new_n516), .ZN(new_n1162));
  AOI211_X1 g0962(.A(G50), .B(new_n1162), .C1(new_n270), .C2(new_n248), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1162), .B1(new_n745), .B2(new_n330), .C1(new_n735), .C2(new_n376), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n739), .A2(new_n471), .B1(new_n741), .B2(G283), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n335), .B2(new_n733), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1164), .B(new_n1166), .C1(G77), .C2(new_n751), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1167), .B1(new_n560), .B2(new_n760), .C1(new_n591), .C2(new_n758), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT58), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1163), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n739), .A2(G137), .B1(G150), .B2(new_n766), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n735), .B2(new_n1127), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n751), .B2(new_n1120), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n817), .A2(G125), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1173), .B(new_n1174), .C1(new_n803), .C2(new_n760), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n270), .B(new_n248), .C1(new_n733), .C2(new_n1023), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G124), .B2(new_n741), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1170), .B1(new_n1169), .B2(new_n1168), .C1(new_n1176), .C2(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1161), .B1(new_n1181), .B2(new_n727), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1160), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1158), .A2(new_n1159), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1183), .ZN(new_n1185));
  OAI21_X1  g0985(.A(KEYINPUT122), .B1(new_n1157), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1147), .A2(new_n1156), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1075), .A2(new_n1080), .B1(new_n1083), .B2(new_n884), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1091), .B1(new_n1107), .B2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1188), .A2(KEYINPUT57), .A3(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1191), .A2(KEYINPUT123), .A3(new_n711), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT57), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1192), .A2(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT123), .B1(new_n1191), .B2(new_n711), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1187), .B1(new_n1196), .B2(new_n1197), .ZN(G375));
  NAND2_X1  g0998(.A1(new_n1189), .A2(new_n1090), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1092), .A2(new_n981), .A3(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n716), .B1(G68), .B2(new_n1112), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n992), .B1(new_n583), .B2(new_n740), .C1(new_n769), .C2(new_n376), .ZN(new_n1202));
  OAI221_X1 g1002(.A(new_n317), .B1(new_n276), .B2(new_n733), .C1(new_n735), .C2(new_n731), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1202), .B(new_n1203), .C1(G97), .C2(new_n751), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n591), .B2(new_n760), .C1(new_n743), .C2(new_n758), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n769), .A2(new_n286), .B1(new_n745), .B2(new_n423), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n273), .B1(new_n335), .B2(new_n733), .C1(new_n735), .C2(new_n805), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(G128), .C2(new_n741), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n761), .A2(new_n1120), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n817), .A2(G132), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n751), .A2(G159), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(KEYINPUT124), .B1(new_n1205), .B2(new_n1212), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1213), .A2(new_n1012), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1205), .A2(KEYINPUT124), .A3(new_n1212), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1201), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n725), .B2(new_n885), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n1189), .B2(new_n713), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1200), .A2(new_n1219), .ZN(G381));
  NOR4_X1   g1020(.A1(G381), .A2(G384), .A3(G396), .A4(G393), .ZN(new_n1221));
  INV_X1    g1021(.A(G387), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1110), .A2(new_n1132), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1109), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  OR4_X1    g1026(.A1(G390), .A2(G375), .A3(new_n1223), .A4(new_n1226), .ZN(G407));
  INV_X1    g1027(.A(G343), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(G213), .ZN(new_n1229));
  OR3_X1    g1029(.A1(G375), .A2(new_n1226), .A3(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(G407), .A2(new_n1230), .A3(G213), .ZN(G409));
  INV_X1    g1031(.A(new_n1064), .ZN(new_n1232));
  AOI21_X1  g1032(.A(KEYINPUT117), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1222), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  XOR2_X1   g1034(.A(G393), .B(G396), .Z(new_n1235));
  NAND3_X1  g1035(.A1(new_n1063), .A2(G387), .A3(new_n1064), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1235), .B1(new_n1234), .B2(new_n1236), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT127), .ZN(new_n1241));
  OAI211_X1 g1041(.A(G378), .B(new_n1187), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1158), .A2(new_n1183), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1193), .A2(new_n980), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1225), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1229), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1189), .A2(KEYINPUT60), .A3(new_n1090), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n711), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1092), .A2(KEYINPUT60), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1249), .B1(new_n1250), .B2(new_n1199), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1251), .A2(new_n1218), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1228), .A2(G213), .A3(G2897), .ZN(new_n1256));
  XOR2_X1   g1056(.A(new_n1256), .B(KEYINPUT126), .Z(new_n1257));
  INV_X1    g1057(.A(KEYINPUT125), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n800), .B2(new_n823), .ZN(new_n1259));
  OAI22_X1  g1059(.A1(new_n1253), .A2(new_n1259), .B1(new_n1251), .B2(new_n1218), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1255), .A2(new_n1257), .A3(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1257), .B1(new_n1255), .B2(new_n1260), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1247), .A2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT61), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1241), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1255), .A2(new_n1260), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1246), .A2(new_n1229), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT62), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n1242), .A2(new_n1245), .B1(G213), .B2(new_n1228), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT62), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1271), .A2(new_n1272), .A3(new_n1268), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1240), .B1(new_n1266), .B2(new_n1274), .ZN(new_n1275));
  AND4_X1   g1075(.A1(KEYINPUT63), .A2(new_n1246), .A3(new_n1229), .A4(new_n1268), .ZN(new_n1276));
  AOI21_X1  g1076(.A(KEYINPUT63), .B1(new_n1271), .B2(new_n1268), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1239), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(KEYINPUT127), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1262), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1255), .A2(new_n1257), .A3(new_n1260), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1280), .A2(new_n1281), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1279), .B(new_n1265), .C1(new_n1282), .C2(new_n1271), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1278), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1275), .A2(new_n1285), .ZN(G405));
  NAND2_X1  g1086(.A1(G375), .A2(new_n1225), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1242), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1268), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1287), .A2(new_n1242), .A3(new_n1267), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(new_n1240), .ZN(G402));
endmodule


