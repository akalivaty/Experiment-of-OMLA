//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G122), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XOR2_X1   g004(.A(KEYINPUT2), .B(G113), .Z(new_n191));
  XNOR2_X1  g005(.A(G116), .B(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT2), .B(G113), .ZN(new_n194));
  INV_X1    g008(.A(G116), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G119), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G116), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n194), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n193), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  INV_X1    g015(.A(G104), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT3), .B1(new_n202), .B2(G107), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT83), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT83), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n205), .B(KEYINPUT3), .C1(new_n202), .C2(G107), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G107), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT84), .B1(new_n208), .B2(G104), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT84), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(new_n202), .A3(G107), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n202), .A2(G107), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT3), .ZN(new_n213));
  AOI22_X1  g027(.A1(new_n209), .A2(new_n211), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n201), .B1(new_n207), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT4), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n200), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT85), .ZN(new_n218));
  INV_X1    g032(.A(new_n206), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n208), .A2(G104), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n205), .B1(new_n220), .B2(KEYINPUT3), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n209), .A2(new_n211), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n212), .A2(new_n213), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n218), .B(G101), .C1(new_n222), .C2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n207), .A2(new_n201), .A3(new_n214), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n226), .A2(KEYINPUT4), .A3(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n215), .A2(new_n218), .ZN(new_n229));
  OAI211_X1 g043(.A(KEYINPUT86), .B(new_n217), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n192), .A2(KEYINPUT5), .ZN(new_n231));
  INV_X1    g045(.A(G113), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT5), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n232), .B1(new_n196), .B2(new_n233), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n231), .A2(new_n234), .B1(new_n191), .B2(new_n192), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n208), .A2(G104), .ZN(new_n236));
  OAI21_X1  g050(.A(G101), .B1(new_n212), .B2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n227), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n230), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(G101), .B1(new_n222), .B2(new_n225), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(KEYINPUT85), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n241), .A2(KEYINPUT4), .A3(new_n226), .A4(new_n227), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT86), .B1(new_n242), .B2(new_n217), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n190), .B1(new_n239), .B2(new_n243), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n217), .B1(new_n228), .B2(new_n229), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT86), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n247), .A2(new_n189), .A3(new_n238), .A4(new_n230), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n244), .A2(KEYINPUT6), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G953), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G224), .ZN(new_n251));
  INV_X1    g065(.A(G146), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G143), .ZN(new_n253));
  INV_X1    g067(.A(G143), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G146), .ZN(new_n255));
  AND2_X1   g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  OR2_X1    g071(.A1(KEYINPUT75), .A2(G125), .ZN(new_n258));
  NAND2_X1  g072(.A1(KEYINPUT75), .A2(G125), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT64), .B1(new_n252), .B2(G143), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT64), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n262), .A2(new_n254), .A3(G146), .ZN(new_n263));
  AOI22_X1  g077(.A1(new_n261), .A2(new_n263), .B1(G143), .B2(new_n252), .ZN(new_n264));
  NOR2_X1   g078(.A1(KEYINPUT0), .A2(G128), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n256), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n257), .B(new_n260), .C1(new_n264), .C2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n269));
  AND4_X1   g083(.A1(new_n269), .A2(new_n253), .A3(new_n255), .A4(G128), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n262), .B1(new_n254), .B2(G146), .ZN(new_n271));
  NOR3_X1   g085(.A1(new_n252), .A2(KEYINPUT64), .A3(G143), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n253), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G128), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT66), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT66), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G128), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n253), .A2(KEYINPUT1), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n270), .B1(new_n273), .B2(new_n280), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n251), .B(new_n268), .C1(new_n281), .C2(new_n260), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n260), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n261), .A2(new_n263), .ZN(new_n285));
  AOI22_X1  g099(.A1(new_n285), .A2(new_n253), .B1(new_n278), .B2(new_n279), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n284), .B1(new_n286), .B2(new_n270), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n251), .B1(new_n287), .B2(new_n268), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT6), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n290), .B(new_n190), .C1(new_n239), .C2(new_n243), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n249), .A2(new_n289), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT7), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n251), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n294), .B1(new_n283), .B2(new_n288), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n287), .A2(new_n268), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(new_n293), .A3(new_n251), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT87), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n238), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n227), .A2(new_n237), .ZN(new_n300));
  INV_X1    g114(.A(new_n235), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n227), .A2(new_n235), .A3(KEYINPUT87), .A4(new_n237), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n299), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n189), .B(KEYINPUT8), .ZN(new_n305));
  AOI22_X1  g119(.A1(new_n295), .A2(new_n297), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n248), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G902), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT88), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT88), .ZN(new_n310));
  AOI211_X1 g124(.A(new_n310), .B(G902), .C1(new_n248), .C2(new_n306), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n292), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(G210), .B1(G237), .B2(G902), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT89), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n312), .A2(new_n316), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n292), .B(new_n315), .C1(new_n309), .C2(new_n311), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n188), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT9), .B(G234), .ZN(new_n320));
  OAI21_X1  g134(.A(G221), .B1(new_n320), .B2(G902), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G469), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(new_n308), .ZN(new_n324));
  INV_X1    g138(.A(new_n257), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(new_n273), .B2(new_n266), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n215), .A2(new_n216), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n326), .B(new_n327), .C1(new_n228), .C2(new_n229), .ZN(new_n328));
  INV_X1    g142(.A(G137), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(G134), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT65), .ZN(new_n331));
  INV_X1    g145(.A(G134), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n331), .B1(new_n332), .B2(G137), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n330), .B1(new_n333), .B2(KEYINPUT11), .ZN(new_n334));
  INV_X1    g148(.A(G131), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT11), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n331), .B(new_n336), .C1(new_n332), .C2(G137), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n335), .B1(new_n334), .B2(new_n337), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n300), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT10), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n281), .A2(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n253), .A2(new_n255), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n274), .B1(new_n253), .B2(KEYINPUT1), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n227), .B(new_n237), .C1(new_n270), .C2(new_n346), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n341), .A2(new_n343), .B1(new_n347), .B2(new_n342), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n328), .A2(new_n340), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n250), .A2(KEYINPUT69), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT69), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G953), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G227), .ZN(new_n354));
  XOR2_X1   g168(.A(G110), .B(G140), .Z(new_n355));
  XNOR2_X1  g169(.A(new_n354), .B(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n349), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n340), .B1(new_n328), .B2(new_n348), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n300), .A2(new_n281), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n340), .B1(new_n362), .B2(new_n347), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n363), .A2(KEYINPUT12), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n363), .A2(KEYINPUT12), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n349), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n359), .A2(new_n361), .B1(new_n366), .B2(new_n356), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n324), .B1(new_n367), .B2(G469), .ZN(new_n368));
  XOR2_X1   g182(.A(KEYINPUT73), .B(G902), .Z(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n349), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n356), .B1(new_n371), .B2(new_n360), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n349), .B(new_n357), .C1(new_n364), .C2(new_n365), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n370), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n323), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n322), .B1(new_n368), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n319), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT20), .ZN(new_n378));
  XNOR2_X1  g192(.A(G113), .B(G122), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n379), .B(new_n202), .ZN(new_n380));
  INV_X1    g194(.A(G237), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n254), .A2(KEYINPUT90), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n353), .A2(G214), .A3(new_n381), .A4(new_n382), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n350), .A2(new_n352), .A3(G214), .A4(new_n381), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(KEYINPUT90), .A3(new_n254), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n386), .A2(KEYINPUT18), .A3(G131), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT18), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n383), .B(new_n385), .C1(new_n388), .C2(new_n335), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n260), .A2(G140), .ZN(new_n390));
  NOR2_X1   g204(.A1(G125), .A2(G140), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(G146), .A3(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G125), .B(G140), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n252), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n393), .A2(KEYINPUT91), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT91), .B1(new_n393), .B2(new_n395), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n387), .B(new_n389), .C1(new_n396), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n386), .A2(G131), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT17), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n383), .A2(new_n385), .A3(new_n335), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n335), .B1(new_n383), .B2(new_n385), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT17), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G140), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n406), .B1(new_n258), .B2(new_n259), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT16), .B1(new_n407), .B2(new_n391), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT16), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n260), .A2(new_n409), .A3(new_n406), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(G146), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT76), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n408), .A2(KEYINPUT76), .A3(G146), .A4(new_n410), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n408), .A2(new_n410), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n252), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n413), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  OAI211_X1 g231(.A(new_n380), .B(new_n398), .C1(new_n405), .C2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n391), .B1(new_n260), .B2(G140), .ZN(new_n419));
  XOR2_X1   g233(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n420));
  AOI22_X1  g234(.A1(new_n419), .A2(KEYINPUT19), .B1(new_n394), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(new_n252), .ZN(new_n422));
  INV_X1    g236(.A(new_n401), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n422), .B(new_n411), .C1(new_n423), .C2(new_n403), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n398), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n380), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n418), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g242(.A1(G475), .A2(G902), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n378), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n429), .ZN(new_n431));
  AOI211_X1 g245(.A(KEYINPUT20), .B(new_n431), .C1(new_n418), .C2(new_n427), .ZN(new_n432));
  AOI21_X1  g246(.A(G146), .B1(new_n408), .B2(new_n410), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n433), .B1(new_n412), .B2(new_n411), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n434), .A2(new_n402), .A3(new_n414), .A4(new_n404), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n398), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n426), .ZN(new_n437));
  AOI21_X1  g251(.A(G902), .B1(new_n437), .B2(new_n418), .ZN(new_n438));
  INV_X1    g252(.A(G475), .ZN(new_n439));
  OAI22_X1  g253(.A1(new_n430), .A2(new_n432), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G217), .ZN(new_n441));
  NOR3_X1   g255(.A1(new_n320), .A2(new_n441), .A3(G953), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(KEYINPUT94), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(G116), .B(G122), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT14), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n195), .A2(KEYINPUT14), .A3(G122), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(G107), .A3(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT93), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n445), .A2(new_n208), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT66), .B(G128), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G143), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n254), .A2(G128), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n455), .A2(G134), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n332), .B1(new_n453), .B2(new_n454), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n450), .B(new_n451), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  XOR2_X1   g272(.A(new_n454), .B(KEYINPUT13), .Z(new_n459));
  INV_X1    g273(.A(new_n453), .ZN(new_n460));
  OAI21_X1  g274(.A(G134), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n445), .B(new_n208), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n461), .B(new_n462), .C1(G134), .C2(new_n455), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n444), .B1(new_n458), .B2(new_n463), .ZN(new_n464));
  XOR2_X1   g278(.A(new_n449), .B(KEYINPUT93), .Z(new_n465));
  OAI21_X1  g279(.A(new_n451), .B1(new_n456), .B2(new_n457), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n463), .B(new_n444), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n369), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(G478), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(KEYINPUT15), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n469), .B(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n440), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n353), .ZN(new_n474));
  NAND2_X1  g288(.A1(G234), .A2(G237), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n474), .A2(new_n370), .A3(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT21), .B(G898), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n475), .A2(G952), .A3(new_n250), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n473), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n377), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(G472), .A2(G902), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n484), .B(KEYINPUT72), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT32), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n200), .ZN(new_n488));
  INV_X1    g302(.A(new_n281), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT68), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n332), .A2(G137), .ZN(new_n492));
  OAI21_X1  g306(.A(G131), .B1(new_n492), .B2(new_n330), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n489), .A2(new_n490), .A3(new_n491), .A4(new_n493), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n491), .B(new_n493), .C1(new_n286), .C2(new_n270), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(KEYINPUT68), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n326), .B1(new_n338), .B2(new_n339), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n494), .A2(KEYINPUT30), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT67), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n495), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT30), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AOI211_X1 g316(.A(KEYINPUT67), .B(KEYINPUT30), .C1(new_n497), .C2(new_n495), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n488), .B(new_n498), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n494), .A2(new_n200), .A3(new_n496), .A4(new_n497), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n353), .A2(G210), .A3(new_n381), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n506), .B(KEYINPUT27), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT26), .B(G101), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n507), .B(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n504), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT31), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT70), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n510), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n200), .B1(new_n497), .B2(new_n495), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT28), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n497), .A2(new_n200), .A3(new_n495), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n518), .B1(new_n516), .B2(new_n505), .ZN(new_n519));
  INV_X1    g333(.A(new_n509), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n513), .A2(new_n514), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT31), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n504), .A2(new_n523), .A3(new_n505), .A4(new_n509), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n524), .B(KEYINPUT71), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n487), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT29), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n518), .B(new_n527), .C1(new_n516), .C2(new_n505), .ZN(new_n528));
  AND2_X1   g342(.A1(new_n528), .A2(new_n509), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n496), .A2(new_n494), .A3(new_n497), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n488), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n516), .B1(new_n531), .B2(new_n505), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n517), .A2(new_n516), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT29), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n370), .B1(new_n529), .B2(new_n535), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n504), .A2(new_n505), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(new_n527), .A3(new_n520), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(G472), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n514), .A2(new_n521), .ZN(new_n541));
  AOI21_X1  g355(.A(KEYINPUT70), .B1(new_n510), .B2(KEYINPUT31), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT71), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n524), .B(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n485), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n526), .B(new_n540), .C1(new_n546), .C2(KEYINPUT32), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n441), .B1(new_n369), .B2(G234), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT74), .B1(new_n197), .B2(G128), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n278), .B2(new_n197), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT24), .B(G110), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n452), .A2(KEYINPUT74), .A3(G119), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n452), .A2(KEYINPUT23), .A3(G119), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT23), .B1(new_n274), .B2(G119), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(new_n197), .B2(G128), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT77), .B(G110), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n554), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n559), .A2(new_n411), .A3(new_n395), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT78), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n559), .A2(KEYINPUT78), .A3(new_n411), .A4(new_n395), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n550), .A2(new_n552), .ZN(new_n565));
  INV_X1    g379(.A(new_n551), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n554), .A2(new_n556), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(G110), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n570), .B1(new_n434), .B2(new_n414), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT79), .B1(new_n564), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n570), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n417), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT79), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n574), .A2(new_n575), .A3(new_n562), .A4(new_n563), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n353), .A2(G221), .A3(G234), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT22), .B(G137), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n572), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n574), .A2(new_n562), .A3(new_n563), .A4(new_n579), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT80), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n572), .A2(KEYINPUT80), .A3(new_n576), .A4(new_n580), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT25), .B1(new_n587), .B2(new_n369), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT25), .ZN(new_n589));
  AOI211_X1 g403(.A(new_n589), .B(new_n370), .C1(new_n585), .C2(new_n586), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n548), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n548), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n308), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT81), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n587), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n547), .A2(new_n596), .A3(KEYINPUT82), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(KEYINPUT82), .B1(new_n547), .B2(new_n596), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n483), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G101), .ZN(G3));
  NAND2_X1  g415(.A1(new_n312), .A2(new_n313), .ZN(new_n602));
  OAI211_X1 g416(.A(new_n292), .B(new_n314), .C1(new_n309), .C2(new_n311), .ZN(new_n603));
  AND4_X1   g417(.A1(KEYINPUT95), .A2(new_n602), .A3(new_n187), .A4(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n188), .B1(new_n312), .B2(new_n313), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT95), .B1(new_n605), .B2(new_n603), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT96), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n607), .B1(new_n608), .B2(new_n443), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  OAI22_X1  g424(.A1(new_n609), .A2(new_n610), .B1(new_n464), .B2(new_n468), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n608), .A2(new_n443), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n612), .A2(new_n607), .A3(KEYINPUT33), .A4(new_n467), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n611), .A2(G478), .A3(new_n369), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n469), .A2(new_n470), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n440), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n481), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n604), .A2(new_n606), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n485), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n621), .B1(new_n522), .B2(new_n525), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n370), .B1(new_n543), .B2(new_n545), .ZN(new_n623));
  INV_X1    g437(.A(G472), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n591), .A2(new_n595), .A3(new_n376), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n620), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT34), .B(G104), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  NAND3_X1  g444(.A1(new_n602), .A2(new_n187), .A3(new_n603), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT95), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n605), .A2(KEYINPUT95), .A3(new_n603), .ZN(new_n634));
  INV_X1    g448(.A(new_n471), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n469), .B(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n440), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n481), .B(KEYINPUT97), .ZN(new_n638));
  AND4_X1   g452(.A1(new_n633), .A2(new_n634), .A3(new_n637), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n627), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G107), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  OAI21_X1  g456(.A(new_n369), .B1(new_n522), .B2(new_n525), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n546), .B1(G472), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n572), .A2(new_n576), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n580), .A2(KEYINPUT36), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n645), .B(new_n646), .Z(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n594), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n482), .B1(new_n591), .B2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n644), .A2(new_n649), .A3(new_n319), .A4(new_n376), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT37), .B(G110), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G12));
  NOR2_X1   g466(.A1(new_n604), .A2(new_n606), .ZN(new_n653));
  INV_X1    g467(.A(new_n376), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n624), .B1(new_n536), .B2(new_n538), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n543), .A2(new_n545), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n655), .B1(new_n656), .B2(new_n487), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n622), .A2(new_n486), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n654), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n591), .A2(new_n648), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n428), .A2(new_n429), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n661), .A2(KEYINPUT20), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n428), .A2(new_n378), .A3(new_n429), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n437), .A2(new_n418), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n308), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(G475), .ZN(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n476), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n480), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n472), .A2(new_n664), .A3(new_n667), .A4(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT98), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n653), .A2(new_n659), .A3(new_n660), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G128), .ZN(G30));
  XOR2_X1   g489(.A(KEYINPUT100), .B(KEYINPUT40), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n670), .B(KEYINPUT39), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n676), .B1(new_n654), .B2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n676), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n376), .A2(new_n677), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n587), .A2(new_n369), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n589), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n587), .A2(KEYINPUT25), .A3(new_n369), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n592), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n648), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n440), .A2(new_n472), .ZN(new_n688));
  NOR4_X1   g502(.A1(new_n686), .A2(new_n687), .A3(new_n188), .A4(new_n688), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n682), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT101), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n537), .A2(new_n520), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n520), .A2(new_n531), .A3(new_n505), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n308), .ZN(new_n694));
  OAI21_X1  g508(.A(G472), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT99), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n658), .A2(new_n697), .A3(new_n526), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n317), .A2(new_n318), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT38), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n690), .A2(new_n691), .A3(new_n698), .A4(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n700), .A2(new_n682), .A3(new_n689), .A4(new_n698), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(KEYINPUT101), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n254), .ZN(G45));
  NAND2_X1  g519(.A1(new_n618), .A2(new_n670), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n653), .A2(new_n659), .A3(new_n660), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  OR2_X1    g523(.A1(new_n374), .A2(new_n323), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n710), .A2(new_n321), .A3(new_n375), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n547), .A2(new_n596), .A3(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n633), .A2(new_n481), .A3(new_n634), .A4(new_n618), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT41), .B(G113), .Z(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G15));
  NAND4_X1  g531(.A1(new_n633), .A2(new_n634), .A3(new_n637), .A4(new_n638), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(new_n195), .ZN(G18));
  NOR3_X1   g534(.A1(new_n604), .A2(new_n606), .A3(new_n711), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n721), .A2(KEYINPUT102), .A3(new_n547), .A4(new_n649), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT102), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n547), .A2(new_n649), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n633), .A2(new_n634), .A3(new_n712), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  NOR2_X1   g542(.A1(new_n711), .A2(new_n688), .ZN(new_n729));
  AND4_X1   g543(.A1(new_n633), .A2(new_n634), .A3(new_n638), .A4(new_n729), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n532), .A2(new_n534), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n520), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n545), .A2(new_n511), .A3(new_n732), .ZN(new_n733));
  AOI22_X1  g547(.A1(new_n643), .A2(G472), .B1(new_n621), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n596), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT103), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n730), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n633), .A2(new_n634), .A3(new_n638), .A4(new_n729), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n596), .A2(new_n734), .ZN(new_n739));
  OAI21_X1  g553(.A(KEYINPUT103), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G122), .ZN(G24));
  AND3_X1   g556(.A1(new_n734), .A2(new_n660), .A3(new_n707), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n721), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G125), .ZN(G27));
  NAND3_X1  g559(.A1(new_n317), .A2(new_n187), .A3(new_n318), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT42), .ZN(new_n747));
  NOR4_X1   g561(.A1(new_n706), .A2(new_n746), .A3(new_n654), .A4(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT104), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n658), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(KEYINPUT32), .B1(new_n656), .B2(new_n621), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n657), .B1(new_n751), .B2(KEYINPUT104), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n748), .B(new_n596), .C1(new_n750), .C2(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n746), .A2(new_n654), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n547), .A2(new_n596), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n747), .B1(new_n755), .B2(new_n706), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G131), .ZN(G33));
  NAND4_X1  g572(.A1(new_n547), .A2(new_n596), .A3(new_n754), .A4(new_n673), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G134), .ZN(G36));
  AOI21_X1  g574(.A(new_n440), .B1(new_n615), .B2(new_n614), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT106), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n762), .B1(new_n440), .B2(new_n763), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n761), .A2(new_n764), .ZN(new_n766));
  AOI22_X1  g580(.A1(new_n765), .A2(new_n766), .B1(new_n591), .B2(new_n648), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(KEYINPUT44), .A3(new_n625), .ZN(new_n768));
  INV_X1    g582(.A(new_n746), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT107), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n366), .A2(new_n356), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n772), .B1(new_n360), .B2(new_n358), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n367), .A2(KEYINPUT45), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n776), .A3(G469), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT105), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n775), .A2(new_n776), .A3(KEYINPUT105), .A4(G469), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n324), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT46), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n375), .B1(new_n781), .B2(KEYINPUT46), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n321), .B(new_n677), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT107), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n768), .A2(new_n787), .A3(new_n769), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT44), .B1(new_n767), .B2(new_n625), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n771), .A2(new_n786), .A3(new_n788), .A4(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G137), .ZN(G39));
  NOR4_X1   g606(.A1(new_n547), .A2(new_n596), .A3(new_n706), .A4(new_n746), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n781), .A2(KEYINPUT46), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n375), .A3(new_n782), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT47), .B1(new_n795), .B2(new_n321), .ZN(new_n796));
  OAI211_X1 g610(.A(KEYINPUT47), .B(new_n321), .C1(new_n783), .C2(new_n784), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n793), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G140), .ZN(G42));
  AND4_X1   g614(.A1(new_n591), .A2(new_n648), .A3(new_n376), .A4(new_n670), .ZN(new_n801));
  INV_X1    g615(.A(new_n688), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n653), .A2(new_n698), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n744), .A2(new_n674), .A3(new_n708), .A4(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n727), .A2(new_n600), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n547), .A2(new_n596), .A3(new_n712), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n808), .B1(new_n639), .B2(new_n620), .ZN(new_n809));
  INV_X1    g623(.A(new_n482), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n810), .B1(new_n686), .B2(new_n687), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n377), .ZN(new_n812));
  OAI21_X1  g626(.A(KEYINPUT109), .B1(new_n440), .B2(new_n636), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT109), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n472), .A2(new_n664), .A3(new_n667), .A4(new_n814), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n813), .A2(new_n815), .A3(new_n638), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n816), .A2(new_n319), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n812), .A2(new_n644), .B1(new_n627), .B2(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n616), .A2(new_n440), .A3(new_n638), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n699), .A2(new_n187), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT108), .ZN(new_n821));
  INV_X1    g635(.A(new_n626), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT108), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n319), .A2(new_n823), .A3(new_n819), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n821), .A2(new_n644), .A3(new_n822), .A4(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n809), .A2(new_n818), .A3(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n736), .B1(new_n730), .B2(new_n735), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n738), .A2(new_n739), .A3(KEYINPUT103), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n807), .A2(new_n826), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n473), .A2(new_n670), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n831), .B1(new_n591), .B2(new_n648), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n547), .A2(new_n832), .A3(new_n376), .A4(new_n769), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n754), .A2(new_n734), .A3(new_n660), .A4(new_n707), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n759), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n753), .B2(new_n756), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n806), .A2(new_n830), .A3(KEYINPUT53), .A4(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT111), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n599), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n597), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n841), .A2(new_n483), .B1(new_n722), .B2(new_n726), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n822), .A2(new_n644), .A3(new_n319), .A4(new_n816), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n825), .A2(new_n650), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n713), .B1(new_n714), .B2(new_n718), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n842), .A2(new_n836), .A3(new_n846), .A4(new_n741), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n633), .A2(new_n634), .A3(new_n660), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n526), .A2(new_n540), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n376), .B1(new_n751), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n851), .A2(new_n673), .B1(new_n721), .B2(new_n743), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n852), .A2(new_n805), .A3(new_n708), .A4(new_n803), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n804), .A2(KEYINPUT52), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n847), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n856), .A2(KEYINPUT111), .A3(KEYINPUT53), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n807), .A2(new_n826), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT110), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n858), .A2(new_n859), .A3(new_n741), .A4(new_n836), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n847), .A2(KEYINPUT110), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n744), .A2(new_n674), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(KEYINPUT52), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n853), .A2(new_n854), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n860), .A2(new_n861), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n839), .A2(new_n857), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT112), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n752), .A2(new_n750), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n591), .A2(new_n595), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n765), .A2(new_n766), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n769), .A2(new_n712), .A3(new_n479), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT48), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(KEYINPUT116), .A3(new_n878), .ZN(new_n879));
  XNOR2_X1  g693(.A(KEYINPUT116), .B(KEYINPUT48), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n873), .A2(new_n876), .A3(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n874), .A2(new_n739), .A3(new_n480), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n721), .ZN(new_n883));
  INV_X1    g697(.A(G952), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n875), .A2(new_n698), .A3(new_n872), .ZN(new_n885));
  AOI211_X1 g699(.A(new_n884), .B(G953), .C1(new_n885), .C2(new_n618), .ZN(new_n886));
  AND4_X1   g700(.A1(new_n879), .A2(new_n881), .A3(new_n883), .A4(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n616), .A2(new_n440), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n734), .A2(new_n660), .ZN(new_n889));
  AOI22_X1  g703(.A1(new_n885), .A2(new_n888), .B1(new_n876), .B2(new_n889), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n700), .A2(new_n187), .A3(new_n711), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT113), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT50), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT114), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n892), .A2(new_n894), .A3(new_n882), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n894), .B1(new_n892), .B2(new_n882), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n890), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n796), .ZN(new_n898));
  INV_X1    g712(.A(new_n375), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n374), .A2(new_n323), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n322), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n898), .A2(new_n797), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n903), .A2(new_n769), .A3(new_n882), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT51), .ZN(new_n905));
  OAI21_X1  g719(.A(new_n887), .B1(new_n897), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n897), .A2(KEYINPUT115), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT115), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n908), .B(new_n890), .C1(new_n895), .C2(new_n896), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(new_n909), .A3(new_n904), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT51), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n906), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT112), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT111), .B1(new_n856), .B2(KEYINPUT53), .ZN(new_n914));
  NOR4_X1   g728(.A1(new_n847), .A2(new_n855), .A3(new_n838), .A4(new_n867), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n847), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n864), .B1(new_n917), .B2(new_n859), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT53), .B1(new_n918), .B2(new_n861), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n913), .B(KEYINPUT54), .C1(new_n916), .C2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n856), .A2(KEYINPUT53), .A3(new_n863), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n867), .B1(new_n847), .B2(new_n855), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n923), .A2(KEYINPUT54), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n870), .A2(new_n912), .A3(new_n920), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n884), .A2(new_n250), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n901), .B(KEYINPUT49), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n929), .A2(new_n187), .A3(new_n321), .A4(new_n761), .ZN(new_n930));
  OR4_X1    g744(.A1(new_n872), .A2(new_n930), .A3(new_n698), .A4(new_n700), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n928), .A2(new_n931), .ZN(G75));
  NAND2_X1  g746(.A1(new_n474), .A2(new_n884), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT119), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n369), .B1(new_n921), .B2(new_n922), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n314), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT56), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n936), .A2(KEYINPUT118), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n249), .A2(new_n291), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT117), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n289), .B(KEYINPUT55), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n934), .B1(new_n938), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n938), .B2(new_n942), .ZN(G51));
  INV_X1    g758(.A(new_n934), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n372), .A2(new_n373), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n923), .B(new_n869), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n324), .B(KEYINPUT57), .Z(new_n948));
  OAI21_X1  g762(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n935), .A2(new_n779), .A3(new_n780), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n945), .B1(new_n949), .B2(new_n950), .ZN(G54));
  AND3_X1   g765(.A1(new_n935), .A2(KEYINPUT58), .A3(G475), .ZN(new_n952));
  INV_X1    g766(.A(new_n428), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n952), .A2(new_n953), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n945), .B1(new_n954), .B2(new_n955), .ZN(G60));
  AND2_X1   g770(.A1(new_n611), .A2(new_n613), .ZN(new_n957));
  NAND2_X1  g771(.A1(G478), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT59), .Z(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n957), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n934), .B1(new_n947), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n870), .A2(new_n920), .A3(new_n925), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n960), .ZN(new_n964));
  INV_X1    g778(.A(new_n957), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(G63));
  OAI21_X1  g780(.A(new_n934), .B1(KEYINPUT121), .B2(KEYINPUT61), .ZN(new_n967));
  XNOR2_X1  g781(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n441), .A2(new_n308), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n923), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n967), .B1(new_n971), .B2(new_n647), .ZN(new_n972));
  NAND2_X1  g786(.A1(KEYINPUT121), .A2(KEYINPUT61), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n923), .A2(new_n970), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n974), .A2(new_n585), .A3(new_n586), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n972), .A2(new_n973), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n973), .B1(new_n972), .B2(new_n975), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(G66));
  INV_X1    g792(.A(new_n477), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n250), .B1(new_n979), .B2(G224), .ZN(new_n980));
  INV_X1    g794(.A(new_n830), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n980), .B1(new_n981), .B2(new_n353), .ZN(new_n982));
  INV_X1    g796(.A(G898), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n940), .B1(new_n983), .B2(new_n474), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n982), .B(new_n984), .ZN(G69));
  AOI21_X1  g799(.A(new_n353), .B1(G227), .B2(G900), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT125), .Z(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n813), .A2(new_n815), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n678), .B1(new_n989), .B2(new_n617), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n841), .A2(new_n754), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n799), .A2(new_n791), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n744), .A2(new_n674), .A3(new_n708), .ZN(new_n993));
  OAI21_X1  g807(.A(KEYINPUT62), .B1(new_n704), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(KEYINPUT123), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT123), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n996), .B(KEYINPUT62), .C1(new_n704), .C2(new_n993), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n992), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n993), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT62), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n999), .A2(new_n1000), .A3(new_n701), .A4(new_n703), .ZN(new_n1001));
  INV_X1    g815(.A(KEYINPUT122), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n998), .A2(KEYINPUT124), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(KEYINPUT124), .B1(new_n998), .B2(new_n1003), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n353), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n498), .B1(new_n502), .B2(new_n503), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(new_n421), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  AND3_X1   g823(.A1(new_n799), .A2(new_n757), .A3(new_n759), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n786), .A2(new_n653), .A3(new_n873), .A4(new_n802), .ZN(new_n1011));
  OR2_X1    g825(.A1(new_n1011), .A2(KEYINPUT126), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n993), .B1(new_n1011), .B2(KEYINPUT126), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1010), .A2(new_n791), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(new_n353), .ZN(new_n1015));
  NOR2_X1   g829(.A1(new_n353), .A2(G900), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1008), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n988), .B1(new_n1009), .B2(new_n1019), .ZN(new_n1020));
  AOI211_X1 g834(.A(new_n987), .B(new_n1018), .C1(new_n1006), .C2(new_n1008), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1020), .A2(new_n1021), .ZN(G72));
  NAND2_X1  g836(.A1(G472), .A2(G902), .ZN(new_n1023));
  XOR2_X1   g837(.A(new_n1023), .B(KEYINPUT63), .Z(new_n1024));
  OAI21_X1  g838(.A(new_n1024), .B1(new_n1014), .B2(new_n981), .ZN(new_n1025));
  INV_X1    g839(.A(new_n537), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1026), .A2(new_n509), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n945), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1027), .ZN(new_n1029));
  INV_X1    g843(.A(new_n692), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n1029), .A2(new_n1030), .A3(new_n1024), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1031), .B(KEYINPUT127), .Z(new_n1032));
  OAI21_X1  g846(.A(new_n1028), .B1(new_n868), .B2(new_n1032), .ZN(new_n1033));
  OR2_X1    g847(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n1024), .B1(new_n1034), .B2(new_n981), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1033), .B1(new_n1035), .B2(new_n692), .ZN(G57));
endmodule


