//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1299, new_n1300, new_n1301, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383,
    new_n1384, new_n1385, new_n1386, new_n1387, new_n1388, new_n1389;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT64), .B(G20), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(new_n201), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G226), .ZN(new_n222));
  INV_X1    g0022(.A(G116), .ZN(new_n223));
  INV_X1    g0023(.A(G270), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n221), .B1(new_n202), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT65), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n227), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n225), .A2(new_n226), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n211), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n214), .B1(new_n218), .B2(new_n220), .C1(new_n232), .C2(KEYINPUT1), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT66), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT67), .ZN(new_n241));
  XOR2_X1   g0041(.A(G264), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n239), .B(new_n243), .Z(G358));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n245), .B(new_n246), .Z(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  AOI22_X1  g0052(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n215), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT72), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n253), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n216), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G13), .ZN(new_n262));
  NOR3_X1   g0062(.A1(new_n262), .A2(new_n209), .A3(G1), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(new_n260), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n202), .B1(new_n208), .B2(G20), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n264), .A2(new_n265), .B1(new_n202), .B2(new_n263), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n267), .B(KEYINPUT9), .ZN(new_n268));
  OR2_X1    g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT70), .ZN(new_n270));
  NAND2_X1  g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(KEYINPUT3), .A2(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  OAI21_X1  g0074(.A(KEYINPUT70), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n276), .A2(G222), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G77), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n276), .A2(G1698), .ZN(new_n280));
  INV_X1    g0080(.A(G223), .ZN(new_n281));
  OAI221_X1 g0081(.A(new_n278), .B1(new_n279), .B2(new_n276), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G1), .A3(G13), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n284), .A2(G274), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G45), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT68), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT68), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G45), .ZN(new_n292));
  INV_X1    g0092(.A(G41), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n290), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n208), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT69), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT69), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n294), .A2(new_n297), .A3(new_n208), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n288), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n284), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n299), .B1(G226), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n286), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT71), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n286), .A2(KEYINPUT71), .A3(new_n303), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n306), .A2(G200), .A3(new_n307), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n306), .A2(new_n307), .ZN(new_n309));
  INV_X1    g0109(.A(G190), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n268), .B(new_n308), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT10), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT76), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n312), .B1(new_n308), .B2(new_n313), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n311), .B(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n306), .A2(new_n307), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n267), .B1(new_n316), .B2(G169), .ZN(new_n317));
  INV_X1    g0117(.A(G179), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n317), .A2(KEYINPUT73), .B1(new_n318), .B2(new_n316), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(KEYINPUT73), .B2(new_n317), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G68), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n252), .A2(G50), .B1(G20), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n256), .B2(new_n279), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n324), .A2(KEYINPUT11), .A3(new_n260), .ZN(new_n325));
  AOI21_X1  g0125(.A(KEYINPUT11), .B1(new_n324), .B2(new_n260), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT79), .B1(new_n263), .B2(new_n322), .ZN(new_n327));
  XNOR2_X1  g0127(.A(new_n327), .B(KEYINPUT12), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n208), .A2(G20), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n264), .A2(G68), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NOR3_X1   g0131(.A1(new_n325), .A2(new_n326), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT14), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT78), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT77), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n301), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n284), .A2(KEYINPUT77), .A3(new_n300), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n337), .A2(G238), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n335), .B1(new_n299), .B2(new_n340), .ZN(new_n341));
  AND3_X1   g0141(.A1(new_n294), .A2(new_n297), .A3(new_n208), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n297), .B1(new_n294), .B2(new_n208), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n287), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(KEYINPUT78), .A3(new_n339), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT13), .ZN(new_n347));
  NAND2_X1  g0147(.A1(G33), .A2(G97), .ZN(new_n348));
  INV_X1    g0148(.A(G232), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n348), .B1(new_n280), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n276), .A2(new_n277), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(new_n222), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n285), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n346), .A2(new_n347), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n347), .B1(new_n346), .B2(new_n353), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n334), .B(G169), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n346), .A2(new_n353), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT13), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n359), .A2(G179), .A3(new_n354), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n354), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n334), .B1(new_n362), .B2(G169), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n333), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(G200), .B1(new_n355), .B2(new_n356), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n359), .A2(G190), .A3(new_n354), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n365), .A2(new_n366), .A3(new_n332), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n364), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n264), .ZN(new_n370));
  INV_X1    g0170(.A(new_n257), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n329), .ZN(new_n372));
  INV_X1    g0172(.A(new_n263), .ZN(new_n373));
  OAI22_X1  g0173(.A1(new_n370), .A2(new_n372), .B1(new_n373), .B2(new_n371), .ZN(new_n374));
  INV_X1    g0174(.A(new_n260), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n252), .A2(G159), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT82), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G58), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(new_n322), .ZN(new_n380));
  OAI21_X1  g0180(.A(G20), .B1(new_n380), .B2(new_n201), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  AND2_X1   g0182(.A1(KEYINPUT80), .A2(G33), .ZN(new_n383));
  NOR2_X1   g0183(.A1(KEYINPUT80), .A2(G33), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT3), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(new_n215), .A3(new_n269), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT7), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g0188(.A(KEYINPUT80), .B(G33), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n274), .B1(new_n389), .B2(KEYINPUT3), .ZN(new_n390));
  OR2_X1    g0190(.A1(KEYINPUT81), .A2(KEYINPUT7), .ZN(new_n391));
  NAND2_X1  g0191(.A1(KEYINPUT81), .A2(KEYINPUT7), .ZN(new_n392));
  AOI21_X1  g0192(.A(G20), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n388), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n382), .B1(new_n395), .B2(G68), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n375), .B1(new_n396), .B2(KEYINPUT16), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT16), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n209), .A2(KEYINPUT64), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT64), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G20), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n402), .A2(new_n387), .A3(new_n273), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(KEYINPUT3), .B2(new_n389), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n391), .A2(new_n392), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n276), .B2(G20), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n322), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n398), .B1(new_n407), .B2(new_n382), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n374), .B1(new_n397), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n281), .A2(new_n277), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n222), .A2(G1698), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n385), .B2(new_n269), .ZN(new_n413));
  INV_X1    g0213(.A(G33), .ZN(new_n414));
  INV_X1    g0214(.A(G87), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n285), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n301), .A2(new_n349), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n344), .A2(new_n417), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(G200), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n344), .A2(new_n310), .A3(new_n417), .A4(new_n419), .ZN(new_n423));
  AND3_X1   g0223(.A1(new_n422), .A2(KEYINPUT83), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT83), .B1(new_n422), .B2(new_n423), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n409), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT17), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n296), .A2(new_n298), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n418), .B1(new_n429), .B2(new_n287), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n430), .A2(G179), .A3(new_n417), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n420), .A2(G169), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(KEYINPUT18), .B1(new_n409), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n397), .A2(new_n408), .ZN(new_n436));
  INV_X1    g0236(.A(new_n374), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n438), .A2(new_n439), .A3(new_n433), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n409), .B(KEYINPUT17), .C1(new_n425), .C2(new_n424), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n428), .A2(new_n435), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT74), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n351), .B2(new_n349), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n276), .A2(KEYINPUT74), .A3(G232), .A4(new_n277), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G238), .ZN(new_n448));
  INV_X1    g0248(.A(G107), .ZN(new_n449));
  OAI22_X1  g0249(.A1(new_n280), .A2(new_n448), .B1(new_n449), .B2(new_n276), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n284), .B1(new_n447), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(G244), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n344), .B1(new_n453), .B2(new_n301), .ZN(new_n454));
  OAI21_X1  g0254(.A(KEYINPUT75), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT75), .ZN(new_n456));
  INV_X1    g0256(.A(new_n454), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n450), .B1(new_n445), .B2(new_n446), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n456), .B(new_n457), .C1(new_n458), .C2(new_n284), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n318), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n371), .A2(new_n252), .B1(G77), .B2(new_n402), .ZN(new_n462));
  XNOR2_X1  g0262(.A(KEYINPUT15), .B(G87), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n464), .A2(G33), .A3(new_n215), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n375), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n264), .A2(G77), .A3(new_n329), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(G77), .B2(new_n373), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(G169), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n455), .A2(new_n471), .A3(new_n459), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n461), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n310), .B1(new_n455), .B2(new_n459), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n455), .A2(G200), .A3(new_n459), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(new_n469), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n443), .B(new_n473), .C1(new_n474), .C2(new_n476), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n321), .A2(new_n369), .A3(new_n477), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n478), .A2(KEYINPUT84), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT84), .ZN(new_n480));
  NOR4_X1   g0280(.A1(new_n321), .A2(new_n477), .A3(new_n480), .A4(new_n369), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n289), .A2(G1), .ZN(new_n483));
  XNOR2_X1  g0283(.A(KEYINPUT5), .B(G41), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n287), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  AND2_X1   g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  NOR2_X1   g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n483), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n284), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n485), .B1(new_n224), .B2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT88), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n277), .A2(G257), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n491), .B1(new_n390), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n385), .A2(new_n269), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n494), .A2(KEYINPUT88), .A3(G257), .A4(new_n277), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n272), .A2(new_n275), .A3(G303), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(G264), .A3(G1698), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n493), .A2(new_n495), .A3(new_n496), .A4(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n490), .B1(new_n498), .B2(new_n285), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G190), .ZN(new_n500));
  INV_X1    g0300(.A(G283), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n215), .B1(new_n414), .B2(new_n501), .ZN(new_n502));
  OR2_X1    g0302(.A1(KEYINPUT85), .A2(G97), .ZN(new_n503));
  NAND2_X1  g0303(.A1(KEYINPUT85), .A2(G97), .ZN(new_n504));
  AOI21_X1  g0304(.A(G33), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OR2_X1    g0305(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT20), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n259), .A2(new_n216), .B1(G20), .B2(new_n223), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n506), .A2(KEYINPUT89), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n373), .A2(G116), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n208), .A2(G33), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n264), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n510), .B1(new_n513), .B2(G116), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n508), .B1(new_n502), .B2(new_n505), .ZN(new_n515));
  OR2_X1    g0315(.A1(new_n507), .A2(KEYINPUT89), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n507), .A2(KEYINPUT89), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n509), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n500), .B(new_n520), .C1(new_n421), .C2(new_n499), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT21), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n519), .A2(G169), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n522), .B1(new_n523), .B2(new_n499), .ZN(new_n524));
  AOI211_X1 g0324(.A(new_n318), .B(new_n490), .C1(new_n498), .C2(new_n285), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n519), .ZN(new_n526));
  INV_X1    g0326(.A(new_n499), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n527), .A2(KEYINPUT21), .A3(G169), .A4(new_n519), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n521), .A2(new_n524), .A3(new_n526), .A4(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT24), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT22), .B1(new_n276), .B2(G87), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT23), .B1(new_n209), .B2(G107), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT90), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(KEYINPUT90), .B(KEYINPUT23), .C1(new_n209), .C2(G107), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n389), .A2(new_n209), .A3(G116), .ZN(new_n537));
  OAI21_X1  g0337(.A(KEYINPUT22), .B1(KEYINPUT23), .B2(G107), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n402), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n531), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(KEYINPUT22), .A2(G87), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n390), .A2(new_n402), .A3(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n530), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  OR2_X1    g0345(.A1(KEYINPUT80), .A2(G33), .ZN(new_n546));
  NAND2_X1  g0346(.A1(KEYINPUT80), .A2(G33), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n223), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n548), .A2(new_n209), .B1(new_n402), .B2(new_n538), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n415), .B1(new_n272), .B2(new_n275), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n549), .B(new_n536), .C1(new_n550), .C2(KEYINPUT22), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n551), .A2(KEYINPUT24), .A3(new_n543), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n260), .B1(new_n545), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(KEYINPUT25), .B1(new_n263), .B2(new_n449), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n263), .A2(KEYINPUT25), .A3(new_n449), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n513), .A2(G107), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(G250), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n277), .ZN(new_n560));
  INV_X1    g0360(.A(G257), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G1698), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n385), .B2(new_n269), .ZN(new_n564));
  INV_X1    g0364(.A(G294), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n546), .B2(new_n547), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n285), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n216), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n484), .A2(new_n483), .B1(new_n568), .B2(new_n283), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT91), .B1(new_n569), .B2(G264), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n488), .A2(G264), .A3(new_n284), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT91), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n567), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT92), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n569), .A2(KEYINPUT91), .A3(G264), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n571), .A2(new_n572), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n579), .A2(KEYINPUT92), .A3(new_n567), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n576), .A2(G179), .A3(new_n485), .A4(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n485), .ZN(new_n582));
  OAI21_X1  g0382(.A(G169), .B1(new_n574), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n558), .A2(new_n584), .ZN(new_n585));
  NOR3_X1   g0385(.A1(new_n574), .A2(G190), .A3(new_n582), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n576), .A2(new_n485), .A3(new_n580), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n586), .B1(new_n587), .B2(new_n421), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n585), .B1(new_n558), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n485), .B1(new_n561), .B2(new_n489), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n277), .A2(KEYINPUT4), .A3(G244), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n559), .B2(new_n277), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n276), .A2(new_n592), .B1(G33), .B2(G283), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT4), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n277), .A2(G244), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n594), .B1(new_n390), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n590), .B1(new_n597), .B2(new_n285), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n318), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n284), .B1(new_n593), .B2(new_n596), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n471), .B1(new_n600), .B2(new_n590), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n404), .A2(new_n406), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(G107), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n503), .A2(new_n504), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n604), .A2(KEYINPUT6), .A3(new_n449), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT6), .ZN(new_n606));
  INV_X1    g0406(.A(G97), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(new_n449), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n606), .B1(new_n608), .B2(new_n205), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n610), .A2(new_n402), .B1(G77), .B2(new_n252), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n375), .B1(new_n603), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n512), .A2(G97), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT86), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n373), .A2(new_n607), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n614), .B1(new_n613), .B2(new_n615), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n599), .B(new_n601), .C1(new_n612), .C2(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n503), .A2(new_n415), .A3(new_n449), .A4(new_n504), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT19), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n215), .B1(new_n621), .B2(new_n348), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n604), .A2(G33), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n620), .A2(new_n622), .B1(new_n623), .B2(new_n621), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n494), .A2(G68), .A3(new_n215), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n375), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n512), .A2(new_n463), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n464), .A2(new_n373), .ZN(new_n628));
  OR3_X1    g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n453), .A2(G1698), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(G238), .B2(G1698), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n269), .B2(new_n385), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n285), .B1(new_n632), .B2(new_n548), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n483), .A2(new_n559), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n287), .A2(new_n483), .B1(new_n284), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n471), .ZN(new_n637));
  INV_X1    g0437(.A(new_n636), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n318), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n629), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n598), .A2(G190), .ZN(new_n641));
  INV_X1    g0441(.A(new_n611), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n449), .B1(new_n404), .B2(new_n406), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n260), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n613), .A2(new_n615), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT86), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(G200), .B1(new_n600), .B2(new_n590), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n641), .A2(new_n644), .A3(new_n648), .A4(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n512), .A2(new_n415), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n626), .A2(new_n628), .A3(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT87), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n636), .B2(new_n310), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n636), .A2(G200), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n633), .A2(KEYINPUT87), .A3(G190), .A4(new_n635), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n652), .A2(new_n654), .A3(new_n655), .A4(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n619), .A2(new_n640), .A3(new_n650), .A4(new_n657), .ZN(new_n658));
  NOR4_X1   g0458(.A1(new_n482), .A2(new_n529), .A3(new_n589), .A4(new_n658), .ZN(G372));
  INV_X1    g0459(.A(KEYINPUT83), .ZN(new_n660));
  AOI21_X1  g0460(.A(G200), .B1(new_n430), .B2(new_n417), .ZN(new_n661));
  INV_X1    g0461(.A(new_n423), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n422), .A2(KEYINPUT83), .A3(new_n423), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(KEYINPUT17), .B1(new_n665), .B2(new_n409), .ZN(new_n666));
  INV_X1    g0466(.A(new_n441), .ZN(new_n667));
  OR2_X1    g0467(.A1(new_n367), .A2(new_n473), .ZN(new_n668));
  AOI211_X1 g0468(.A(new_n666), .B(new_n667), .C1(new_n668), .C2(new_n364), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n440), .A2(new_n435), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n315), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n671), .A2(new_n320), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n619), .A2(new_n650), .ZN(new_n673));
  AOI21_X1  g0473(.A(KEYINPUT93), .B1(new_n636), .B2(new_n471), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n636), .A2(KEYINPUT93), .A3(new_n471), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n629), .B(new_n639), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n652), .B(new_n655), .C1(new_n310), .C2(new_n636), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT94), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT94), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n676), .A2(new_n680), .A3(new_n677), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n673), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n588), .A2(new_n558), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n524), .A2(new_n528), .A3(new_n526), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n683), .B1(new_n685), .B2(new_n585), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n676), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n640), .A2(new_n657), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(new_n619), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(KEYINPUT26), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n619), .ZN(new_n693));
  INV_X1    g0493(.A(new_n681), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n680), .B1(new_n676), .B2(new_n677), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n693), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT26), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n692), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n688), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n672), .B1(new_n482), .B2(new_n699), .ZN(G369));
  NAND3_X1  g0500(.A1(new_n215), .A2(new_n208), .A3(G13), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(KEYINPUT27), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G213), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(G343), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n520), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n684), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n529), .B2(new_n708), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G330), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n589), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n558), .A2(new_n706), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n585), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n706), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n712), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n685), .A2(new_n706), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n720), .A2(new_n713), .B1(new_n716), .B2(new_n707), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n719), .A2(new_n721), .ZN(G399));
  INV_X1    g0522(.A(new_n212), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G41), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n620), .A2(G116), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(G1), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n220), .B2(new_n725), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT28), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n707), .B1(new_n688), .B2(new_n698), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT29), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n676), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n733), .B1(new_n690), .B2(new_n697), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT96), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n673), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n619), .A2(KEYINPUT96), .A3(new_n650), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n736), .B(new_n737), .C1(new_n694), .C2(new_n695), .ZN(new_n738));
  OAI22_X1  g0538(.A1(new_n716), .A2(new_n684), .B1(new_n558), .B2(new_n588), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n734), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n696), .A2(KEYINPUT26), .ZN(new_n741));
  OAI211_X1 g0541(.A(KEYINPUT29), .B(new_n707), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n732), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n706), .A2(KEYINPUT31), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n576), .A2(new_n598), .A3(new_n580), .A4(new_n638), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n499), .A2(G179), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n598), .A2(new_n638), .A3(G179), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(new_n527), .A3(new_n587), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(KEYINPUT95), .ZN(new_n752));
  AND3_X1   g0552(.A1(new_n579), .A2(KEYINPUT92), .A3(new_n567), .ZN(new_n753));
  AOI21_X1  g0553(.A(KEYINPUT92), .B1(new_n579), .B2(new_n567), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n600), .A2(new_n636), .A3(new_n590), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n755), .A2(new_n525), .A3(KEYINPUT30), .A4(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n752), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n751), .A2(KEYINPUT95), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n744), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n529), .ZN(new_n762));
  INV_X1    g0562(.A(new_n658), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n713), .A2(new_n762), .A3(new_n763), .A4(new_n707), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n748), .A2(new_n750), .A3(new_n757), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(new_n706), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT31), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(G330), .B1(new_n761), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n743), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n729), .B1(new_n772), .B2(G1), .ZN(G364));
  NOR2_X1   g0573(.A1(new_n402), .A2(new_n262), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G45), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT97), .Z(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n777), .A2(new_n208), .A3(new_n724), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n712), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(G330), .B2(new_n710), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G13), .A2(G33), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n216), .B1(G20), .B2(new_n471), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n723), .A2(new_n494), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n290), .A2(new_n292), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(new_n220), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n247), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n788), .B1(G45), .B2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n276), .A2(new_n212), .ZN(new_n791));
  INV_X1    g0591(.A(G355), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n791), .A2(new_n792), .B1(G116), .B2(new_n212), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n785), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n778), .ZN(new_n795));
  INV_X1    g0595(.A(new_n276), .ZN(new_n796));
  INV_X1    g0596(.A(G303), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n421), .A2(G179), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n798), .A2(G20), .A3(G190), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G179), .A2(G200), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G190), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n402), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n796), .B1(new_n797), .B2(new_n799), .C1(new_n803), .C2(new_n565), .ZN(new_n804));
  NOR4_X1   g0604(.A1(new_n215), .A2(new_n318), .A3(G190), .A4(G200), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G311), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n402), .A2(new_n310), .A3(new_n798), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n806), .A2(new_n807), .B1(new_n501), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n318), .A2(new_n421), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n402), .A2(G190), .A3(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI211_X1 g0612(.A(new_n804), .B(new_n809), .C1(G326), .C2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n402), .A2(new_n310), .A3(new_n810), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(KEYINPUT33), .B(G317), .ZN(new_n816));
  NOR3_X1   g0616(.A1(new_n318), .A2(new_n310), .A3(G200), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n402), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n815), .A2(new_n816), .B1(new_n819), .B2(G322), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT101), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n402), .A2(new_n310), .A3(new_n800), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT100), .Z(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(G329), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n813), .A2(new_n821), .A3(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n276), .B1(new_n415), .B2(new_n799), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n202), .A2(new_n811), .B1(new_n808), .B2(new_n449), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n826), .B(new_n827), .C1(G58), .C2(new_n819), .ZN(new_n828));
  INV_X1    g0628(.A(G159), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n822), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT32), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n806), .A2(KEYINPUT98), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n806), .A2(KEYINPUT98), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n828), .B(new_n831), .C1(new_n279), .C2(new_n834), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n803), .A2(new_n607), .B1(new_n814), .B2(new_n322), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT99), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n825), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n795), .B1(new_n838), .B2(new_n784), .ZN(new_n839));
  INV_X1    g0639(.A(new_n783), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n839), .B1(new_n710), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n780), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G396));
  NAND2_X1  g0643(.A1(new_n696), .A2(new_n697), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n691), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n733), .B1(new_n682), .B2(new_n686), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n706), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n470), .A2(new_n706), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n476), .B2(new_n474), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n473), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n461), .A2(new_n470), .A3(new_n472), .A4(new_n707), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n847), .B(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n778), .B1(new_n854), .B2(new_n770), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n770), .B2(new_n854), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n784), .A2(new_n781), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT102), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n778), .B1(G77), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n834), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n860), .A2(G116), .B1(G311), .B2(new_n823), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n803), .A2(new_n607), .B1(new_n818), .B2(new_n565), .ZN(new_n862));
  INV_X1    g0662(.A(new_n799), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n276), .B(new_n862), .C1(G107), .C2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n808), .A2(new_n415), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n811), .A2(new_n797), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n865), .B(new_n866), .C1(G283), .C2(new_n815), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n861), .A2(new_n864), .A3(new_n867), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n812), .A2(G137), .B1(new_n819), .B2(G143), .ZN(new_n869));
  INV_X1    g0669(.A(G150), .ZN(new_n870));
  OAI221_X1 g0670(.A(new_n869), .B1(new_n870), .B2(new_n814), .C1(new_n834), .C2(new_n829), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n871), .B(KEYINPUT34), .Z(new_n872));
  NOR2_X1   g0672(.A1(new_n808), .A2(new_n322), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n494), .B1(new_n202), .B2(new_n799), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n873), .B(new_n874), .C1(G58), .C2(new_n802), .ZN(new_n875));
  INV_X1    g0675(.A(G132), .ZN(new_n876));
  INV_X1    g0676(.A(new_n823), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n868), .B1(new_n872), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n859), .B1(new_n879), .B2(new_n784), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n853), .B2(new_n782), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n856), .A2(new_n881), .ZN(G384));
  AOI211_X1 g0682(.A(new_n223), .B(new_n218), .C1(new_n610), .C2(KEYINPUT35), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(KEYINPUT35), .B2(new_n610), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n884), .B(KEYINPUT36), .Z(new_n885));
  OR3_X1    g0685(.A1(new_n220), .A2(new_n279), .A3(new_n380), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n202), .A2(G68), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n208), .B(G13), .C1(new_n886), .C2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n851), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(new_n847), .B2(new_n853), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n333), .A2(new_n706), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n364), .A2(new_n368), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(G169), .B1(new_n355), .B2(new_n356), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT14), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n895), .A2(new_n360), .A3(new_n357), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n333), .B(new_n706), .C1(new_n896), .C2(new_n367), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n893), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT103), .B1(new_n891), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n851), .B1(new_n730), .B2(new_n852), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT103), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n893), .A2(new_n897), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT38), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n395), .A2(G68), .ZN(new_n905));
  INV_X1    g0705(.A(new_n382), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(KEYINPUT16), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n260), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n396), .A2(KEYINPUT16), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n437), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n704), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n667), .A2(new_n666), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n440), .A2(new_n435), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT37), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n431), .A2(new_n432), .A3(new_n704), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n910), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n916), .B1(new_n426), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n438), .A2(new_n917), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n920), .A2(new_n426), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n919), .B1(new_n921), .B2(new_n916), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n904), .B1(new_n915), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n920), .A2(new_n426), .A3(new_n916), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n426), .A2(new_n918), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n924), .B1(new_n925), .B2(new_n916), .ZN(new_n926));
  OAI211_X1 g0726(.A(KEYINPUT38), .B(new_n926), .C1(new_n443), .C2(new_n912), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n923), .A2(KEYINPUT104), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT104), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n929), .B(new_n904), .C1(new_n915), .C2(new_n922), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n899), .A2(new_n903), .A3(new_n932), .ZN(new_n933));
  AND3_X1   g0733(.A1(new_n442), .A2(new_n438), .A3(new_n911), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n916), .B1(new_n920), .B2(new_n426), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(KEYINPUT105), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT105), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n924), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n936), .B1(new_n938), .B2(new_n935), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n904), .B1(new_n934), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT39), .B1(new_n940), .B2(new_n927), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n941), .B1(new_n931), .B2(KEYINPUT39), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n896), .A2(new_n333), .A3(new_n707), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n670), .A2(new_n704), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n933), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  OAI211_X1 g0747(.A(new_n732), .B(new_n742), .C1(new_n479), .C2(new_n481), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n672), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n947), .B(new_n949), .Z(new_n950));
  INV_X1    g0750(.A(G330), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT106), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n765), .A2(KEYINPUT31), .A3(new_n706), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n764), .A2(new_n952), .A3(new_n768), .A4(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n768), .A2(new_n953), .ZN(new_n955));
  NOR4_X1   g0755(.A1(new_n589), .A2(new_n529), .A3(new_n658), .A4(new_n706), .ZN(new_n956));
  OAI21_X1  g0756(.A(KEYINPUT106), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n482), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n954), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n852), .B1(new_n893), .B2(new_n897), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n928), .A2(new_n930), .A3(new_n959), .A4(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT40), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n959), .A2(new_n960), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n962), .B1(new_n940), .B2(new_n927), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n961), .A2(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n951), .B1(new_n958), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n965), .B2(new_n958), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n950), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n208), .B2(new_n774), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n950), .A2(new_n967), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n889), .B1(new_n969), .B2(new_n970), .ZN(G367));
  OAI21_X1  g0771(.A(new_n706), .B1(new_n612), .B2(new_n618), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n736), .A2(new_n737), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n693), .A2(new_n706), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(KEYINPUT107), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT107), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n981), .A2(new_n719), .ZN(new_n982));
  INV_X1    g0782(.A(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n980), .A2(new_n716), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n706), .B1(new_n984), .B2(new_n619), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n720), .A2(new_n713), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n976), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT42), .Z(new_n988));
  NOR2_X1   g0788(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT108), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(KEYINPUT108), .B1(new_n985), .B2(new_n988), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n652), .A2(new_n707), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n679), .B2(new_n681), .ZN(new_n994));
  NOR3_X1   g0794(.A1(new_n676), .A2(new_n652), .A3(new_n707), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT43), .Z(new_n997));
  NAND3_X1  g0797(.A1(new_n991), .A2(new_n992), .A3(new_n997), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n991), .A2(new_n992), .ZN(new_n999));
  INV_X1    g0799(.A(new_n996), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n1000), .A2(KEYINPUT43), .ZN(new_n1001));
  OAI211_X1 g0801(.A(new_n983), .B(new_n998), .C1(new_n999), .C2(new_n1001), .ZN(new_n1002));
  AND3_X1   g0802(.A1(new_n991), .A2(new_n992), .A3(new_n997), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1001), .B1(new_n991), .B2(new_n992), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n982), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n777), .A2(new_n208), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n721), .A2(new_n975), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT45), .Z(new_n1008));
  NOR2_X1   g0808(.A1(new_n721), .A2(new_n975), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT44), .ZN(new_n1010));
  AND3_X1   g0810(.A1(new_n1008), .A2(new_n719), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n719), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n986), .B1(new_n718), .B2(new_n720), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(new_n712), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n771), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n724), .B(KEYINPUT41), .Z(new_n1017));
  OAI21_X1  g0817(.A(new_n1006), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1002), .A2(new_n1005), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n786), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n243), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n785), .B1(new_n212), .B2(new_n463), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n778), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n822), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(G311), .A2(new_n812), .B1(new_n1024), .B2(G317), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n604), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1025), .B1(new_n1026), .B2(new_n808), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n863), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT46), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n799), .B2(new_n223), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1028), .B(new_n1030), .C1(new_n449), .C2(new_n803), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n390), .B1(new_n818), .B2(new_n797), .C1(new_n565), .C2(new_n814), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n1027), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n501), .B2(new_n834), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n802), .A2(G68), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n870), .B2(new_n818), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n796), .B(new_n1036), .C1(G58), .C2(new_n863), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n808), .A2(new_n279), .ZN(new_n1038));
  INV_X1    g0838(.A(G143), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n1039), .A2(new_n811), .B1(new_n814), .B2(new_n829), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n1038), .B(new_n1040), .C1(G137), .C2(new_n1024), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1037), .B(new_n1041), .C1(new_n202), .C2(new_n834), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1034), .A2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT47), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1023), .B1(new_n1044), .B2(new_n784), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n1000), .B2(new_n840), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1019), .A2(new_n1046), .ZN(G387));
  INV_X1    g0847(.A(new_n1006), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n791), .A2(new_n726), .B1(G107), .B2(new_n212), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n726), .ZN(new_n1050));
  AOI211_X1 g0850(.A(G45), .B(new_n1050), .C1(G68), .C2(G77), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n257), .A2(G50), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT50), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1020), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1054), .A2(KEYINPUT109), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n239), .B2(new_n787), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(KEYINPUT109), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1049), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n785), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n778), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n802), .A2(new_n464), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n202), .B2(new_n818), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n390), .B(new_n1062), .C1(G77), .C2(new_n863), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n806), .A2(new_n322), .B1(new_n870), .B2(new_n822), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G159), .B2(new_n812), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n808), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(G97), .A2(new_n1066), .B1(new_n815), .B2(new_n371), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1063), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n494), .B1(new_n1024), .B2(G326), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n803), .A2(new_n501), .B1(new_n565), .B2(new_n799), .ZN(new_n1070));
  INV_X1    g0870(.A(G317), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n814), .A2(new_n807), .B1(new_n818), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G322), .B2(new_n812), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n834), .B2(new_n797), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT48), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1070), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n1075), .B2(new_n1074), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT49), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1069), .B1(new_n223), .B2(new_n808), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1068), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT110), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n784), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1060), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n715), .A2(new_n717), .A3(new_n783), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1015), .A2(new_n1048), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n772), .A2(new_n1015), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1089), .A2(new_n724), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n772), .A2(new_n1015), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1088), .B1(new_n1090), .B2(new_n1091), .ZN(G393));
  INV_X1    g0892(.A(new_n1089), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n725), .B1(new_n1093), .B2(new_n1013), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n1093), .B2(new_n1013), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n785), .B1(new_n212), .B2(new_n1026), .C1(new_n1020), .C2(new_n250), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n796), .B1(new_n501), .B2(new_n799), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G303), .A2(new_n815), .B1(new_n1024), .B2(G322), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n1098), .B1(new_n449), .B2(new_n808), .C1(new_n565), .C2(new_n806), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1097), .B(new_n1099), .C1(G116), .C2(new_n802), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n811), .A2(new_n1071), .B1(new_n818), .B2(new_n807), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT52), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n494), .B1(new_n322), .B2(new_n799), .C1(new_n803), .C2(new_n279), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n865), .B1(G50), .B2(new_n815), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n1039), .B2(new_n822), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1103), .B(new_n1105), .C1(new_n860), .C2(new_n371), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n811), .A2(new_n870), .B1(new_n818), .B2(new_n829), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT51), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1100), .A2(new_n1102), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n778), .B(new_n1096), .C1(new_n1109), .C2(new_n1084), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(new_n981), .B2(new_n783), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n1013), .B2(new_n1048), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1095), .A2(new_n1112), .ZN(G390));
  OAI211_X1 g0913(.A(new_n707), .B(new_n850), .C1(new_n740), .C2(new_n741), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n851), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n902), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n940), .A2(new_n927), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n943), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n770), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n960), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n944), .B1(new_n900), .B2(new_n902), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1118), .B(new_n1120), .C1(new_n1121), .C2(new_n942), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n898), .B1(new_n851), .B2(new_n1114), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1117), .A2(new_n943), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n931), .A2(KEYINPUT39), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n941), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n943), .B1(new_n891), .B2(new_n898), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1125), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT111), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n951), .B1(new_n957), .B2(new_n954), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n960), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1131), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1132), .A2(KEYINPUT111), .A3(new_n960), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1122), .B1(new_n1130), .B2(new_n1137), .ZN(new_n1138));
  OR2_X1    g0938(.A1(new_n1138), .A2(new_n1006), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n778), .B1(new_n371), .B2(new_n858), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n819), .A2(G116), .B1(new_n802), .B2(G77), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT113), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n834), .B2(new_n1026), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n276), .B(new_n873), .C1(G87), .C2(new_n863), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(G107), .A2(new_n815), .B1(new_n812), .B2(G283), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1144), .B(new_n1145), .C1(new_n877), .C2(new_n565), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT54), .B(G143), .ZN(new_n1147));
  INV_X1    g0947(.A(G125), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n834), .A2(new_n1147), .B1(new_n877), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n276), .B1(new_n818), .B2(new_n876), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(G159), .B2(new_n802), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n863), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT53), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n799), .B2(new_n870), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1152), .A2(new_n1154), .B1(new_n815), .B2(G137), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(G50), .A2(new_n1066), .B1(new_n812), .B2(G128), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1151), .A2(new_n1155), .A3(new_n1156), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n1143), .A2(new_n1146), .B1(new_n1149), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1140), .B1(new_n1158), .B2(new_n784), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n942), .B2(new_n782), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1139), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(KEYINPUT114), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1115), .B1(new_n1119), .B2(new_n960), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n898), .B1(new_n1133), .B2(new_n852), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT112), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n851), .B(new_n1114), .C1(new_n1134), .C2(new_n770), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n902), .B1(new_n1132), .B2(new_n853), .ZN(new_n1168));
  OAI21_X1  g0968(.A(KEYINPUT112), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1166), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n898), .B1(new_n770), .B2(new_n852), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1135), .A2(new_n1136), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n900), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1132), .B1(new_n479), .B2(new_n481), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n948), .A2(new_n672), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1174), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n725), .B1(new_n1178), .B2(new_n1138), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1179), .B1(new_n1138), .B2(new_n1178), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT114), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1139), .A2(new_n1181), .A3(new_n1160), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1162), .A2(new_n1180), .A3(new_n1182), .ZN(G378));
  INV_X1    g0983(.A(new_n947), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n951), .B1(new_n963), .B2(new_n964), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n961), .A2(new_n962), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT115), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1187), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1189));
  XNOR2_X1  g0989(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n267), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1192), .A2(new_n704), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n315), .A2(new_n320), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1194), .B1(new_n315), .B2(new_n320), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1191), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1197), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1199), .A2(new_n1195), .A3(new_n1190), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n1188), .A2(new_n1189), .A3(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1185), .A2(new_n1201), .A3(new_n1186), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1184), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n942), .A2(new_n944), .B1(new_n670), .B2(new_n704), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1206), .A2(new_n1203), .A3(new_n933), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(KEYINPUT115), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1201), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1208), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1006), .B1(new_n1205), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1211), .A2(new_n781), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n778), .B1(G50), .B2(new_n858), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n803), .A2(new_n870), .B1(new_n799), .B2(new_n1147), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G137), .A2(new_n805), .B1(new_n815), .B2(G132), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n1148), .B2(new_n811), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1218), .B(new_n1220), .C1(G128), .C2(new_n819), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1222), .A2(KEYINPUT59), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1222), .A2(KEYINPUT59), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n414), .B(new_n293), .C1(new_n808), .C2(new_n829), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G124), .B2(new_n1024), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1223), .A2(new_n1224), .A3(new_n1226), .ZN(new_n1227));
  OAI22_X1  g1027(.A1(new_n607), .A2(new_n814), .B1(new_n811), .B2(new_n223), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1035), .B1(new_n279), .B2(new_n799), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1228), .B(new_n1229), .C1(G107), .C2(new_n819), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n390), .A2(new_n293), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n808), .A2(new_n379), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n1231), .B(new_n1232), .C1(new_n464), .C2(new_n805), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n1230), .B(new_n1233), .C1(new_n501), .C2(new_n877), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT58), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1231), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1227), .A2(new_n1236), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1217), .B1(new_n1239), .B2(new_n784), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1216), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(KEYINPUT116), .B1(new_n1215), .B2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n947), .B1(new_n1213), .B2(new_n1203), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1189), .A2(new_n1201), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1207), .B1(new_n1212), .B2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1048), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT116), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n1248), .A3(new_n1241), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1243), .A2(new_n1249), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1166), .A2(new_n1169), .B1(new_n1172), .B2(new_n900), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1177), .B1(new_n1138), .B2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT57), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n725), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT117), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1202), .A2(new_n1256), .A3(new_n1207), .ZN(new_n1257));
  AOI21_X1  g1057(.A(KEYINPUT117), .B1(new_n1208), .B2(new_n1213), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1205), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1252), .A2(KEYINPUT57), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1255), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1250), .A2(new_n1262), .ZN(G375));
  OAI21_X1  g1063(.A(KEYINPUT118), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1017), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT118), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1251), .A2(new_n1266), .A3(new_n1176), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1264), .A2(new_n1265), .A3(new_n1178), .A4(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1174), .A2(KEYINPUT119), .A3(new_n1048), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n778), .B1(G68), .B2(new_n858), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1038), .B1(G294), .B2(new_n812), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1271), .B1(new_n223), .B2(new_n814), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n796), .B1(new_n607), .B2(new_n799), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1061), .B1(new_n501), .B2(new_n818), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1272), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  OAI221_X1 g1075(.A(new_n1275), .B1(new_n449), .B2(new_n834), .C1(new_n797), .C2(new_n877), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n494), .B1(new_n829), .B2(new_n799), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n803), .A2(new_n202), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n1277), .B(new_n1278), .C1(G137), .C2(new_n819), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n823), .A2(G128), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1232), .B1(G132), .B2(new_n812), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1147), .ZN(new_n1282));
  AOI22_X1  g1082(.A1(G150), .A2(new_n805), .B1(new_n815), .B2(new_n1282), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1279), .A2(new_n1280), .A3(new_n1281), .A4(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1276), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1270), .B1(new_n1285), .B2(new_n784), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1286), .B1(new_n902), .B2(new_n782), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT119), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1288), .B1(new_n1251), .B2(new_n1006), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1268), .A2(new_n1269), .A3(new_n1287), .A4(new_n1289), .ZN(new_n1290));
  XOR2_X1   g1090(.A(new_n1290), .B(KEYINPUT120), .Z(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(G381));
  INV_X1    g1092(.A(G378), .ZN(new_n1293));
  AND2_X1   g1093(.A1(new_n1019), .A2(new_n1046), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(G393), .A2(G396), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(G390), .A2(G384), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1293), .A2(new_n1294), .A3(new_n1295), .A4(new_n1296), .ZN(new_n1297));
  OR3_X1    g1097(.A1(G381), .A2(G375), .A3(new_n1297), .ZN(G407));
  NAND2_X1  g1098(.A1(new_n705), .A2(G213), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1299), .B(KEYINPUT121), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1293), .A2(new_n1300), .ZN(new_n1301));
  OAI211_X1 g1101(.A(G407), .B(G213), .C1(G375), .C2(new_n1301), .ZN(G409));
  INV_X1    g1102(.A(G390), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(G387), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(KEYINPUT125), .ZN(new_n1305));
  XNOR2_X1  g1105(.A(G393), .B(new_n842), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1294), .A2(G390), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n1305), .A2(new_n1306), .B1(new_n1307), .B2(new_n1304), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(G387), .A2(new_n1303), .ZN(new_n1309));
  AOI21_X1  g1109(.A(G390), .B1(new_n1019), .B2(new_n1046), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1306), .ZN(new_n1311));
  NOR4_X1   g1111(.A1(new_n1309), .A2(new_n1310), .A3(KEYINPUT125), .A4(new_n1311), .ZN(new_n1312));
  NOR2_X1   g1112(.A1(new_n1308), .A2(new_n1312), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1300), .ZN(new_n1315));
  AND3_X1   g1115(.A1(new_n1250), .A2(G378), .A3(new_n1262), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT122), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1259), .A2(new_n1317), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1256), .B1(new_n1202), .B2(new_n1207), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1208), .A2(new_n1213), .A3(KEYINPUT117), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1244), .B1(new_n1319), .B2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(KEYINPUT122), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1318), .A2(new_n1322), .A3(new_n1048), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n1252), .B(new_n1265), .C1(new_n1244), .C2(new_n1246), .ZN(new_n1324));
  AND2_X1   g1124(.A1(new_n1324), .A2(new_n1241), .ZN(new_n1325));
  AOI21_X1  g1125(.A(G378), .B1(new_n1323), .B2(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1315), .B1(new_n1316), .B2(new_n1326), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1300), .A2(G2897), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT124), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(G384), .A2(new_n1330), .ZN(new_n1331));
  XNOR2_X1  g1131(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1332), .B1(new_n1251), .B2(new_n1176), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1264), .A2(new_n1333), .A3(new_n1267), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1174), .A2(new_n1177), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n725), .B1(new_n1335), .B2(KEYINPUT60), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1334), .A2(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n856), .A2(KEYINPUT124), .A3(new_n881), .ZN(new_n1338));
  AND4_X1   g1138(.A1(new_n1269), .A2(new_n1289), .A3(new_n1338), .A4(new_n1287), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1331), .B1(new_n1337), .B2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1337), .A2(new_n1339), .A3(new_n1331), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1329), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1342), .ZN(new_n1344));
  NOR3_X1   g1144(.A1(new_n1344), .A2(new_n1340), .A3(new_n1328), .ZN(new_n1345));
  NOR2_X1   g1145(.A1(new_n1343), .A2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1327), .A2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT61), .ZN(new_n1348));
  AOI21_X1  g1148(.A(KEYINPUT126), .B1(new_n1347), .B2(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1350));
  OAI211_X1 g1150(.A(new_n1315), .B(new_n1350), .C1(new_n1316), .C2(new_n1326), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(KEYINPUT62), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1048), .B1(new_n1321), .B2(KEYINPUT122), .ZN(new_n1353));
  AOI211_X1 g1153(.A(new_n1317), .B(new_n1244), .C1(new_n1319), .C2(new_n1320), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1325), .B1(new_n1353), .B2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1355), .A2(new_n1293), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1250), .A2(new_n1262), .A3(G378), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1300), .B1(new_n1356), .B2(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT62), .ZN(new_n1359));
  NAND3_X1  g1159(.A1(new_n1358), .A2(new_n1359), .A3(new_n1350), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1352), .A2(new_n1360), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1314), .B1(new_n1349), .B2(new_n1361), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1356), .A2(new_n1357), .ZN(new_n1363));
  AND4_X1   g1163(.A1(KEYINPUT63), .A2(new_n1363), .A3(new_n1315), .A4(new_n1350), .ZN(new_n1364));
  AOI21_X1  g1164(.A(KEYINPUT63), .B1(new_n1358), .B2(new_n1350), .ZN(new_n1365));
  OAI21_X1  g1165(.A(new_n1313), .B1(new_n1364), .B2(new_n1365), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT126), .ZN(new_n1367));
  OAI21_X1  g1167(.A(new_n1367), .B1(new_n1308), .B2(new_n1312), .ZN(new_n1368));
  OR2_X1    g1168(.A1(new_n1343), .A2(new_n1345), .ZN(new_n1369));
  OAI211_X1 g1169(.A(new_n1368), .B(new_n1348), .C1(new_n1369), .C2(new_n1358), .ZN(new_n1370));
  INV_X1    g1170(.A(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1366), .A2(new_n1371), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1362), .A2(new_n1372), .ZN(G405));
  NAND2_X1  g1173(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1307), .A2(new_n1304), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1374), .A2(new_n1375), .ZN(new_n1376));
  NAND4_X1  g1176(.A1(new_n1305), .A2(new_n1304), .A3(new_n1307), .A4(new_n1306), .ZN(new_n1377));
  NAND4_X1  g1177(.A1(new_n1376), .A2(new_n1377), .A3(new_n1341), .A4(new_n1342), .ZN(new_n1378));
  OAI21_X1  g1178(.A(new_n1350), .B1(new_n1308), .B2(new_n1312), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1378), .A2(new_n1379), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1380), .A2(KEYINPUT127), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(G375), .A2(new_n1293), .ZN(new_n1382));
  INV_X1    g1182(.A(KEYINPUT127), .ZN(new_n1383));
  NAND3_X1  g1183(.A1(new_n1378), .A2(new_n1383), .A3(new_n1379), .ZN(new_n1384));
  NAND4_X1  g1184(.A1(new_n1381), .A2(new_n1357), .A3(new_n1382), .A4(new_n1384), .ZN(new_n1385));
  NAND2_X1  g1185(.A1(new_n1382), .A2(new_n1357), .ZN(new_n1386));
  AND3_X1   g1186(.A1(new_n1378), .A2(new_n1383), .A3(new_n1379), .ZN(new_n1387));
  AOI21_X1  g1187(.A(new_n1383), .B1(new_n1378), .B2(new_n1379), .ZN(new_n1388));
  OAI21_X1  g1188(.A(new_n1386), .B1(new_n1387), .B2(new_n1388), .ZN(new_n1389));
  NAND2_X1  g1189(.A1(new_n1385), .A2(new_n1389), .ZN(G402));
endmodule


