//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n770, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n858, new_n859, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT6), .ZN(new_n206));
  INV_X1    g005(.A(new_n205), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT5), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT82), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT80), .ZN(new_n212));
  INV_X1    g011(.A(G155gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT79), .ZN(new_n214));
  INV_X1    g013(.A(G162gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n213), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT2), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n212), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AND2_X1   g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G148gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT78), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT78), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G148gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n227), .A3(G141gat), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n224), .A2(G141gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n223), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n217), .ZN(new_n232));
  NOR2_X1   g031(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n233));
  OAI21_X1  g032(.A(G155gat), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(KEYINPUT80), .A3(KEYINPUT2), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n220), .A2(new_n231), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(G141gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n237), .A2(G148gat), .ZN(new_n238));
  OAI22_X1  g037(.A1(new_n229), .A2(new_n238), .B1(new_n219), .B2(new_n221), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n223), .A2(KEYINPUT77), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n223), .A2(KEYINPUT77), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n239), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n236), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G134gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G127gat), .ZN(new_n245));
  INV_X1    g044(.A(G127gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G134gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G120gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(G113gat), .ZN(new_n250));
  INV_X1    g049(.A(G113gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G120gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n250), .A2(new_n252), .A3(KEYINPUT68), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT68), .B1(new_n250), .B2(new_n252), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n248), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  OR2_X1    g056(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(KEYINPUT69), .A2(G113gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(G120gat), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(new_n250), .ZN(new_n261));
  INV_X1    g060(.A(new_n248), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n261), .A2(new_n254), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n211), .B1(new_n243), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT81), .ZN(new_n266));
  XNOR2_X1  g065(.A(G113gat), .B(G120gat), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT1), .B1(new_n267), .B2(KEYINPUT68), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n250), .A2(new_n252), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT68), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n262), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n245), .A2(new_n247), .A3(new_n254), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n273), .B1(new_n250), .B2(new_n260), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n266), .B1(new_n272), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n257), .A2(KEYINPUT81), .A3(new_n263), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n243), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n268), .A2(new_n271), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n274), .B1(new_n278), .B2(new_n248), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n279), .A2(KEYINPUT82), .A3(new_n242), .A4(new_n236), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G225gat), .A2(G233gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n210), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n265), .A2(new_n285), .A3(new_n280), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n243), .A2(KEYINPUT3), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT3), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n236), .A2(new_n242), .A3(new_n288), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n287), .A2(new_n289), .A3(new_n275), .A4(new_n276), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n243), .A2(new_n264), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT4), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n286), .A2(new_n290), .A3(new_n282), .A4(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n284), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n290), .A2(new_n210), .A3(new_n282), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n285), .B1(new_n265), .B2(new_n280), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n291), .A2(KEYINPUT4), .ZN(new_n297));
  NOR3_X1   g096(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n206), .B(new_n209), .C1(new_n294), .C2(new_n298), .ZN(new_n299));
  AND2_X1   g098(.A1(new_n290), .A2(new_n282), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n265), .A2(new_n280), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT4), .ZN(new_n302));
  INV_X1    g101(.A(new_n297), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n300), .A2(new_n210), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n284), .A2(new_n293), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n304), .A2(new_n305), .A3(new_n208), .A4(new_n207), .ZN(new_n306));
  XNOR2_X1  g105(.A(G197gat), .B(G204gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT22), .ZN(new_n308));
  INV_X1    g107(.A(G211gat), .ZN(new_n309));
  INV_X1    g108(.A(G218gat), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G211gat), .B(G218gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n307), .A3(new_n311), .ZN(new_n316));
  AND3_X1   g115(.A1(new_n315), .A2(KEYINPUT75), .A3(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT75), .B1(new_n315), .B2(new_n316), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G226gat), .A2(G233gat), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G169gat), .ZN(new_n322));
  INV_X1    g121(.A(G176gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT26), .ZN(new_n325));
  NAND2_X1  g124(.A1(G169gat), .A2(G176gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(G183gat), .A2(G190gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(G169gat), .A2(G176gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT26), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n327), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT27), .B(G183gat), .ZN(new_n333));
  INV_X1    g132(.A(G190gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(KEYINPUT28), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT28), .B1(new_n333), .B2(new_n334), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n332), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OR2_X1    g137(.A1(G183gat), .A2(G190gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n340));
  AND2_X1   g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT24), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n328), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT64), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT64), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n341), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n323), .A2(KEYINPUT23), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n326), .A2(KEYINPUT23), .ZN(new_n354));
  AOI22_X1  g153(.A1(new_n352), .A2(new_n353), .B1(new_n354), .B2(new_n324), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT25), .B1(new_n348), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n322), .A2(new_n323), .A3(KEYINPUT23), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT25), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n329), .B1(KEYINPUT23), .B2(new_n326), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT66), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n328), .A2(new_n360), .ZN(new_n361));
  OR2_X1    g160(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n362));
  NAND3_X1  g161(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n361), .A2(new_n362), .A3(new_n363), .A4(new_n364), .ZN(new_n365));
  AOI211_X1 g164(.A(new_n358), .B(new_n359), .C1(new_n341), .C2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n338), .B1(new_n356), .B2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n321), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n324), .ZN(new_n370));
  INV_X1    g169(.A(new_n351), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n353), .A2(new_n371), .A3(new_n349), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n339), .B(new_n340), .C1(new_n345), .C2(new_n346), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n343), .A2(KEYINPUT64), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n370), .B(new_n372), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT25), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n365), .A2(new_n341), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n359), .A2(new_n358), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n320), .B1(new_n381), .B2(new_n338), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n319), .B1(new_n369), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n321), .ZN(new_n384));
  OR2_X1    g183(.A1(new_n317), .A2(new_n318), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT29), .B1(new_n381), .B2(new_n338), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n384), .B(new_n385), .C1(new_n386), .C2(new_n321), .ZN(new_n387));
  XNOR2_X1  g186(.A(G8gat), .B(G36gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(G64gat), .B(G92gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n391), .A2(KEYINPUT37), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n392), .B(KEYINPUT38), .Z(new_n393));
  AND3_X1   g192(.A1(new_n383), .A2(new_n387), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n383), .A2(new_n387), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n390), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n299), .A2(new_n306), .A3(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G78gat), .B(G106gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT31), .B(G50gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(G22gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n289), .A2(new_n368), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(KEYINPUT83), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT83), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n289), .A2(new_n406), .A3(new_n368), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n385), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G228gat), .A2(G233gat), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n243), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n315), .A2(new_n316), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT3), .B1(new_n412), .B2(new_n368), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n410), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n408), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n404), .A2(new_n385), .ZN(new_n417));
  INV_X1    g216(.A(new_n413), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(new_n243), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(new_n409), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n403), .B1(new_n416), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n319), .B1(new_n404), .B2(KEYINPUT83), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n414), .B1(new_n423), .B2(new_n407), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n410), .B1(new_n417), .B2(new_n419), .ZN(new_n425));
  NOR3_X1   g224(.A1(new_n424), .A2(new_n425), .A3(G22gat), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n402), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n416), .A2(new_n421), .A3(new_n403), .ZN(new_n428));
  OAI21_X1  g227(.A(G22gat), .B1(new_n424), .B2(new_n425), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n429), .A3(new_n401), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n398), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT40), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n302), .A2(new_n303), .A3(new_n290), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT39), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n283), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n205), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n265), .A2(new_n277), .A3(new_n280), .A4(new_n282), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT39), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n439), .B1(new_n434), .B2(new_n283), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n433), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n383), .A2(new_n390), .A3(new_n387), .ZN(new_n442));
  AND2_X1   g241(.A1(new_n442), .A2(KEYINPUT76), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT76), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n383), .A2(new_n387), .A3(new_n444), .A4(new_n390), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT30), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n447), .B1(new_n395), .B2(new_n391), .ZN(new_n448));
  AOI211_X1 g247(.A(KEYINPUT30), .B(new_n390), .C1(new_n383), .C2(new_n387), .ZN(new_n449));
  OAI22_X1  g248(.A1(new_n443), .A2(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n283), .ZN(new_n451));
  INV_X1    g250(.A(new_n439), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n453), .A2(KEYINPUT40), .A3(new_n205), .A4(new_n436), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n304), .A2(new_n305), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n207), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n441), .A2(new_n450), .A3(new_n454), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n395), .A2(new_n391), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT30), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n395), .A2(new_n447), .A3(new_n391), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n442), .A2(KEYINPUT76), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n459), .A2(new_n460), .B1(new_n461), .B2(new_n445), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n455), .A2(new_n206), .A3(new_n209), .ZN(new_n463));
  INV_X1    g262(.A(new_n306), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(new_n431), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n432), .A2(new_n457), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT36), .ZN(new_n468));
  AOI22_X1  g267(.A1(new_n375), .A2(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n469));
  INV_X1    g268(.A(new_n337), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n331), .B1(new_n470), .B2(new_n335), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n279), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n264), .B(new_n338), .C1(new_n356), .C2(new_n366), .ZN(new_n473));
  INV_X1    g272(.A(G227gat), .ZN(new_n474));
  INV_X1    g273(.A(G233gat), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n472), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  XOR2_X1   g276(.A(G71gat), .B(G99gat), .Z(new_n478));
  XNOR2_X1  g277(.A(G15gat), .B(G43gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  XNOR2_X1  g279(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n482), .A2(KEYINPUT71), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n477), .A2(KEYINPUT32), .A3(new_n483), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n472), .A2(new_n473), .A3(new_n476), .A4(new_n480), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT71), .B1(new_n485), .B2(new_n482), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n477), .A2(KEYINPUT32), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n484), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n489));
  INV_X1    g288(.A(new_n476), .ZN(new_n490));
  XNOR2_X1  g289(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n491), .B1(new_n489), .B2(new_n490), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n488), .A2(KEYINPUT73), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(KEYINPUT73), .B1(new_n488), .B2(new_n494), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n477), .A2(KEYINPUT32), .A3(new_n483), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n485), .A2(new_n482), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT71), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n477), .A2(KEYINPUT32), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n492), .A2(new_n493), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(KEYINPUT74), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT74), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n506), .B1(new_n488), .B2(new_n494), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n468), .B1(new_n497), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT73), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n510), .B1(new_n503), .B2(new_n504), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n488), .A2(KEYINPUT73), .A3(new_n494), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n503), .A2(new_n504), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(KEYINPUT36), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n509), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n513), .A2(new_n431), .A3(new_n514), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT35), .B1(new_n517), .B2(new_n465), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n497), .A2(new_n508), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n450), .B1(new_n306), .B2(new_n299), .ZN(new_n520));
  XOR2_X1   g319(.A(KEYINPUT84), .B(KEYINPUT35), .Z(new_n521));
  AOI21_X1  g320(.A(new_n521), .B1(new_n427), .B2(new_n430), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n467), .A2(new_n516), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT88), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G1gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n525), .A2(new_n526), .A3(G1gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT16), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n529), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(G8gat), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(G43gat), .B(G50gat), .Z(new_n536));
  INV_X1    g335(.A(KEYINPUT15), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT86), .B(G36gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(G29gat), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(G29gat), .A2(G36gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT14), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n538), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(KEYINPUT87), .ZN(new_n545));
  INV_X1    g344(.A(new_n538), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n536), .A2(new_n537), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(new_n540), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n544), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT17), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI211_X1 g350(.A(KEYINPUT17), .B(new_n544), .C1(new_n545), .C2(new_n548), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n535), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(G229gat), .A2(G233gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n534), .A2(new_n549), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT18), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n553), .A2(KEYINPUT18), .A3(new_n554), .A4(new_n555), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n534), .B(new_n549), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n554), .B(KEYINPUT13), .Z(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n558), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G113gat), .B(G141gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(G197gat), .ZN(new_n565));
  XOR2_X1   g364(.A(KEYINPUT11), .B(G169gat), .Z(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(KEYINPUT12), .ZN(new_n568));
  AND3_X1   g367(.A1(new_n563), .A2(KEYINPUT85), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n568), .B1(new_n563), .B2(KEYINPUT85), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n524), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(G230gat), .A2(G233gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(G71gat), .A2(G78gat), .ZN(new_n575));
  NOR2_X1   g374(.A1(G71gat), .A2(G78gat), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT9), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n575), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(KEYINPUT89), .B(G57gat), .Z(new_n580));
  AND2_X1   g379(.A1(new_n580), .A2(G64gat), .ZN(new_n581));
  INV_X1    g380(.A(G57gat), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n582), .A2(G64gat), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n579), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G57gat), .B(G64gat), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n575), .B(new_n577), .C1(new_n585), .C2(new_n578), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(KEYINPUT92), .A2(G85gat), .A3(G92gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT7), .ZN(new_n589));
  XOR2_X1   g388(.A(G99gat), .B(G106gat), .Z(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G99gat), .A2(G106gat), .ZN(new_n592));
  INV_X1    g391(.A(G85gat), .ZN(new_n593));
  INV_X1    g392(.A(G92gat), .ZN(new_n594));
  AOI22_X1  g393(.A1(KEYINPUT8), .A2(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  AND3_X1   g394(.A1(new_n589), .A2(new_n591), .A3(new_n595), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n591), .B1(new_n589), .B2(new_n595), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n587), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n586), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n600), .B1(new_n596), .B2(new_n597), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n599), .A2(KEYINPUT94), .A3(new_n601), .ZN(new_n602));
  OR3_X1    g401(.A1(new_n587), .A2(new_n598), .A3(KEYINPUT94), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT10), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT10), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n574), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n574), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n602), .A2(new_n603), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT95), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT96), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT96), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n610), .A2(KEYINPUT95), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G120gat), .B(G148gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(G176gat), .B(G204gat), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n615), .B(new_n616), .Z(new_n617));
  NAND3_X1  g416(.A1(new_n612), .A2(new_n614), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n617), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n613), .B1(new_n610), .B2(KEYINPUT95), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT95), .ZN(new_n621));
  AOI211_X1 g420(.A(new_n621), .B(KEYINPUT96), .C1(new_n607), .C2(new_n609), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n619), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n587), .A2(KEYINPUT21), .ZN(new_n625));
  AND2_X1   g424(.A1(G231gat), .A2(G233gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(new_n246), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n534), .B1(KEYINPUT21), .B2(new_n587), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n627), .B(G127gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n629), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT90), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G155gat), .ZN(new_n636));
  XOR2_X1   g435(.A(G183gat), .B(G211gat), .Z(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n630), .A2(new_n633), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n638), .B1(new_n630), .B2(new_n633), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT91), .ZN(new_n643));
  XNOR2_X1  g442(.A(G134gat), .B(G162gat), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G190gat), .B(G218gat), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n646), .A2(KEYINPUT93), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n551), .B(new_n552), .C1(new_n596), .C2(new_n597), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(KEYINPUT93), .ZN(new_n650));
  NAND3_X1  g449(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n652), .B1(new_n549), .B2(new_n598), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n648), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n649), .A2(new_n648), .A3(new_n653), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n645), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n655), .A2(new_n645), .A3(new_n656), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR3_X1   g459(.A1(new_n624), .A2(new_n641), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n573), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n463), .A2(new_n464), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT97), .B(G1gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(G1324gat));
  INV_X1    g466(.A(new_n662), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n450), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n669), .A2(G8gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(KEYINPUT16), .B(G8gat), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT42), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n673), .B1(KEYINPUT42), .B2(new_n672), .ZN(G1325gat));
  XNOR2_X1  g473(.A(new_n516), .B(KEYINPUT98), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(G15gat), .B1(new_n662), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n519), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n678), .A2(G15gat), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n677), .B1(new_n662), .B2(new_n679), .ZN(G1326gat));
  NAND2_X1  g479(.A1(new_n668), .A2(new_n466), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT99), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT43), .B(G22gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1327gat));
  INV_X1    g483(.A(new_n624), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n641), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(new_n572), .ZN(new_n687));
  INV_X1    g486(.A(new_n660), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n524), .A2(new_n688), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(G29gat), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n690), .A2(new_n691), .A3(new_n663), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT45), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n695), .B1(new_n524), .B2(new_n688), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n457), .A2(new_n431), .A3(new_n398), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n465), .A2(new_n466), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n516), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n518), .A2(new_n523), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(KEYINPUT44), .A3(new_n660), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n696), .A2(new_n687), .A3(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT100), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n696), .A2(new_n702), .A3(new_n687), .A4(KEYINPUT100), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n694), .B1(new_n707), .B2(new_n664), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(G29gat), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n707), .A2(new_n694), .A3(new_n664), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n693), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT102), .Z(G1328gat));
  NOR2_X1   g511(.A1(new_n462), .A2(new_n539), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n690), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g513(.A(new_n714), .B(KEYINPUT46), .Z(new_n715));
  OAI21_X1  g514(.A(new_n539), .B1(new_n707), .B2(new_n462), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(G1329gat));
  INV_X1    g516(.A(G43gat), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n690), .A2(new_n718), .A3(new_n519), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n696), .A2(new_n702), .ZN(new_n720));
  INV_X1    g519(.A(new_n516), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n721), .A3(new_n687), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(KEYINPUT104), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(G43gat), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n722), .A2(KEYINPUT104), .ZN(new_n725));
  OAI211_X1 g524(.A(KEYINPUT47), .B(new_n719), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  XOR2_X1   g525(.A(new_n719), .B(KEYINPUT103), .Z(new_n727));
  NAND3_X1  g526(.A1(new_n705), .A2(new_n675), .A3(new_n706), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n727), .B1(new_n728), .B2(G43gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n726), .B1(new_n729), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR4_X1   g529(.A1(new_n686), .A2(G50gat), .A3(new_n431), .A4(new_n688), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n731), .A2(new_n573), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G50gat), .B1(new_n703), .B2(new_n431), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(KEYINPUT48), .A3(new_n734), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT107), .Z(new_n736));
  NAND3_X1  g535(.A1(new_n705), .A2(new_n466), .A3(new_n706), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G50gat), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT105), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n732), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n737), .A2(KEYINPUT105), .A3(G50gat), .ZN(new_n741));
  AOI211_X1 g540(.A(KEYINPUT106), .B(KEYINPUT48), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n738), .A2(new_n739), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(new_n741), .A3(new_n733), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT48), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n743), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n736), .B1(new_n742), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT108), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT108), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n750), .B(new_n736), .C1(new_n742), .C2(new_n747), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(G1331gat));
  INV_X1    g551(.A(new_n641), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n688), .ZN(new_n754));
  NOR4_X1   g553(.A1(new_n524), .A2(new_n754), .A3(new_n685), .A4(new_n571), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n663), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT109), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(new_n580), .ZN(G1332gat));
  AOI21_X1  g557(.A(new_n462), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n759), .B(KEYINPUT110), .Z(new_n760));
  NAND2_X1  g559(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n762));
  XOR2_X1   g561(.A(new_n761), .B(new_n762), .Z(G1333gat));
  NAND3_X1  g562(.A1(new_n755), .A2(G71gat), .A3(new_n675), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT111), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n519), .B(KEYINPUT112), .Z(new_n766));
  AND2_X1   g565(.A1(new_n755), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(G71gat), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g568(.A1(new_n755), .A2(new_n466), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g570(.A1(new_n685), .A2(new_n571), .A3(new_n753), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n720), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(G85gat), .B1(new_n773), .B2(new_n664), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n689), .A2(new_n572), .A3(new_n641), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT51), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT113), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT113), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT51), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n775), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n777), .A2(new_n624), .A3(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n663), .A2(new_n593), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n774), .B1(new_n781), .B2(new_n782), .ZN(G1336gat));
  OAI21_X1  g582(.A(G92gat), .B1(new_n773), .B2(new_n462), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n624), .A2(new_n594), .A3(new_n450), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n776), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT52), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n781), .A2(G92gat), .A3(new_n462), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n784), .A2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n787), .B1(new_n788), .B2(new_n790), .ZN(G1337gat));
  OR2_X1    g590(.A1(new_n678), .A2(G99gat), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n720), .A2(new_n675), .A3(new_n772), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G99gat), .ZN(new_n797));
  OAI22_X1  g596(.A1(new_n781), .A2(new_n792), .B1(new_n795), .B2(new_n797), .ZN(G1338gat));
  NOR2_X1   g597(.A1(new_n773), .A2(new_n431), .ZN(new_n799));
  INV_X1    g598(.A(G106gat), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n624), .A2(new_n800), .A3(new_n466), .ZN(new_n801));
  OAI22_X1  g600(.A1(new_n799), .A2(new_n800), .B1(new_n776), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT53), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n777), .A2(new_n780), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n804), .B1(new_n805), .B2(new_n801), .ZN(new_n806));
  OAI21_X1  g605(.A(G106gat), .B1(new_n799), .B2(KEYINPUT115), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n807), .B1(KEYINPUT115), .B2(new_n799), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n803), .B1(new_n806), .B2(new_n808), .ZN(G1339gat));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n810), .B(new_n574), .C1(new_n604), .C2(new_n606), .ZN(new_n811));
  AND2_X1   g610(.A1(new_n811), .A2(new_n619), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n602), .A2(new_n603), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n606), .B1(new_n813), .B2(new_n605), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n608), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n815), .A2(KEYINPUT54), .A3(new_n607), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n607), .A2(new_n609), .A3(new_n617), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n812), .A2(new_n816), .A3(KEYINPUT55), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n571), .A2(new_n819), .A3(new_n820), .A4(new_n821), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n558), .A2(new_n559), .A3(new_n562), .A4(new_n568), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n560), .A2(new_n561), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n554), .B1(new_n553), .B2(new_n555), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n567), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n618), .A2(new_n623), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n660), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n660), .A2(new_n827), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n821), .A2(new_n820), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT55), .B1(new_n812), .B2(new_n816), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n641), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n661), .A2(new_n572), .ZN(new_n835));
  AND3_X1   g634(.A1(new_n834), .A2(new_n835), .A3(KEYINPUT116), .ZN(new_n836));
  AOI21_X1  g635(.A(KEYINPUT116), .B1(new_n834), .B2(new_n835), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n663), .A2(new_n462), .ZN(new_n840));
  NOR4_X1   g639(.A1(new_n839), .A2(new_n678), .A3(new_n466), .A4(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G113gat), .B1(new_n842), .B2(new_n572), .ZN(new_n843));
  NOR3_X1   g642(.A1(new_n836), .A2(new_n837), .A3(new_n664), .ZN(new_n844));
  INV_X1    g643(.A(new_n517), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT117), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n844), .A2(KEYINPUT117), .A3(new_n845), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n450), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n571), .A2(new_n258), .A3(new_n259), .ZN(new_n851));
  XNOR2_X1  g650(.A(new_n851), .B(KEYINPUT118), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n843), .A2(new_n853), .ZN(G1340gat));
  AOI21_X1  g653(.A(G120gat), .B1(new_n850), .B2(new_n624), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n842), .A2(new_n249), .A3(new_n685), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(G1341gat));
  NAND3_X1  g656(.A1(new_n850), .A2(new_n246), .A3(new_n753), .ZN(new_n858));
  OAI21_X1  g657(.A(G127gat), .B1(new_n842), .B2(new_n641), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1342gat));
  AOI21_X1  g659(.A(new_n244), .B1(new_n841), .B2(new_n660), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n660), .A2(new_n244), .ZN(new_n862));
  AOI211_X1 g661(.A(new_n450), .B(new_n862), .C1(new_n848), .C2(new_n849), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT56), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n863), .A2(new_n864), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(KEYINPUT119), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT119), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n863), .A2(new_n868), .A3(new_n864), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n865), .B1(new_n867), .B2(new_n869), .ZN(G1343gat));
  NAND4_X1  g669(.A1(new_n844), .A2(new_n462), .A3(new_n466), .A4(new_n676), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n237), .B1(new_n871), .B2(new_n572), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n721), .A2(new_n840), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT120), .Z(new_n874));
  AOI21_X1  g673(.A(KEYINPUT57), .B1(new_n838), .B2(new_n466), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n466), .A2(KEYINPUT57), .ZN(new_n876));
  OAI21_X1  g675(.A(KEYINPUT121), .B1(new_n831), .B2(new_n832), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n819), .A2(new_n878), .A3(new_n820), .A4(new_n821), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n877), .A2(new_n571), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n660), .B1(new_n880), .B2(new_n828), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n641), .B1(new_n881), .B2(new_n833), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT122), .ZN(new_n883));
  AOI22_X1  g682(.A1(new_n882), .A2(new_n883), .B1(new_n572), .B2(new_n661), .ZN(new_n884));
  OAI211_X1 g683(.A(KEYINPUT122), .B(new_n641), .C1(new_n881), .C2(new_n833), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n876), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n874), .B1(new_n875), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n571), .A2(G141gat), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n872), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  XOR2_X1   g688(.A(new_n889), .B(KEYINPUT58), .Z(G1344gat));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n838), .A2(KEYINPUT57), .A3(new_n466), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n882), .A2(new_n835), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n466), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n874), .A2(new_n624), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n891), .B1(new_n899), .B2(G148gat), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n624), .B(new_n874), .C1(new_n875), .C2(new_n886), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT59), .B1(new_n225), .B2(new_n227), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n901), .A2(KEYINPUT123), .A3(new_n902), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n900), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n225), .A2(new_n227), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n871), .A2(new_n908), .A3(new_n685), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT124), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT124), .ZN(new_n911));
  INV_X1    g710(.A(new_n909), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n901), .A2(KEYINPUT123), .A3(new_n902), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT123), .B1(new_n901), .B2(new_n902), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n911), .B(new_n912), .C1(new_n915), .C2(new_n900), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n910), .A2(new_n916), .ZN(G1345gat));
  OAI21_X1  g716(.A(G155gat), .B1(new_n887), .B2(new_n641), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n753), .A2(new_n213), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n871), .B2(new_n919), .ZN(G1346gat));
  NAND2_X1  g719(.A1(new_n216), .A2(new_n217), .ZN(new_n921));
  OR3_X1    g720(.A1(new_n871), .A2(new_n921), .A3(new_n688), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n887), .A2(new_n688), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n923), .A2(KEYINPUT125), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n921), .B1(new_n923), .B2(KEYINPUT125), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(G1347gat));
  NOR2_X1   g725(.A1(new_n663), .A2(new_n462), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n838), .A2(new_n431), .A3(new_n766), .A4(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G169gat), .B1(new_n928), .B2(new_n572), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n839), .A2(new_n663), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(new_n450), .A3(new_n845), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n571), .A2(new_n352), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1348gat));
  OAI21_X1  g732(.A(G176gat), .B1(new_n928), .B2(new_n685), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n624), .A2(new_n323), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n934), .B1(new_n931), .B2(new_n935), .ZN(G1349gat));
  OAI21_X1  g735(.A(G183gat), .B1(new_n928), .B2(new_n641), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n753), .A2(new_n333), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n931), .B2(new_n938), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g739(.A(G190gat), .B1(new_n928), .B2(new_n688), .ZN(new_n941));
  OR2_X1    g740(.A1(new_n941), .A2(KEYINPUT126), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(KEYINPUT126), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n942), .A2(KEYINPUT61), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n660), .A2(new_n334), .ZN(new_n945));
  OAI221_X1 g744(.A(new_n944), .B1(KEYINPUT61), .B2(new_n943), .C1(new_n931), .C2(new_n945), .ZN(G1351gat));
  NOR3_X1   g745(.A1(new_n675), .A2(new_n462), .A3(new_n431), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n930), .A2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(G197gat), .B1(new_n949), .B2(new_n571), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n897), .A2(new_n676), .A3(new_n927), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n571), .A2(G197gat), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(G1352gat));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n624), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(G204gat), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n685), .A2(G204gat), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(KEYINPUT62), .B1(new_n948), .B2(new_n957), .ZN(new_n958));
  OR3_X1    g757(.A1(new_n948), .A2(KEYINPUT62), .A3(new_n957), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n955), .A2(new_n958), .A3(new_n959), .ZN(G1353gat));
  NAND3_X1  g759(.A1(new_n949), .A2(new_n309), .A3(new_n753), .ZN(new_n961));
  OAI21_X1  g760(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n962), .B1(new_n951), .B2(new_n753), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n963), .A2(KEYINPUT127), .A3(KEYINPUT63), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n963), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(G1354gat));
  NAND3_X1  g765(.A1(new_n949), .A2(new_n310), .A3(new_n660), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n951), .A2(new_n660), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n967), .B1(new_n968), .B2(new_n310), .ZN(G1355gat));
endmodule


