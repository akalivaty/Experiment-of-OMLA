//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT76), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207));
  INV_X1    g006(.A(G211gat), .ZN(new_n208));
  INV_X1    g007(.A(G218gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n207), .B1(KEYINPUT22), .B2(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(G211gat), .B(G218gat), .Z(new_n212));
  XNOR2_X1  g011(.A(new_n211), .B(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G226gat), .A2(G233gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G183gat), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT24), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n219), .A2(G183gat), .A3(G190gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(KEYINPUT66), .B(G183gat), .Z(new_n222));
  OAI21_X1  g021(.A(new_n221), .B1(new_n222), .B2(G190gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT23), .ZN(new_n225));
  INV_X1    g024(.A(G169gat), .ZN(new_n226));
  INV_X1    g025(.A(G176gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT23), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n223), .A2(KEYINPUT25), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT25), .ZN(new_n232));
  OR2_X1    g031(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n233), .A2(KEYINPUT23), .A3(new_n227), .A4(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n229), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n218), .A2(new_n220), .B1(new_n216), .B2(new_n217), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n232), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n231), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT26), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n228), .A2(new_n240), .A3(new_n224), .ZN(new_n241));
  NOR2_X1   g040(.A1(G169gat), .A2(G176gat), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n242), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT28), .ZN(new_n245));
  OAI21_X1  g044(.A(KEYINPUT67), .B1(new_n216), .B2(KEYINPUT27), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT27), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n248), .A3(G183gat), .ZN(new_n249));
  AND4_X1   g048(.A1(new_n245), .A2(new_n246), .A3(new_n249), .A4(new_n217), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT66), .B(G183gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(KEYINPUT27), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n244), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT27), .B(G183gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT68), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT68), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n216), .A2(KEYINPUT27), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n248), .A2(G183gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(G190gat), .B1(new_n255), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n253), .B1(new_n245), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n239), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT29), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n215), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n255), .A2(new_n259), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT28), .B1(new_n265), .B2(G190gat), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n266), .A2(new_n253), .B1(new_n231), .B2(new_n238), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n267), .A2(new_n214), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT75), .B1(new_n264), .B2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n214), .B1(new_n267), .B2(KEYINPUT29), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT75), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n213), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n262), .A2(new_n215), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n213), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n206), .B1(new_n273), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n271), .B1(new_n270), .B2(new_n274), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n264), .A2(KEYINPUT75), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n276), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n275), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n213), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(new_n283), .A3(new_n205), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n278), .A2(new_n284), .A3(KEYINPUT30), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n273), .A2(new_n277), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT30), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(new_n287), .A3(new_n205), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT2), .ZN(new_n289));
  INV_X1    g088(.A(G155gat), .ZN(new_n290));
  INV_X1    g089(.A(G162gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293));
  INV_X1    g092(.A(G141gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n294), .A2(G148gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT77), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n292), .A2(new_n293), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G141gat), .B(G148gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT77), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G148gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(G141gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n289), .B1(new_n295), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n290), .A2(new_n291), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n304), .A2(new_n293), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n300), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT3), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n297), .A2(new_n299), .B1(new_n303), .B2(new_n305), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT3), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT69), .ZN(new_n312));
  INV_X1    g111(.A(G113gat), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n312), .B1(new_n313), .B2(G120gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT70), .ZN(new_n315));
  INV_X1    g114(.A(G120gat), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n315), .B1(new_n316), .B2(G113gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n313), .A2(KEYINPUT70), .A3(G120gat), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n314), .A2(new_n317), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT1), .ZN(new_n321));
  XNOR2_X1  g120(.A(G127gat), .B(G134gat), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n313), .A2(G120gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n316), .A2(G113gat), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n321), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n322), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n323), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n308), .A2(new_n311), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT4), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(new_n329), .B2(new_n307), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n323), .A2(new_n328), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n333), .A2(KEYINPUT4), .A3(new_n309), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n330), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G225gat), .A2(G233gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n329), .A2(new_n307), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n328), .A2(new_n323), .B1(new_n300), .B2(new_n306), .ZN(new_n340));
  OR2_X1    g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n338), .B(KEYINPUT39), .C1(new_n337), .C2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G1gat), .B(G29gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n343), .B(KEYINPUT0), .ZN(new_n344));
  XNOR2_X1  g143(.A(G57gat), .B(G85gat), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n344), .B(new_n345), .Z(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT83), .B(KEYINPUT39), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n335), .A2(new_n337), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n342), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT40), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n330), .A2(new_n334), .A3(new_n336), .A4(new_n332), .ZN(new_n352));
  OR2_X1    g151(.A1(new_n352), .A2(KEYINPUT5), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n337), .B1(new_n339), .B2(new_n340), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g155(.A(KEYINPUT78), .B(new_n337), .C1(new_n339), .C2(new_n340), .ZN(new_n357));
  NAND4_X1  g156(.A1(new_n356), .A2(new_n352), .A3(KEYINPUT5), .A4(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n346), .B1(new_n353), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n359), .B1(new_n349), .B2(new_n350), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n285), .A2(new_n288), .A3(new_n351), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(G228gat), .A2(G233gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n213), .A2(new_n263), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n309), .B1(new_n363), .B2(new_n310), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n213), .B1(new_n311), .B2(new_n263), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n362), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  OR2_X1    g165(.A1(new_n363), .A2(KEYINPUT81), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT3), .B1(new_n363), .B2(KEYINPUT81), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n309), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OR2_X1    g168(.A1(new_n365), .A2(new_n362), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n366), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G78gat), .B(G106gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(KEYINPUT31), .B(G50gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT82), .ZN(new_n375));
  INV_X1    g174(.A(G22gat), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n377), .B1(new_n376), .B2(new_n374), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n371), .B(new_n378), .ZN(new_n379));
  AND2_X1   g178(.A1(new_n361), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT85), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT37), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n286), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n281), .A2(new_n382), .A3(new_n283), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT85), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT84), .B1(new_n282), .B2(new_n213), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n269), .A2(new_n213), .A3(new_n272), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT84), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n275), .A2(new_n389), .A3(new_n276), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n387), .A2(new_n388), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT38), .B1(new_n391), .B2(KEYINPUT37), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n386), .A2(new_n206), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n353), .A2(new_n358), .ZN(new_n394));
  INV_X1    g193(.A(new_n346), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n353), .A2(new_n358), .A3(new_n346), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT79), .B(KEYINPUT6), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n398), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n359), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n402), .B1(new_n286), .B2(new_n205), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n393), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT38), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n205), .B1(new_n383), .B2(new_n385), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT37), .B1(new_n273), .B2(new_n277), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n380), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(G15gat), .B(G43gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(KEYINPUT72), .ZN(new_n411));
  XOR2_X1   g210(.A(G71gat), .B(G99gat), .Z(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(G227gat), .A2(G233gat), .ZN(new_n414));
  XOR2_X1   g213(.A(new_n414), .B(KEYINPUT64), .Z(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n333), .B1(new_n239), .B2(new_n261), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT71), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n239), .A2(new_n261), .A3(new_n333), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n239), .A2(new_n261), .A3(KEYINPUT71), .A4(new_n333), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n416), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT32), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n423), .A2(KEYINPUT33), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n413), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n419), .A2(new_n418), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n262), .A2(new_n329), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n426), .A2(new_n421), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n415), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n423), .B1(new_n413), .B2(KEYINPUT33), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT73), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT73), .ZN(new_n432));
  INV_X1    g231(.A(new_n430), .ZN(new_n433));
  AOI211_X1 g232(.A(new_n432), .B(new_n433), .C1(new_n428), .C2(new_n415), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n425), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n426), .A2(new_n427), .A3(new_n416), .A4(new_n421), .ZN(new_n436));
  XNOR2_X1  g235(.A(new_n436), .B(KEYINPUT34), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n436), .B(KEYINPUT34), .Z(new_n439));
  OAI211_X1 g238(.A(new_n439), .B(new_n425), .C1(new_n431), .C2(new_n434), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT36), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT74), .ZN(new_n443));
  OR2_X1    g242(.A1(new_n442), .A2(KEYINPUT74), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n438), .A2(new_n440), .A3(KEYINPUT74), .A4(new_n442), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n399), .A2(KEYINPUT80), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT80), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n396), .A2(new_n449), .A3(new_n397), .A4(new_n398), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n448), .A2(new_n450), .A3(new_n401), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n285), .A2(new_n288), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n379), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n409), .A2(new_n447), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n438), .A2(new_n440), .A3(new_n379), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT35), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n441), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT35), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n402), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n459), .A2(new_n462), .A3(new_n452), .A4(new_n379), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n456), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(G71gat), .A2(G78gat), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT9), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OR2_X1    g267(.A1(G57gat), .A2(G64gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(G57gat), .A2(G64gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G71gat), .B(G78gat), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT92), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n473), .B1(G71gat), .B2(G78gat), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n471), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n472), .B1(new_n471), .B2(new_n474), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT21), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(G231gat), .A2(G233gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(G127gat), .ZN(new_n482));
  XOR2_X1   g281(.A(G183gat), .B(G211gat), .Z(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  OR2_X1    g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n482), .A2(new_n484), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n376), .A2(G15gat), .ZN(new_n488));
  INV_X1    g287(.A(G15gat), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(G22gat), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT16), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n488), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(G1gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(G8gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(G15gat), .B(G22gat), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n495), .B1(new_n496), .B2(KEYINPUT89), .ZN(new_n497));
  AND4_X1   g296(.A1(KEYINPUT89), .A2(new_n488), .A3(new_n490), .A4(new_n495), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n488), .A2(new_n490), .A3(KEYINPUT89), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(G8gat), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n496), .A2(KEYINPUT89), .A3(new_n495), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n501), .A2(new_n502), .A3(new_n493), .A4(new_n492), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n504), .B1(new_n477), .B2(new_n478), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n505), .B(KEYINPUT93), .Z(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(new_n290), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n506), .B(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n487), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n487), .A2(new_n510), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G43gat), .B(G50gat), .ZN(new_n516));
  INV_X1    g315(.A(G29gat), .ZN(new_n517));
  INV_X1    g316(.A(G36gat), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT14), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT14), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n520), .B1(G29gat), .B2(G36gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n517), .A2(new_n518), .ZN(new_n523));
  OAI211_X1 g322(.A(KEYINPUT15), .B(new_n516), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(KEYINPUT87), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT87), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n519), .A2(new_n521), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT15), .ZN(new_n529));
  INV_X1    g328(.A(G43gat), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n530), .A2(G50gat), .ZN(new_n531));
  INV_X1    g330(.A(G50gat), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n532), .A2(G43gat), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n529), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n523), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n532), .A2(G43gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n530), .A2(G50gat), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(new_n537), .A3(KEYINPUT15), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n534), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  OAI211_X1 g338(.A(KEYINPUT17), .B(new_n524), .C1(new_n528), .C2(new_n539), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n540), .A2(new_n504), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n523), .B1(new_n516), .B2(KEYINPUT15), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n542), .A2(new_n525), .A3(new_n534), .A4(new_n527), .ZN(new_n543));
  AOI211_X1 g342(.A(KEYINPUT88), .B(KEYINPUT17), .C1(new_n543), .C2(new_n524), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT88), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n524), .B1(new_n528), .B2(new_n539), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n541), .B1(new_n544), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n546), .A2(new_n503), .A3(new_n499), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  XOR2_X1   g351(.A(KEYINPUT90), .B(KEYINPUT18), .Z(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n549), .A2(KEYINPUT18), .A3(new_n550), .A4(new_n551), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n519), .A2(new_n521), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n538), .B1(new_n556), .B2(new_n535), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n538), .A2(new_n535), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n516), .A2(KEYINPUT15), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n519), .A2(new_n521), .A3(new_n526), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n526), .B1(new_n519), .B2(new_n521), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n557), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n504), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n551), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(new_n550), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n554), .A2(new_n555), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G113gat), .B(G141gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G169gat), .B(G197gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT12), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n570), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n554), .A2(new_n555), .A3(new_n569), .A4(new_n576), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G134gat), .B(G162gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT94), .ZN(new_n583));
  AND2_X1   g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(KEYINPUT41), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n583), .B(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(G85gat), .A2(G92gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT7), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT7), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n592), .A2(G85gat), .A3(G92gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT95), .ZN(new_n595));
  INV_X1    g394(.A(G85gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(G92gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(KEYINPUT95), .A2(G85gat), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(G99gat), .ZN(new_n601));
  INV_X1    g400(.A(G106gat), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT8), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n594), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G99gat), .B(G106gat), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n594), .A2(new_n600), .A3(new_n605), .A4(new_n603), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n540), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n610), .B1(new_n544), .B2(new_n548), .ZN(new_n611));
  INV_X1    g410(.A(new_n609), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n612), .A2(new_n546), .B1(KEYINPUT41), .B2(new_n584), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n589), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n587), .B1(new_n614), .B2(KEYINPUT96), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n540), .A2(new_n609), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT88), .B1(new_n564), .B2(KEYINPUT17), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n546), .A2(new_n545), .A3(new_n547), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n613), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n588), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT97), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n611), .A2(new_n589), .A3(new_n613), .ZN(new_n623));
  AND3_X1   g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n622), .B1(new_n621), .B2(new_n623), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n615), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n619), .A2(new_n620), .A3(new_n588), .ZN(new_n627));
  OAI21_X1  g426(.A(KEYINPUT97), .B1(new_n627), .B2(new_n614), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT96), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n586), .B1(new_n621), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n628), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n609), .A2(new_n477), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  OAI211_X1 g434(.A(new_n607), .B(new_n608), .C1(new_n476), .C2(new_n475), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n477), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n612), .A2(new_n638), .A3(KEYINPUT10), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(G176gat), .B(G204gat), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n643), .B(new_n644), .Z(new_n645));
  NAND2_X1  g444(.A1(new_n634), .A2(new_n636), .ZN(new_n646));
  INV_X1    g445(.A(new_n641), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT98), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n641), .B1(new_n634), .B2(new_n636), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT98), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AND4_X1   g451(.A1(new_n642), .A2(new_n645), .A3(new_n649), .A4(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n645), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n647), .B1(new_n637), .B2(new_n639), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n655), .B1(new_n656), .B2(new_n650), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NOR4_X1   g457(.A1(new_n515), .A2(new_n581), .A3(new_n633), .A4(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n465), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n451), .B(KEYINPUT99), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(new_n493), .ZN(G1324gat));
  INV_X1    g463(.A(new_n452), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT16), .B(G8gat), .Z(new_n666));
  NAND4_X1  g465(.A1(new_n465), .A2(new_n665), .A3(new_n659), .A4(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT42), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT100), .ZN(new_n670));
  OAI21_X1  g469(.A(G8gat), .B1(new_n660), .B2(new_n452), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n670), .B(new_n671), .C1(new_n668), .C2(new_n667), .ZN(G1325gat));
  OAI21_X1  g471(.A(G15gat), .B1(new_n660), .B2(new_n447), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n459), .A2(new_n489), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n673), .B1(new_n660), .B2(new_n674), .ZN(G1326gat));
  NOR2_X1   g474(.A1(new_n660), .A2(new_n379), .ZN(new_n676));
  XOR2_X1   g475(.A(KEYINPUT43), .B(G22gat), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(G1327gat));
  NOR3_X1   g477(.A1(new_n514), .A2(new_n581), .A3(new_n658), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n465), .A2(new_n633), .A3(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n680), .A2(new_n517), .A3(new_n661), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT45), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n465), .A2(KEYINPUT44), .A3(new_n633), .ZN(new_n683));
  INV_X1    g482(.A(new_n633), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n685));
  AOI22_X1  g484(.A1(new_n399), .A2(KEYINPUT80), .B1(new_n400), .B2(new_n359), .ZN(new_n686));
  AOI22_X1  g485(.A1(new_n686), .A2(new_n450), .B1(new_n288), .B2(new_n285), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n438), .A2(new_n440), .A3(new_n379), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n460), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n452), .A2(new_n379), .A3(new_n438), .A4(new_n440), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n690), .A2(new_n461), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n685), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n458), .A2(new_n463), .A3(KEYINPUT102), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT101), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n695), .B1(new_n687), .B2(new_n379), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n453), .A2(KEYINPUT101), .A3(new_n454), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n409), .A2(new_n447), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n684), .B1(new_n694), .B2(new_n698), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n683), .B(new_n679), .C1(new_n699), .C2(KEYINPUT44), .ZN(new_n700));
  OAI21_X1  g499(.A(G29gat), .B1(new_n700), .B2(new_n662), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n682), .A2(new_n701), .ZN(G1328gat));
  NAND3_X1  g501(.A1(new_n680), .A2(new_n518), .A3(new_n665), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(KEYINPUT46), .Z(new_n704));
  OAI21_X1  g503(.A(G36gat), .B1(new_n700), .B2(new_n452), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(G1329gat));
  OAI21_X1  g505(.A(G43gat), .B1(new_n700), .B2(new_n447), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT103), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n708), .A2(KEYINPUT47), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n441), .A2(G43gat), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n709), .B1(new_n680), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n708), .A2(KEYINPUT47), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n713), .B(KEYINPUT104), .Z(new_n714));
  XOR2_X1   g513(.A(new_n712), .B(new_n714), .Z(G1330gat));
  OAI21_X1  g514(.A(G50gat), .B1(new_n700), .B2(new_n379), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n680), .A2(new_n532), .A3(new_n454), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(KEYINPUT48), .B1(new_n717), .B2(KEYINPUT105), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1331gat));
  NAND4_X1  g519(.A1(new_n514), .A2(new_n581), .A3(new_n684), .A4(new_n658), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n721), .B1(new_n694), .B2(new_n698), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n661), .B(KEYINPUT106), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g524(.A1(new_n722), .A2(new_n665), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n727));
  XOR2_X1   g526(.A(KEYINPUT49), .B(G64gat), .Z(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n726), .B2(new_n728), .ZN(G1333gat));
  XNOR2_X1  g528(.A(new_n441), .B(KEYINPUT107), .ZN(new_n730));
  AOI21_X1  g529(.A(G71gat), .B1(new_n722), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(G71gat), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n447), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n731), .B1(new_n722), .B2(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g534(.A1(new_n722), .A2(new_n454), .ZN(new_n736));
  XNOR2_X1  g535(.A(KEYINPUT108), .B(G78gat), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1335gat));
  NAND2_X1  g537(.A1(new_n597), .A2(new_n599), .ZN(new_n739));
  INV_X1    g538(.A(new_n658), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n514), .A2(new_n580), .A3(new_n740), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n683), .B(new_n741), .C1(new_n699), .C2(KEYINPUT44), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n739), .B1(new_n742), .B2(new_n662), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n514), .A2(new_n580), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n699), .A2(KEYINPUT51), .A3(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(KEYINPUT51), .B1(new_n699), .B2(new_n744), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n661), .A2(new_n597), .A3(new_n599), .A4(new_n658), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n743), .B1(new_n748), .B2(new_n749), .ZN(G1336gat));
  OAI21_X1  g549(.A(G92gat), .B1(new_n742), .B2(new_n452), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n452), .A2(G92gat), .A3(new_n740), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n689), .A2(new_n691), .A3(new_n685), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT102), .B1(new_n458), .B2(new_n463), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n698), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n756), .A2(new_n633), .A3(new_n744), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT51), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n753), .B1(new_n759), .B2(new_n745), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n751), .B1(new_n760), .B2(KEYINPUT109), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n762));
  AOI211_X1 g561(.A(new_n762), .B(new_n753), .C1(new_n759), .C2(new_n745), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT52), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n760), .A2(KEYINPUT52), .ZN(new_n765));
  AOI21_X1  g564(.A(KEYINPUT110), .B1(new_n765), .B2(new_n751), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n752), .B1(new_n746), .B2(new_n747), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768));
  AND4_X1   g567(.A1(KEYINPUT110), .A2(new_n767), .A3(new_n751), .A4(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n764), .B1(new_n766), .B2(new_n769), .ZN(G1337gat));
  OAI21_X1  g569(.A(G99gat), .B1(new_n742), .B2(new_n447), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n459), .A2(new_n601), .A3(new_n658), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n771), .B1(new_n748), .B2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(G1338gat));
  INV_X1    g574(.A(KEYINPUT53), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n454), .A2(new_n602), .A3(new_n658), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT112), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n746), .B2(new_n747), .ZN(new_n779));
  OAI21_X1  g578(.A(KEYINPUT113), .B1(new_n742), .B2(new_n379), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(G106gat), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n742), .A2(KEYINPUT113), .A3(new_n379), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n776), .B(new_n779), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(G106gat), .B1(new_n742), .B2(new_n379), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n779), .A2(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n783), .B1(new_n776), .B2(new_n785), .ZN(G1339gat));
  NAND3_X1  g585(.A1(new_n637), .A2(new_n639), .A3(new_n647), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n642), .A2(KEYINPUT54), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g587(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n645), .B1(new_n656), .B2(new_n789), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n788), .A2(KEYINPUT55), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n788), .A2(new_n790), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n653), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n555), .A2(new_n569), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n576), .B1(new_n796), .B2(new_n554), .ZN(new_n797));
  AND4_X1   g596(.A1(new_n554), .A2(new_n555), .A3(new_n569), .A4(new_n576), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n792), .B(new_n795), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n550), .B1(new_n549), .B2(new_n551), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n566), .A2(new_n568), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n575), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n658), .A2(new_n579), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n633), .B1(new_n799), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n579), .A2(new_n802), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT55), .B1(new_n788), .B2(new_n790), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n791), .A2(new_n806), .A3(new_n653), .ZN(new_n807));
  AND3_X1   g606(.A1(new_n633), .A2(new_n805), .A3(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT115), .B1(new_n804), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT115), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n633), .A2(new_n807), .A3(new_n805), .ZN(new_n811));
  AOI22_X1  g610(.A1(new_n807), .A2(new_n580), .B1(new_n805), .B2(new_n658), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n810), .B(new_n811), .C1(new_n812), .C2(new_n633), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n809), .A2(new_n515), .A3(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n514), .A2(new_n581), .A3(new_n684), .A4(new_n740), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n815), .B1(new_n814), .B2(new_n816), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n662), .A2(new_n665), .A3(new_n441), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n819), .A2(new_n379), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(G113gat), .B1(new_n821), .B2(new_n581), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n814), .A2(new_n816), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT116), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n825));
  AND3_X1   g624(.A1(new_n824), .A2(new_n723), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(new_n690), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n580), .A2(new_n313), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n822), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  XOR2_X1   g629(.A(new_n830), .B(KEYINPUT117), .Z(G1340gat));
  NOR3_X1   g630(.A1(new_n821), .A2(new_n316), .A3(new_n740), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n826), .A2(new_n827), .A3(new_n658), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(new_n316), .B2(new_n833), .ZN(G1341gat));
  OAI21_X1  g633(.A(G127gat), .B1(new_n821), .B2(new_n515), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n515), .A2(G127gat), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n835), .B1(new_n828), .B2(new_n836), .ZN(G1342gat));
  OR2_X1    g636(.A1(new_n821), .A2(new_n684), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n684), .A2(G134gat), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n828), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT56), .ZN(new_n841));
  AOI22_X1  g640(.A1(new_n838), .A2(G134gat), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n840), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(new_n844), .A3(KEYINPUT56), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n844), .B1(new_n843), .B2(KEYINPUT56), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n842), .B1(new_n846), .B2(new_n847), .ZN(G1343gat));
  NOR2_X1   g647(.A1(new_n804), .A2(new_n808), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n816), .B1(new_n514), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n379), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n817), .A2(new_n818), .A3(new_n379), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(KEYINPUT57), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n447), .A2(new_n452), .A3(new_n661), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(KEYINPUT119), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n447), .A2(new_n858), .A3(new_n661), .A4(new_n452), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n855), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(G141gat), .B1(new_n862), .B2(new_n581), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n447), .A2(new_n454), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n665), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n581), .A2(G141gat), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n826), .A2(new_n865), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  NAND4_X1  g668(.A1(new_n824), .A2(new_n723), .A3(new_n825), .A4(new_n867), .ZN(new_n870));
  INV_X1    g669(.A(new_n868), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT120), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g672(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n863), .A2(new_n864), .A3(new_n873), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n873), .A2(new_n875), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n824), .A2(new_n454), .A3(new_n825), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n851), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n860), .B1(new_n879), .B2(new_n853), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n294), .B1(new_n880), .B2(new_n580), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT122), .B1(new_n877), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n870), .A2(new_n871), .ZN(new_n883));
  OAI21_X1  g682(.A(KEYINPUT58), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n876), .A2(new_n882), .A3(new_n884), .ZN(G1344gat));
  NAND3_X1  g684(.A1(new_n855), .A2(new_n658), .A3(new_n861), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n301), .A2(KEYINPUT59), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n857), .A2(new_n658), .A3(new_n859), .ZN(new_n888));
  INV_X1    g687(.A(new_n852), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n817), .A2(new_n818), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT57), .B1(new_n850), .B2(new_n454), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(G148gat), .ZN(new_n893));
  XOR2_X1   g692(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n894));
  AOI22_X1  g693(.A1(new_n886), .A2(new_n887), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n658), .A2(new_n301), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n870), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT124), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT124), .ZN(new_n899));
  INV_X1    g698(.A(new_n897), .ZN(new_n900));
  INV_X1    g699(.A(new_n887), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n901), .B1(new_n880), .B2(new_n658), .ZN(new_n902));
  INV_X1    g701(.A(new_n894), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n903), .B1(new_n892), .B2(G148gat), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n899), .B(new_n900), .C1(new_n902), .C2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n898), .A2(new_n905), .ZN(G1345gat));
  OAI21_X1  g705(.A(G155gat), .B1(new_n862), .B2(new_n515), .ZN(new_n907));
  INV_X1    g706(.A(new_n870), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n290), .A3(new_n514), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1346gat));
  AOI21_X1  g709(.A(G162gat), .B1(new_n908), .B2(new_n633), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n684), .A2(new_n291), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(new_n880), .B2(new_n912), .ZN(G1347gat));
  NOR2_X1   g712(.A1(new_n723), .A2(new_n452), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n819), .A2(new_n914), .A3(new_n379), .A4(new_n730), .ZN(new_n915));
  OAI21_X1  g714(.A(G169gat), .B1(new_n915), .B2(new_n581), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n817), .A2(new_n818), .A3(new_n661), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n457), .A2(new_n452), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n580), .A2(new_n233), .A3(new_n234), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(G1348gat));
  OAI21_X1  g720(.A(G176gat), .B1(new_n915), .B2(new_n740), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n658), .A2(new_n227), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n919), .B2(new_n923), .ZN(G1349gat));
  OAI21_X1  g723(.A(new_n222), .B1(new_n915), .B2(new_n515), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n515), .A2(new_n265), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n919), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT60), .ZN(G1350gat));
  OR2_X1    g727(.A1(new_n915), .A2(new_n684), .ZN(new_n929));
  XNOR2_X1  g728(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n929), .A2(G190gat), .A3(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n930), .B1(new_n929), .B2(G190gat), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n633), .A2(new_n217), .ZN(new_n934));
  OAI22_X1  g733(.A1(new_n932), .A2(new_n933), .B1(new_n919), .B2(new_n934), .ZN(G1351gat));
  NOR2_X1   g734(.A1(new_n866), .A2(new_n452), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n917), .A2(new_n936), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n937), .A2(G197gat), .A3(new_n581), .ZN(new_n938));
  XOR2_X1   g737(.A(new_n938), .B(KEYINPUT126), .Z(new_n939));
  NOR2_X1   g738(.A1(new_n890), .A2(new_n891), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n914), .A2(new_n447), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n580), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(G197gat), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n939), .A2(new_n944), .ZN(G1352gat));
  INV_X1    g744(.A(new_n941), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n946), .B(new_n658), .C1(new_n891), .C2(new_n890), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(G204gat), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n740), .A2(G204gat), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(KEYINPUT62), .B1(new_n937), .B2(new_n950), .ZN(new_n951));
  OR3_X1    g750(.A1(new_n937), .A2(KEYINPUT62), .A3(new_n950), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n948), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT127), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n948), .A2(new_n955), .A3(new_n951), .A4(new_n952), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1353gat));
  INV_X1    g756(.A(new_n937), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n958), .A2(new_n208), .A3(new_n514), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n514), .ZN(new_n960));
  AND3_X1   g759(.A1(new_n960), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n961));
  AOI21_X1  g760(.A(KEYINPUT63), .B1(new_n960), .B2(G211gat), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n959), .B1(new_n961), .B2(new_n962), .ZN(G1354gat));
  NAND3_X1  g762(.A1(new_n958), .A2(new_n209), .A3(new_n633), .ZN(new_n964));
  NOR3_X1   g763(.A1(new_n940), .A2(new_n684), .A3(new_n941), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(new_n209), .ZN(G1355gat));
endmodule


