

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730;

  NOR2_X1 U368 ( .A1(n627), .A2(n727), .ZN(n585) );
  INV_X1 U369 ( .A(G143), .ZN(n451) );
  OR2_X1 U370 ( .A1(n685), .A2(G902), .ZN(n417) );
  XNOR2_X2 U371 ( .A(n428), .B(n542), .ZN(n570) );
  XNOR2_X2 U372 ( .A(n417), .B(n416), .ZN(n547) );
  XOR2_X1 U373 ( .A(KEYINPUT68), .B(G101), .Z(n489) );
  XOR2_X2 U374 ( .A(G146), .B(G125), .Z(n471) );
  AND2_X2 U375 ( .A1(n604), .A2(n603), .ZN(n699) );
  XNOR2_X1 U376 ( .A(n560), .B(KEYINPUT48), .ZN(n405) );
  AND2_X1 U377 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U378 ( .A1(n420), .A2(n555), .ZN(n550) );
  NOR2_X2 U379 ( .A1(n523), .A2(n600), .ZN(n429) );
  XNOR2_X1 U380 ( .A(n463), .B(n462), .ZN(n386) );
  NAND2_X1 U381 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X2 U382 ( .A(KEYINPUT0), .B(n571), .ZN(n578) );
  XNOR2_X1 U383 ( .A(n386), .B(n362), .ZN(n718) );
  XNOR2_X1 U384 ( .A(n486), .B(n363), .ZN(n362) );
  XNOR2_X1 U385 ( .A(n364), .B(G137), .ZN(n363) );
  INV_X1 U386 ( .A(KEYINPUT4), .ZN(n364) );
  XNOR2_X1 U387 ( .A(n718), .B(n487), .ZN(n385) );
  INV_X1 U388 ( .A(G146), .ZN(n487) );
  INV_X1 U389 ( .A(KEYINPUT6), .ZN(n442) );
  NAND2_X1 U390 ( .A1(n346), .A2(n370), .ZN(n369) );
  INV_X1 U391 ( .A(n631), .ZN(n370) );
  NOR2_X1 U392 ( .A1(n633), .A2(n545), .ZN(n546) );
  NOR2_X1 U393 ( .A1(G237), .A2(G902), .ZN(n494) );
  XNOR2_X1 U394 ( .A(n448), .B(n447), .ZN(n490) );
  XNOR2_X1 U395 ( .A(n446), .B(G113), .ZN(n447) );
  INV_X1 U396 ( .A(G119), .ZN(n446) );
  INV_X1 U397 ( .A(KEYINPUT1), .ZN(n415) );
  XNOR2_X1 U398 ( .A(n472), .B(n473), .ZN(n717) );
  XOR2_X1 U399 ( .A(KEYINPUT71), .B(KEYINPUT10), .Z(n473) );
  XNOR2_X1 U400 ( .A(n385), .B(n501), .ZN(n685) );
  XOR2_X1 U401 ( .A(KEYINPUT83), .B(G140), .Z(n498) );
  NAND2_X1 U402 ( .A1(n590), .A2(n351), .ZN(n413) );
  OR2_X1 U403 ( .A1(n400), .A2(n441), .ZN(n381) );
  INV_X1 U404 ( .A(KEYINPUT50), .ZN(n380) );
  NOR2_X1 U405 ( .A1(n643), .A2(n404), .ZN(n403) );
  INV_X1 U406 ( .A(n644), .ZN(n404) );
  NOR2_X1 U407 ( .A1(n369), .A2(n367), .ZN(n558) );
  XNOR2_X1 U408 ( .A(G113), .B(G122), .ZN(n476) );
  OR2_X1 U409 ( .A1(n698), .A2(G902), .ZN(n411) );
  XNOR2_X1 U410 ( .A(n444), .B(n350), .ZN(n443) );
  XNOR2_X1 U411 ( .A(n490), .B(n492), .ZN(n444) );
  AND2_X1 U412 ( .A1(n405), .A2(n403), .ZN(n437) );
  XOR2_X1 U413 ( .A(KEYINPUT82), .B(G110), .Z(n507) );
  XNOR2_X1 U414 ( .A(G128), .B(G137), .ZN(n506) );
  XNOR2_X1 U415 ( .A(G119), .B(KEYINPUT24), .ZN(n504) );
  XOR2_X1 U416 ( .A(KEYINPUT95), .B(KEYINPUT23), .Z(n505) );
  XNOR2_X1 U417 ( .A(n467), .B(KEYINPUT102), .ZN(n423) );
  XNOR2_X1 U418 ( .A(G116), .B(G107), .ZN(n467) );
  INV_X1 U419 ( .A(G134), .ZN(n462) );
  XNOR2_X1 U420 ( .A(n469), .B(n468), .ZN(n412) );
  XNOR2_X1 U421 ( .A(KEYINPUT87), .B(KEYINPUT8), .ZN(n468) );
  XNOR2_X1 U422 ( .A(n529), .B(KEYINPUT39), .ZN(n532) );
  XOR2_X1 U423 ( .A(n400), .B(KEYINPUT92), .Z(n573) );
  NAND2_X1 U424 ( .A1(n398), .A2(n354), .ZN(n561) );
  AND2_X1 U425 ( .A1(n552), .A2(n351), .ZN(n398) );
  NOR2_X1 U426 ( .A1(n587), .A2(n581), .ZN(n392) );
  XNOR2_X1 U427 ( .A(n410), .B(n408), .ZN(n407) );
  INV_X1 U428 ( .A(KEYINPUT28), .ZN(n408) );
  AND2_X1 U429 ( .A1(n552), .A2(n649), .ZN(n410) );
  INV_X1 U430 ( .A(G469), .ZN(n416) );
  INV_X1 U431 ( .A(KEYINPUT22), .ZN(n434) );
  BUF_X1 U432 ( .A(n579), .Z(n400) );
  XNOR2_X1 U433 ( .A(n481), .B(n348), .ZN(n482) );
  XNOR2_X1 U434 ( .A(n461), .B(n460), .ZN(n606) );
  AND2_X1 U435 ( .A1(n376), .A2(n375), .ZN(n680) );
  INV_X1 U436 ( .A(n676), .ZN(n375) );
  NAND2_X1 U437 ( .A1(n418), .A2(n419), .ZN(n368) );
  INV_X1 U438 ( .A(n573), .ZN(n418) );
  XNOR2_X1 U439 ( .A(n371), .B(KEYINPUT36), .ZN(n419) );
  NOR2_X1 U440 ( .A1(n561), .A2(n563), .ZN(n371) );
  XNOR2_X1 U441 ( .A(n368), .B(n553), .ZN(n367) );
  XNOR2_X1 U442 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n454) );
  XOR2_X1 U443 ( .A(KEYINPUT18), .B(KEYINPUT93), .Z(n455) );
  XNOR2_X1 U444 ( .A(n381), .B(n380), .ZN(n653) );
  XOR2_X1 U445 ( .A(KEYINPUT5), .B(KEYINPUT97), .Z(n488) );
  INV_X1 U446 ( .A(KEYINPUT44), .ZN(n361) );
  XNOR2_X1 U447 ( .A(n705), .B(n430), .ZN(n500) );
  XNOR2_X1 U448 ( .A(n489), .B(n431), .ZN(n430) );
  INV_X1 U449 ( .A(KEYINPUT74), .ZN(n431) );
  NAND2_X1 U450 ( .A1(G234), .A2(G237), .ZN(n512) );
  XOR2_X1 U451 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n513) );
  XNOR2_X1 U452 ( .A(n394), .B(KEYINPUT77), .ZN(n590) );
  NOR2_X1 U453 ( .A1(n646), .A2(n535), .ZN(n536) );
  XNOR2_X1 U454 ( .A(n526), .B(n525), .ZN(n527) );
  INV_X1 U455 ( .A(KEYINPUT85), .ZN(n525) );
  XNOR2_X1 U456 ( .A(G953), .B(KEYINPUT64), .ZN(n516) );
  XNOR2_X1 U457 ( .A(n449), .B(n432), .ZN(n705) );
  XNOR2_X1 U458 ( .A(G104), .B(G107), .ZN(n449) );
  XNOR2_X1 U459 ( .A(n433), .B(G110), .ZN(n432) );
  INV_X1 U460 ( .A(KEYINPUT79), .ZN(n433) );
  XNOR2_X1 U461 ( .A(KEYINPUT16), .B(G122), .ZN(n395) );
  AND2_X1 U462 ( .A1(n405), .A2(n345), .ZN(n439) );
  NOR2_X1 U463 ( .A1(G237), .A2(G953), .ZN(n480) );
  XNOR2_X1 U464 ( .A(n365), .B(KEYINPUT72), .ZN(n486) );
  INV_X1 U465 ( .A(G131), .ZN(n365) );
  XNOR2_X1 U466 ( .A(G143), .B(G104), .ZN(n474) );
  AND2_X1 U467 ( .A1(n521), .A2(n520), .ZN(n556) );
  NOR2_X1 U468 ( .A1(n586), .A2(n519), .ZN(n520) );
  XNOR2_X1 U469 ( .A(n485), .B(n399), .ZN(n554) );
  XNOR2_X1 U470 ( .A(n484), .B(G475), .ZN(n399) );
  XNOR2_X1 U471 ( .A(n493), .B(G472), .ZN(n588) );
  INV_X1 U472 ( .A(n721), .ZN(n366) );
  XNOR2_X1 U473 ( .A(n373), .B(n372), .ZN(n698) );
  XNOR2_X1 U474 ( .A(n445), .B(n347), .ZN(n372) );
  XNOR2_X1 U475 ( .A(n717), .B(n374), .ZN(n373) );
  XNOR2_X1 U476 ( .A(n424), .B(n421), .ZN(n696) );
  XNOR2_X1 U477 ( .A(n466), .B(n423), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n533), .B(KEYINPUT40), .ZN(n730) );
  NAND2_X1 U479 ( .A1(n532), .A2(n544), .ZN(n533) );
  NAND2_X1 U480 ( .A1(n388), .A2(n387), .ZN(n583) );
  NAND2_X1 U481 ( .A1(n393), .A2(n392), .ZN(n387) );
  AND2_X1 U482 ( .A1(n389), .A2(n390), .ZN(n388) );
  XNOR2_X1 U483 ( .A(n427), .B(n425), .ZN(n727) );
  XNOR2_X1 U484 ( .A(n426), .B(KEYINPUT32), .ZN(n425) );
  INV_X1 U485 ( .A(KEYINPUT66), .ZN(n426) );
  OR2_X1 U486 ( .A1(n407), .A2(n406), .ZN(n633) );
  NAND2_X1 U487 ( .A1(n570), .A2(n409), .ZN(n406) );
  XNOR2_X1 U488 ( .A(n550), .B(n549), .ZN(n635) );
  INV_X1 U489 ( .A(n400), .ZN(n651) );
  AND2_X1 U490 ( .A1(n614), .A2(n613), .ZN(n617) );
  NOR2_X1 U491 ( .A1(n694), .A2(n703), .ZN(n396) );
  XNOR2_X1 U492 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U493 ( .A(n689), .B(n688), .ZN(n402) );
  NOR2_X1 U494 ( .A1(n607), .A2(n703), .ZN(n397) );
  XNOR2_X1 U495 ( .A(n382), .B(KEYINPUT121), .ZN(n684) );
  INV_X1 U496 ( .A(n368), .ZN(n640) );
  AND2_X1 U497 ( .A1(n403), .A2(n600), .ZN(n345) );
  XNOR2_X1 U498 ( .A(n546), .B(KEYINPUT47), .ZN(n346) );
  XOR2_X1 U499 ( .A(n505), .B(n504), .Z(n347) );
  AND2_X1 U500 ( .A1(n491), .A2(G214), .ZN(n348) );
  AND2_X1 U501 ( .A1(n438), .A2(n437), .ZN(n349) );
  INV_X1 U502 ( .A(n547), .ZN(n409) );
  XOR2_X1 U503 ( .A(n489), .B(n488), .Z(n350) );
  INV_X1 U504 ( .A(n652), .ZN(n441) );
  XOR2_X1 U505 ( .A(n588), .B(n442), .Z(n351) );
  AND2_X1 U506 ( .A1(n599), .A2(n618), .ZN(n352) );
  XNOR2_X1 U507 ( .A(KEYINPUT119), .B(n675), .ZN(n353) );
  AND2_X1 U508 ( .A1(n551), .A2(n663), .ZN(n354) );
  XNOR2_X1 U509 ( .A(KEYINPUT34), .B(KEYINPUT84), .ZN(n581) );
  XNOR2_X1 U510 ( .A(G902), .B(KEYINPUT15), .ZN(n522) );
  XNOR2_X1 U511 ( .A(n490), .B(n395), .ZN(n704) );
  NOR2_X1 U512 ( .A1(n720), .A2(G952), .ZN(n703) );
  INV_X1 U513 ( .A(G953), .ZN(n683) );
  AND2_X2 U514 ( .A1(n355), .A2(n352), .ZN(n358) );
  NAND2_X1 U515 ( .A1(n356), .A2(KEYINPUT44), .ZN(n355) );
  NAND2_X1 U516 ( .A1(n584), .A2(n585), .ZN(n356) );
  NAND2_X2 U517 ( .A1(n358), .A2(n357), .ZN(n414) );
  NAND2_X1 U518 ( .A1(n360), .A2(n359), .ZN(n357) );
  AND2_X1 U519 ( .A1(n585), .A2(n361), .ZN(n359) );
  XNOR2_X1 U520 ( .A(n726), .B(KEYINPUT69), .ZN(n360) );
  XNOR2_X2 U521 ( .A(n451), .B(G128), .ZN(n463) );
  XNOR2_X1 U522 ( .A(n547), .B(n415), .ZN(n579) );
  NAND2_X1 U523 ( .A1(n595), .A2(n574), .ZN(n427) );
  XNOR2_X1 U524 ( .A(n437), .B(n366), .ZN(n719) );
  NAND2_X1 U525 ( .A1(n412), .A2(G221), .ZN(n374) );
  XNOR2_X1 U526 ( .A(n377), .B(KEYINPUT52), .ZN(n376) );
  NAND2_X1 U527 ( .A1(n378), .A2(n353), .ZN(n377) );
  XNOR2_X1 U528 ( .A(n661), .B(n379), .ZN(n378) );
  INV_X1 U529 ( .A(KEYINPUT115), .ZN(n379) );
  NAND2_X1 U530 ( .A1(n384), .A2(n383), .ZN(n382) );
  XNOR2_X1 U531 ( .A(n681), .B(KEYINPUT120), .ZN(n383) );
  NOR2_X1 U532 ( .A1(n682), .A2(G953), .ZN(n384) );
  XNOR2_X1 U533 ( .A(n385), .B(n443), .ZN(n610) );
  XNOR2_X1 U534 ( .A(n386), .B(n422), .ZN(n421) );
  NAND2_X1 U535 ( .A1(n678), .A2(n581), .ZN(n389) );
  AND2_X1 U536 ( .A1(n391), .A2(n582), .ZN(n390) );
  NAND2_X1 U537 ( .A1(n587), .A2(n581), .ZN(n391) );
  INV_X1 U538 ( .A(n678), .ZN(n393) );
  XNOR2_X2 U539 ( .A(n413), .B(n580), .ZN(n678) );
  XNOR2_X1 U540 ( .A(n605), .B(n606), .ZN(n607) );
  NAND2_X1 U541 ( .A1(n579), .A2(n441), .ZN(n394) );
  XNOR2_X1 U542 ( .A(n396), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U543 ( .A(n397), .B(n609), .ZN(G51) );
  XNOR2_X1 U544 ( .A(n483), .B(n482), .ZN(n691) );
  INV_X1 U545 ( .A(n438), .ZN(n711) );
  NAND2_X1 U546 ( .A1(n438), .A2(n439), .ZN(n440) );
  XNOR2_X2 U547 ( .A(n414), .B(KEYINPUT45), .ZN(n438) );
  NAND2_X1 U548 ( .A1(n402), .A2(n613), .ZN(n401) );
  XNOR2_X1 U549 ( .A(n401), .B(KEYINPUT123), .ZN(G54) );
  NOR2_X1 U550 ( .A1(n407), .A2(n547), .ZN(n543) );
  XNOR2_X2 U551 ( .A(n411), .B(n511), .ZN(n646) );
  NAND2_X1 U552 ( .A1(n412), .A2(G217), .ZN(n424) );
  INV_X1 U553 ( .A(n555), .ZN(n531) );
  INV_X1 U554 ( .A(n550), .ZN(n544) );
  INV_X1 U555 ( .A(n554), .ZN(n420) );
  XNOR2_X1 U556 ( .A(n440), .B(KEYINPUT88), .ZN(n602) );
  NAND2_X1 U557 ( .A1(n548), .A2(n663), .ZN(n428) );
  XNOR2_X2 U558 ( .A(n429), .B(n527), .ZN(n548) );
  INV_X1 U559 ( .A(n578), .ZN(n591) );
  XNOR2_X1 U560 ( .A(n435), .B(n434), .ZN(n575) );
  NOR2_X1 U561 ( .A1(n578), .A2(n436), .ZN(n435) );
  NAND2_X1 U562 ( .A1(n572), .A2(n645), .ZN(n436) );
  XOR2_X1 U563 ( .A(n507), .B(n506), .Z(n445) );
  INV_X1 U564 ( .A(KEYINPUT90), .ZN(n553) );
  INV_X1 U565 ( .A(n534), .ZN(n519) );
  INV_X1 U566 ( .A(KEYINPUT105), .ZN(n549) );
  INV_X1 U567 ( .A(KEYINPUT106), .ZN(n615) );
  XNOR2_X1 U568 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U569 ( .A(n615), .B(KEYINPUT63), .ZN(n616) );
  XNOR2_X1 U570 ( .A(n617), .B(n616), .ZN(G57) );
  INV_X1 U571 ( .A(n516), .ZN(n720) );
  XOR2_X1 U572 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n461) );
  XNOR2_X1 U573 ( .A(KEYINPUT3), .B(G116), .ZN(n448) );
  INV_X1 U574 ( .A(n500), .ZN(n450) );
  XNOR2_X1 U575 ( .A(n704), .B(n450), .ZN(n459) );
  XOR2_X1 U576 ( .A(n463), .B(n471), .Z(n453) );
  NAND2_X1 U577 ( .A1(G224), .A2(n720), .ZN(n452) );
  XNOR2_X1 U578 ( .A(n453), .B(n452), .ZN(n457) );
  XNOR2_X1 U579 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U580 ( .A(n457), .B(n456), .Z(n458) );
  XNOR2_X1 U581 ( .A(n459), .B(n458), .ZN(n523) );
  XNOR2_X1 U582 ( .A(n523), .B(KEYINPUT86), .ZN(n460) );
  XOR2_X1 U583 ( .A(KEYINPUT9), .B(KEYINPUT103), .Z(n465) );
  XNOR2_X1 U584 ( .A(G122), .B(KEYINPUT7), .ZN(n464) );
  XNOR2_X1 U585 ( .A(n465), .B(n464), .ZN(n466) );
  NAND2_X1 U586 ( .A1(n720), .A2(G234), .ZN(n469) );
  NOR2_X1 U587 ( .A1(G902), .A2(n696), .ZN(n470) );
  XNOR2_X1 U588 ( .A(G478), .B(n470), .ZN(n555) );
  XNOR2_X1 U589 ( .A(n471), .B(G140), .ZN(n472) );
  XNOR2_X1 U590 ( .A(n486), .B(n717), .ZN(n483) );
  XOR2_X1 U591 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n475) );
  XNOR2_X1 U592 ( .A(n475), .B(n474), .ZN(n479) );
  XOR2_X1 U593 ( .A(KEYINPUT11), .B(KEYINPUT99), .Z(n477) );
  XNOR2_X1 U594 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U595 ( .A(n479), .B(n478), .Z(n481) );
  XNOR2_X1 U596 ( .A(n480), .B(KEYINPUT80), .ZN(n491) );
  NOR2_X1 U597 ( .A1(G902), .A2(n691), .ZN(n485) );
  XNOR2_X1 U598 ( .A(KEYINPUT13), .B(KEYINPUT101), .ZN(n484) );
  NAND2_X1 U599 ( .A1(n531), .A2(n554), .ZN(n637) );
  INV_X1 U600 ( .A(KEYINPUT30), .ZN(n496) );
  NAND2_X1 U601 ( .A1(n491), .A2(G210), .ZN(n492) );
  NOR2_X1 U602 ( .A1(n610), .A2(G902), .ZN(n493) );
  INV_X1 U603 ( .A(n588), .ZN(n649) );
  XOR2_X1 U604 ( .A(KEYINPUT78), .B(n494), .Z(n524) );
  NAND2_X1 U605 ( .A1(n524), .A2(G214), .ZN(n663) );
  NAND2_X1 U606 ( .A1(n649), .A2(n663), .ZN(n495) );
  XNOR2_X1 U607 ( .A(n496), .B(n495), .ZN(n521) );
  NAND2_X1 U608 ( .A1(G227), .A2(n720), .ZN(n497) );
  XNOR2_X1 U609 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U610 ( .A(n500), .B(n499), .ZN(n501) );
  NAND2_X1 U611 ( .A1(n522), .A2(G234), .ZN(n502) );
  XNOR2_X1 U612 ( .A(n502), .B(KEYINPUT20), .ZN(n508) );
  NAND2_X1 U613 ( .A1(G221), .A2(n508), .ZN(n503) );
  XOR2_X1 U614 ( .A(KEYINPUT21), .B(n503), .Z(n645) );
  XOR2_X1 U615 ( .A(KEYINPUT25), .B(KEYINPUT96), .Z(n510) );
  NAND2_X1 U616 ( .A1(G217), .A2(n508), .ZN(n509) );
  XNOR2_X1 U617 ( .A(n510), .B(n509), .ZN(n511) );
  NAND2_X1 U618 ( .A1(n645), .A2(n646), .ZN(n652) );
  OR2_X1 U619 ( .A1(n547), .A2(n652), .ZN(n586) );
  XNOR2_X1 U620 ( .A(n513), .B(n512), .ZN(n515) );
  NAND2_X1 U621 ( .A1(G952), .A2(n515), .ZN(n676) );
  NOR2_X1 U622 ( .A1(G953), .A2(n676), .ZN(n514) );
  XOR2_X1 U623 ( .A(KEYINPUT94), .B(n514), .Z(n568) );
  NAND2_X1 U624 ( .A1(G902), .A2(n515), .ZN(n565) );
  NOR2_X1 U625 ( .A1(G900), .A2(n565), .ZN(n517) );
  NAND2_X1 U626 ( .A1(n517), .A2(n516), .ZN(n518) );
  NAND2_X1 U627 ( .A1(n568), .A2(n518), .ZN(n534) );
  XNOR2_X1 U628 ( .A(KEYINPUT38), .B(KEYINPUT76), .ZN(n528) );
  INV_X1 U629 ( .A(n522), .ZN(n600) );
  NAND2_X1 U630 ( .A1(n524), .A2(G210), .ZN(n526) );
  XOR2_X1 U631 ( .A(n528), .B(n548), .Z(n662) );
  NAND2_X1 U632 ( .A1(n556), .A2(n662), .ZN(n529) );
  INV_X1 U633 ( .A(n532), .ZN(n530) );
  NOR2_X1 U634 ( .A1(n637), .A2(n530), .ZN(n643) );
  NAND2_X1 U635 ( .A1(n645), .A2(n534), .ZN(n535) );
  XOR2_X1 U636 ( .A(n536), .B(KEYINPUT73), .Z(n552) );
  NAND2_X1 U637 ( .A1(n555), .A2(n554), .ZN(n666) );
  NAND2_X1 U638 ( .A1(n663), .A2(n662), .ZN(n669) );
  NOR2_X1 U639 ( .A1(n666), .A2(n669), .ZN(n537) );
  XNOR2_X1 U640 ( .A(KEYINPUT41), .B(n537), .ZN(n677) );
  INV_X1 U641 ( .A(n677), .ZN(n659) );
  NAND2_X1 U642 ( .A1(n543), .A2(n659), .ZN(n538) );
  XNOR2_X1 U643 ( .A(KEYINPUT42), .B(n538), .ZN(n728) );
  NAND2_X1 U644 ( .A1(n730), .A2(n728), .ZN(n540) );
  XNOR2_X1 U645 ( .A(KEYINPUT65), .B(KEYINPUT46), .ZN(n539) );
  XNOR2_X1 U646 ( .A(n540), .B(n539), .ZN(n559) );
  XNOR2_X1 U647 ( .A(KEYINPUT19), .B(KEYINPUT67), .ZN(n541) );
  XNOR2_X1 U648 ( .A(n541), .B(KEYINPUT81), .ZN(n542) );
  NAND2_X1 U649 ( .A1(n550), .A2(n637), .ZN(n668) );
  NAND2_X1 U650 ( .A1(KEYINPUT70), .A2(n668), .ZN(n545) );
  INV_X1 U651 ( .A(n548), .ZN(n563) );
  INV_X1 U652 ( .A(n635), .ZN(n551) );
  NOR2_X1 U653 ( .A1(n555), .A2(n554), .ZN(n582) );
  NAND2_X1 U654 ( .A1(n556), .A2(n582), .ZN(n557) );
  NOR2_X1 U655 ( .A1(n563), .A2(n557), .ZN(n631) );
  OR2_X1 U656 ( .A1(n400), .A2(n561), .ZN(n562) );
  XNOR2_X1 U657 ( .A(n562), .B(KEYINPUT43), .ZN(n564) );
  NAND2_X1 U658 ( .A1(n564), .A2(n563), .ZN(n644) );
  INV_X1 U659 ( .A(n565), .ZN(n566) );
  NOR2_X1 U660 ( .A1(G898), .A2(n683), .ZN(n707) );
  NAND2_X1 U661 ( .A1(n566), .A2(n707), .ZN(n567) );
  NAND2_X1 U662 ( .A1(n568), .A2(n567), .ZN(n569) );
  INV_X1 U663 ( .A(n666), .ZN(n572) );
  NOR2_X2 U664 ( .A1(n575), .A2(n351), .ZN(n595) );
  NOR2_X1 U665 ( .A1(n573), .A2(n646), .ZN(n574) );
  NOR2_X1 U666 ( .A1(n649), .A2(n575), .ZN(n576) );
  INV_X1 U667 ( .A(n646), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n576), .A2(n597), .ZN(n577) );
  NOR2_X1 U669 ( .A1(n400), .A2(n577), .ZN(n627) );
  BUF_X1 U670 ( .A(n578), .Z(n587) );
  XOR2_X1 U671 ( .A(KEYINPUT104), .B(KEYINPUT33), .Z(n580) );
  XNOR2_X2 U672 ( .A(n583), .B(KEYINPUT35), .ZN(n726) );
  NOR2_X1 U673 ( .A1(n726), .A2(KEYINPUT69), .ZN(n584) );
  NOR2_X1 U674 ( .A1(n587), .A2(n586), .ZN(n589) );
  NAND2_X1 U675 ( .A1(n589), .A2(n588), .ZN(n622) );
  XOR2_X1 U676 ( .A(KEYINPUT98), .B(KEYINPUT31), .Z(n593) );
  AND2_X1 U677 ( .A1(n590), .A2(n649), .ZN(n657) );
  NAND2_X1 U678 ( .A1(n657), .A2(n591), .ZN(n592) );
  XNOR2_X1 U679 ( .A(n593), .B(n592), .ZN(n638) );
  NAND2_X1 U680 ( .A1(n622), .A2(n638), .ZN(n594) );
  NAND2_X1 U681 ( .A1(n594), .A2(n668), .ZN(n599) );
  XNOR2_X1 U682 ( .A(KEYINPUT91), .B(n595), .ZN(n596) );
  NOR2_X1 U683 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U684 ( .A1(n651), .A2(n598), .ZN(n618) );
  NAND2_X1 U685 ( .A1(KEYINPUT2), .A2(n600), .ZN(n601) );
  NAND2_X1 U686 ( .A1(n602), .A2(n601), .ZN(n604) );
  NAND2_X1 U687 ( .A1(KEYINPUT2), .A2(n349), .ZN(n603) );
  NAND2_X1 U688 ( .A1(n699), .A2(G210), .ZN(n605) );
  INV_X1 U689 ( .A(KEYINPUT89), .ZN(n608) );
  XNOR2_X1 U690 ( .A(n608), .B(KEYINPUT56), .ZN(n609) );
  NAND2_X1 U691 ( .A1(n699), .A2(G472), .ZN(n612) );
  XOR2_X1 U692 ( .A(n610), .B(KEYINPUT62), .Z(n611) );
  XNOR2_X1 U693 ( .A(n612), .B(n611), .ZN(n614) );
  INV_X1 U694 ( .A(n703), .ZN(n613) );
  XNOR2_X1 U695 ( .A(G101), .B(n618), .ZN(G3) );
  NOR2_X1 U696 ( .A1(n635), .A2(n622), .ZN(n620) );
  XNOR2_X1 U697 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n619) );
  XNOR2_X1 U698 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U699 ( .A(G104), .B(n621), .ZN(G6) );
  NOR2_X1 U700 ( .A1(n622), .A2(n637), .ZN(n626) );
  XOR2_X1 U701 ( .A(KEYINPUT26), .B(KEYINPUT109), .Z(n624) );
  XNOR2_X1 U702 ( .A(G107), .B(KEYINPUT27), .ZN(n623) );
  XNOR2_X1 U703 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U704 ( .A(n626), .B(n625), .ZN(G9) );
  XOR2_X1 U705 ( .A(G110), .B(n627), .Z(G12) );
  NOR2_X1 U706 ( .A1(n637), .A2(n633), .ZN(n629) );
  XNOR2_X1 U707 ( .A(KEYINPUT110), .B(KEYINPUT29), .ZN(n628) );
  XNOR2_X1 U708 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U709 ( .A(G128), .B(n630), .ZN(G30) );
  XNOR2_X1 U710 ( .A(G143), .B(n631), .ZN(n632) );
  XNOR2_X1 U711 ( .A(n632), .B(KEYINPUT111), .ZN(G45) );
  NOR2_X1 U712 ( .A1(n635), .A2(n633), .ZN(n634) );
  XOR2_X1 U713 ( .A(G146), .B(n634), .Z(G48) );
  NOR2_X1 U714 ( .A1(n638), .A2(n635), .ZN(n636) );
  XOR2_X1 U715 ( .A(G113), .B(n636), .Z(G15) );
  NOR2_X1 U716 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U717 ( .A(G116), .B(n639), .Z(G18) );
  XNOR2_X1 U718 ( .A(n640), .B(KEYINPUT37), .ZN(n641) );
  XNOR2_X1 U719 ( .A(n641), .B(KEYINPUT112), .ZN(n642) );
  XNOR2_X1 U720 ( .A(G125), .B(n642), .ZN(G27) );
  XOR2_X1 U721 ( .A(G134), .B(n643), .Z(G36) );
  XNOR2_X1 U722 ( .A(G140), .B(n644), .ZN(G42) );
  NOR2_X1 U723 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U724 ( .A(KEYINPUT49), .B(n647), .Z(n648) );
  NOR2_X1 U725 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U726 ( .A(KEYINPUT113), .B(n650), .ZN(n654) );
  NOR2_X1 U727 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U728 ( .A(n655), .B(KEYINPUT114), .ZN(n656) );
  NOR2_X1 U729 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U730 ( .A(KEYINPUT51), .B(n658), .ZN(n660) );
  NAND2_X1 U731 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U733 ( .A(n664), .B(KEYINPUT116), .ZN(n665) );
  NOR2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U735 ( .A(KEYINPUT117), .B(n667), .Z(n673) );
  INV_X1 U736 ( .A(n668), .ZN(n670) );
  NOR2_X1 U737 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U738 ( .A(KEYINPUT118), .B(n671), .ZN(n672) );
  NOR2_X1 U739 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U740 ( .A1(n678), .A2(n674), .ZN(n675) );
  NOR2_X1 U741 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U742 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U743 ( .A(KEYINPUT2), .B(n349), .Z(n682) );
  XNOR2_X1 U744 ( .A(KEYINPUT53), .B(n684), .ZN(G75) );
  NAND2_X1 U745 ( .A1(n699), .A2(G469), .ZN(n689) );
  XNOR2_X1 U746 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n687) );
  XNOR2_X1 U747 ( .A(n685), .B(KEYINPUT57), .ZN(n686) );
  XNOR2_X1 U748 ( .A(n687), .B(n686), .ZN(n688) );
  NAND2_X1 U749 ( .A1(n699), .A2(G475), .ZN(n693) );
  XOR2_X1 U750 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n690) );
  NAND2_X1 U751 ( .A1(G478), .A2(n699), .ZN(n695) );
  XNOR2_X1 U752 ( .A(n696), .B(n695), .ZN(n697) );
  NOR2_X1 U753 ( .A1(n703), .A2(n697), .ZN(G63) );
  XOR2_X1 U754 ( .A(n698), .B(KEYINPUT125), .Z(n701) );
  NAND2_X1 U755 ( .A1(n699), .A2(G217), .ZN(n700) );
  XNOR2_X1 U756 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U757 ( .A1(n703), .A2(n702), .ZN(G66) );
  XOR2_X1 U758 ( .A(n705), .B(G101), .Z(n706) );
  XNOR2_X1 U759 ( .A(n704), .B(n706), .ZN(n708) );
  NOR2_X1 U760 ( .A1(n708), .A2(n707), .ZN(n715) );
  NAND2_X1 U761 ( .A1(G953), .A2(G224), .ZN(n709) );
  XNOR2_X1 U762 ( .A(n709), .B(KEYINPUT61), .ZN(n710) );
  NAND2_X1 U763 ( .A1(n710), .A2(G898), .ZN(n713) );
  OR2_X1 U764 ( .A1(G953), .A2(n711), .ZN(n712) );
  NAND2_X1 U765 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U766 ( .A(n715), .B(n714), .ZN(n716) );
  XNOR2_X1 U767 ( .A(KEYINPUT126), .B(n716), .ZN(G69) );
  XNOR2_X1 U768 ( .A(n718), .B(n717), .ZN(n721) );
  NAND2_X1 U769 ( .A1(n720), .A2(n719), .ZN(n725) );
  XNOR2_X1 U770 ( .A(G227), .B(n721), .ZN(n722) );
  NAND2_X1 U771 ( .A1(n722), .A2(G900), .ZN(n723) );
  NAND2_X1 U772 ( .A1(G953), .A2(n723), .ZN(n724) );
  NAND2_X1 U773 ( .A1(n725), .A2(n724), .ZN(G72) );
  XOR2_X1 U774 ( .A(n726), .B(G122), .Z(G24) );
  XOR2_X1 U775 ( .A(G119), .B(n727), .Z(G21) );
  XOR2_X1 U776 ( .A(G137), .B(n728), .Z(n729) );
  XNOR2_X1 U777 ( .A(KEYINPUT127), .B(n729), .ZN(G39) );
  XNOR2_X1 U778 ( .A(G131), .B(n730), .ZN(G33) );
endmodule

