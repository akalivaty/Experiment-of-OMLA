//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1242, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0006(.A(G250), .ZN(new_n207));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  INV_X1    g0014(.A(G264), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n207), .B(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT65), .B(KEYINPUT0), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n209), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G50), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(new_n216), .A2(new_n217), .B1(new_n219), .B2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n225), .B1(new_n216), .B2(new_n217), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  INV_X1    g0027(.A(G238), .ZN(new_n228));
  INV_X1    g0028(.A(G87), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n227), .B1(new_n221), .B2(new_n228), .C1(new_n229), .C2(new_n207), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n231));
  INV_X1    g0031(.A(G77), .ZN(new_n232));
  INV_X1    g0032(.A(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G107), .ZN(new_n234));
  OAI221_X1 g0034(.A(new_n231), .B1(new_n232), .B2(new_n233), .C1(new_n234), .C2(new_n215), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n211), .B1(new_n230), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT1), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n226), .A2(new_n237), .ZN(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT66), .B(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n202), .A2(G68), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n221), .A2(G50), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G58), .B(G77), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n250), .B(new_n255), .ZN(G351));
  AOI21_X1  g0056(.A(new_n218), .B1(G33), .B2(G41), .ZN(new_n257));
  INV_X1    g0057(.A(G274), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n259));
  NOR3_X1   g0059(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  INV_X1    g0062(.A(G45), .ZN(new_n263));
  AOI21_X1  g0063(.A(G1), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n261), .B1(new_n228), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  OAI211_X1 g0068(.A(G1), .B(G13), .C1(new_n268), .C2(new_n262), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  INV_X1    g0070(.A(G226), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n270), .B(new_n273), .C1(G232), .C2(new_n272), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G97), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n269), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n267), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT13), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n277), .B(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G169), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT14), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n277), .A2(new_n278), .ZN(new_n282));
  OR2_X1    g0082(.A1(new_n282), .A2(KEYINPUT74), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(KEYINPUT74), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n277), .A2(new_n278), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n283), .A2(new_n284), .A3(G179), .A4(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT14), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n279), .A2(new_n287), .A3(G169), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n281), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n221), .A2(G20), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n209), .A2(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n209), .A2(new_n268), .ZN(new_n292));
  OAI221_X1 g0092(.A(new_n290), .B1(new_n291), .B2(new_n232), .C1(new_n202), .C2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n218), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT11), .ZN(new_n297));
  INV_X1    g0097(.A(G13), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n298), .A2(new_n209), .A3(G1), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n221), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT12), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  AOI211_X1 g0102(.A(new_n295), .B(new_n299), .C1(new_n208), .C2(G20), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(new_n221), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n296), .A2(KEYINPUT11), .ZN(new_n306));
  NOR3_X1   g0106(.A1(new_n302), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n289), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND4_X1  g0110(.A1(new_n283), .A2(new_n284), .A3(G190), .A4(new_n285), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n279), .A2(G200), .ZN(new_n312));
  AND3_X1   g0112(.A1(new_n311), .A2(new_n307), .A3(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n310), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n270), .A2(G232), .A3(new_n272), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(new_n234), .B2(new_n270), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n270), .A2(G1698), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT67), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n317), .B(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n316), .B1(new_n319), .B2(G238), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(new_n269), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n261), .B1(new_n233), .B2(new_n266), .ZN(new_n322));
  OR2_X1    g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G169), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n321), .A2(new_n322), .ZN(new_n326));
  INV_X1    g0126(.A(G179), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(G20), .A2(G77), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT15), .B(G87), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT8), .B(G58), .ZN(new_n331));
  OAI221_X1 g0131(.A(new_n329), .B1(new_n330), .B2(new_n291), .C1(new_n292), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n295), .ZN(new_n333));
  OR2_X1    g0133(.A1(new_n333), .A2(KEYINPUT69), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(KEYINPUT69), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n299), .A2(new_n232), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n304), .B2(new_n232), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT70), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n336), .A2(KEYINPUT70), .A3(new_n339), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n325), .B(new_n328), .C1(new_n340), .C2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n323), .A2(G200), .ZN(new_n344));
  INV_X1    g0144(.A(new_n340), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n326), .A2(G190), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n344), .A2(new_n345), .A3(new_n341), .A4(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n303), .A2(G50), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n299), .A2(new_n202), .ZN(new_n350));
  INV_X1    g0150(.A(new_n295), .ZN(new_n351));
  INV_X1    g0151(.A(G150), .ZN(new_n352));
  OAI22_X1  g0152(.A1(new_n331), .A2(new_n291), .B1(new_n352), .B2(new_n292), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(G20), .B2(new_n203), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n349), .B(new_n350), .C1(new_n351), .C2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n270), .A2(G222), .A3(new_n272), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n232), .B2(new_n270), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(new_n319), .B2(G223), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n358), .A2(new_n269), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n261), .B1(new_n271), .B2(new_n266), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n355), .B1(new_n361), .B2(G169), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT68), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT68), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n364), .B(new_n355), .C1(new_n361), .C2(G169), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n361), .A2(new_n327), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  OR2_X1    g0167(.A1(new_n358), .A2(new_n269), .ZN(new_n368));
  INV_X1    g0168(.A(new_n360), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(G190), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT71), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT71), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n361), .A2(new_n373), .A3(G190), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G200), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(new_n368), .B2(new_n369), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT10), .B1(new_n377), .B2(KEYINPUT72), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n355), .A2(KEYINPUT9), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n355), .A2(KEYINPUT9), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n370), .A2(G200), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n375), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n378), .B1(new_n375), .B2(new_n381), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n348), .B(new_n367), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n314), .B1(new_n385), .B2(KEYINPUT73), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT73), .ZN(new_n387));
  AND3_X1   g0187(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n388));
  INV_X1    g0188(.A(new_n374), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n373), .B1(new_n361), .B2(G190), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n381), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n378), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n388), .B1(new_n393), .B2(new_n382), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n387), .B1(new_n394), .B2(new_n348), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT7), .ZN(new_n396));
  NOR3_X1   g0196(.A1(new_n270), .A2(new_n396), .A3(G20), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n268), .A2(KEYINPUT3), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT3), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G33), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT7), .B1(new_n401), .B2(new_n209), .ZN(new_n402));
  OAI21_X1  g0202(.A(G68), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT79), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AND2_X1   g0205(.A1(G58), .A2(G68), .ZN(new_n406));
  OAI21_X1  g0206(.A(G20), .B1(new_n406), .B2(new_n201), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT77), .ZN(new_n408));
  INV_X1    g0208(.A(G159), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n407), .A2(new_n408), .B1(new_n409), .B2(new_n292), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G58), .A2(G68), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n222), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT77), .B1(new_n412), .B2(G20), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n396), .B1(new_n270), .B2(G20), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n401), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n221), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT79), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n405), .A2(new_n414), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT16), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n351), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT75), .B1(new_n399), .B2(G33), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT75), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n423), .A2(new_n268), .A3(KEYINPUT3), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n422), .A2(new_n424), .A3(new_n400), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n209), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n396), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n425), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(KEYINPUT76), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT7), .B1(new_n425), .B2(new_n209), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT76), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n221), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  AND4_X1   g0233(.A1(KEYINPUT78), .A2(new_n433), .A3(KEYINPUT16), .A4(new_n414), .ZN(new_n434));
  OR2_X1    g0234(.A1(new_n410), .A2(new_n413), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(new_n429), .B2(new_n432), .ZN(new_n436));
  AOI21_X1  g0236(.A(KEYINPUT78), .B1(new_n436), .B2(KEYINPUT16), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n421), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n331), .A2(new_n299), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n304), .B2(new_n331), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n260), .B1(G232), .B2(new_n265), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT80), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  AOI211_X1 g0244(.A(KEYINPUT80), .B(new_n260), .C1(G232), .C2(new_n265), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n271), .A2(G1698), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(G223), .B2(G1698), .ZN(new_n448));
  OAI22_X1  g0248(.A1(new_n425), .A2(new_n448), .B1(new_n268), .B2(new_n229), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n257), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n446), .A2(new_n371), .A3(new_n450), .ZN(new_n451));
  AND2_X1   g0251(.A1(new_n442), .A2(new_n450), .ZN(new_n452));
  OR2_X1    g0252(.A1(new_n452), .A2(G200), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  AND3_X1   g0254(.A1(new_n438), .A2(new_n441), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT17), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n452), .A2(G169), .ZN(new_n457));
  AOI21_X1  g0257(.A(G179), .B1(new_n449), .B2(new_n257), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n457), .B1(new_n446), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n414), .B1(new_n417), .B2(KEYINPUT79), .ZN(new_n460));
  AOI211_X1 g0260(.A(new_n404), .B(new_n221), .C1(new_n415), .C2(new_n416), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n420), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n295), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n425), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n464));
  NOR3_X1   g0264(.A1(new_n464), .A2(new_n430), .A3(new_n431), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n426), .A2(new_n431), .A3(new_n396), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G68), .ZN(new_n467));
  OAI211_X1 g0267(.A(KEYINPUT16), .B(new_n414), .C1(new_n465), .C2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT78), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n436), .A2(KEYINPUT78), .A3(KEYINPUT16), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n463), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n459), .B1(new_n472), .B2(new_n440), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(KEYINPUT18), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n446), .A2(new_n458), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(G169), .B2(new_n452), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n476), .B1(new_n438), .B2(new_n441), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT18), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n438), .A2(new_n441), .A3(new_n454), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT17), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n456), .A2(new_n474), .A3(new_n479), .A4(new_n482), .ZN(new_n483));
  NOR3_X1   g0283(.A1(new_n386), .A2(new_n395), .A3(new_n483), .ZN(new_n484));
  AND3_X1   g0284(.A1(new_n422), .A2(new_n424), .A3(new_n400), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(new_n209), .A3(G68), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT19), .ZN(new_n487));
  NOR2_X1   g0287(.A1(G97), .A2(G107), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n229), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n275), .A2(new_n209), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n487), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(G97), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n291), .A2(KEYINPUT19), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n486), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n494), .A2(new_n295), .B1(new_n299), .B2(new_n330), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n268), .A2(G1), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n299), .A2(new_n295), .A3(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n495), .B1(new_n229), .B2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT82), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n485), .A2(new_n500), .A3(G244), .A4(G1698), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n422), .A2(new_n424), .A3(G244), .A4(new_n400), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT82), .B1(new_n502), .B2(new_n272), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(G116), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n268), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n228), .A2(G1698), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n422), .A2(new_n424), .A3(new_n400), .A4(new_n508), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n509), .A2(KEYINPUT81), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n509), .A2(KEYINPUT81), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(KEYINPUT83), .B1(new_n504), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT81), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n485), .A2(new_n514), .A3(new_n508), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n509), .A2(KEYINPUT81), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n506), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n501), .A2(new_n503), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT83), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n513), .A2(new_n520), .A3(new_n257), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n257), .A2(new_n258), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n263), .A2(G1), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n269), .B(G250), .C1(G1), .C2(new_n263), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n521), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n499), .B1(new_n528), .B2(G200), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n517), .A2(new_n518), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n269), .B1(new_n530), .B2(KEYINPUT83), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n526), .B1(new_n531), .B2(new_n520), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT86), .B1(new_n532), .B2(G190), .ZN(new_n533));
  AND4_X1   g0333(.A1(KEYINPUT86), .A2(new_n521), .A3(G190), .A4(new_n527), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n529), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT84), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n521), .A2(G179), .A3(new_n527), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n324), .B1(new_n521), .B2(new_n527), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n537), .B(KEYINPUT84), .C1(new_n324), .C2(new_n532), .ZN(new_n541));
  OR2_X1    g0341(.A1(new_n498), .A2(new_n330), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n495), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT85), .ZN(new_n544));
  XNOR2_X1  g0344(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n540), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n214), .A2(G1698), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n547), .B1(G250), .B2(G1698), .ZN(new_n548));
  INV_X1    g0348(.A(G294), .ZN(new_n549));
  OAI22_X1  g0349(.A1(new_n425), .A2(new_n548), .B1(new_n268), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n257), .ZN(new_n551));
  XNOR2_X1  g0351(.A(KEYINPUT5), .B(G41), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n257), .B1(new_n523), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G264), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n551), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n552), .A2(new_n269), .A3(G274), .A4(new_n523), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n324), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT23), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n209), .B2(G107), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n234), .A2(KEYINPUT23), .A3(G20), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n560), .A2(new_n561), .B1(new_n506), .B2(new_n209), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n401), .A2(G20), .A3(new_n229), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n562), .B1(new_n563), .B2(KEYINPUT22), .ZN(new_n564));
  NAND2_X1  g0364(.A1(KEYINPUT22), .A2(G87), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n425), .A2(G20), .A3(new_n565), .ZN(new_n566));
  OR3_X1    g0366(.A1(new_n564), .A2(new_n566), .A3(KEYINPUT24), .ZN(new_n567));
  OAI21_X1  g0367(.A(KEYINPUT24), .B1(new_n564), .B2(new_n566), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n351), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT25), .B1(new_n299), .B2(new_n234), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n299), .A2(KEYINPUT25), .A3(new_n234), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n571), .A2(new_n572), .B1(new_n497), .B2(G107), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI221_X1 g0374(.A(new_n558), .B1(G179), .B2(new_n557), .C1(new_n569), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n401), .A2(G303), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n214), .A2(new_n272), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n215), .A2(G1698), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n576), .B1(new_n425), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT87), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT87), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n576), .B(new_n582), .C1(new_n425), .C2(new_n579), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n257), .ZN(new_n585));
  NAND2_X1  g0385(.A1(G33), .A2(G283), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n586), .B(new_n209), .C1(G33), .C2(new_n492), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n505), .A2(G20), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n587), .A2(new_n295), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT20), .ZN(new_n590));
  XNOR2_X1  g0390(.A(new_n589), .B(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n299), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n592), .A2(G116), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n497), .B2(G116), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(KEYINPUT5), .A2(G41), .ZN(new_n596));
  NOR2_X1   g0396(.A1(KEYINPUT5), .A2(G41), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n523), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n598), .A2(G270), .A3(new_n269), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n599), .A2(new_n556), .A3(G179), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n585), .A2(new_n595), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n269), .B1(new_n581), .B2(new_n583), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n599), .A2(new_n556), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n595), .A2(G169), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT21), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n324), .B1(new_n591), .B2(new_n594), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT21), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n607), .B(new_n608), .C1(new_n602), .C2(new_n603), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n601), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT88), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n595), .B1(new_n604), .B2(G190), .ZN(new_n612));
  OAI21_X1  g0412(.A(G200), .B1(new_n602), .B2(new_n603), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n603), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n585), .A2(G190), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n595), .ZN(new_n617));
  AND4_X1   g0417(.A1(new_n611), .A2(new_n616), .A3(new_n617), .A4(new_n613), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n575), .B(new_n610), .C1(new_n614), .C2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n553), .A2(G257), .ZN(new_n620));
  NAND2_X1  g0420(.A1(G250), .A2(G1698), .ZN(new_n621));
  NAND2_X1  g0421(.A1(KEYINPUT4), .A2(G244), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n621), .B1(new_n622), .B2(G1698), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n586), .B1(new_n624), .B2(new_n401), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n424), .A2(new_n400), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n626), .A2(G244), .A3(new_n272), .A4(new_n422), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT4), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n620), .B1(new_n629), .B2(new_n269), .ZN(new_n630));
  INV_X1    g0430(.A(new_n556), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n327), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n299), .A2(new_n492), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n498), .B2(new_n492), .ZN(new_n635));
  OAI21_X1  g0435(.A(G107), .B1(new_n397), .B2(new_n402), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT6), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n492), .A2(new_n234), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n637), .B1(new_n638), .B2(new_n488), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n234), .A2(KEYINPUT6), .A3(G97), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G20), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n636), .B(new_n642), .C1(new_n232), .C2(new_n292), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n635), .B1(new_n643), .B2(new_n295), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n633), .B(new_n645), .C1(G169), .C2(new_n632), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n632), .A2(G190), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n647), .B(new_n644), .C1(new_n376), .C2(new_n632), .ZN(new_n648));
  INV_X1    g0448(.A(new_n569), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n555), .A2(G190), .A3(new_n556), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n557), .A2(G200), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n649), .A2(new_n573), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n646), .A2(new_n648), .A3(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n619), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n484), .A2(new_n535), .A3(new_n546), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT89), .ZN(G372));
  OAI21_X1  g0456(.A(new_n545), .B1(new_n538), .B2(new_n539), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT26), .ZN(new_n658));
  INV_X1    g0458(.A(new_n646), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n535), .A2(new_n657), .A3(new_n658), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n657), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n546), .A2(new_n535), .A3(new_n659), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n661), .B1(KEYINPUT26), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT90), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n535), .A2(new_n657), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n664), .B1(new_n665), .B2(new_n653), .ZN(new_n666));
  INV_X1    g0466(.A(new_n653), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n667), .A2(new_n535), .A3(KEYINPUT90), .A4(new_n657), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n575), .A2(new_n610), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n666), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n663), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n484), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n309), .B1(new_n343), .B2(new_n313), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n480), .B(KEYINPUT17), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n474), .A2(new_n479), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n393), .A2(new_n382), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n388), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n672), .A2(new_n679), .ZN(G369));
  NAND3_X1  g0480(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(KEYINPUT27), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G213), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n595), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g0487(.A(new_n687), .B(KEYINPUT91), .Z(new_n688));
  OAI211_X1 g0488(.A(new_n610), .B(new_n688), .C1(new_n614), .C2(new_n618), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n610), .B2(new_n688), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n569), .A2(new_n574), .ZN(new_n693));
  INV_X1    g0493(.A(new_n686), .ZN(new_n694));
  OAI211_X1 g0494(.A(new_n575), .B(new_n652), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n575), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n575), .A2(new_n686), .ZN(new_n698));
  INV_X1    g0498(.A(new_n695), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n610), .A2(new_n686), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n697), .A2(new_n701), .ZN(G399));
  NOR2_X1   g0502(.A1(new_n213), .A2(G41), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n489), .A2(G116), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(G1), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n223), .B2(new_n704), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n535), .A2(new_n657), .A3(KEYINPUT26), .A4(new_n659), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n710), .B1(new_n658), .B2(new_n662), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n667), .A2(new_n535), .A3(new_n657), .A4(new_n669), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n657), .ZN(new_n713));
  OAI211_X1 g0513(.A(KEYINPUT29), .B(new_n694), .C1(new_n711), .C2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n686), .B1(new_n663), .B2(new_n670), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n714), .B1(new_n715), .B2(KEYINPUT29), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT31), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n600), .A2(new_n551), .A3(new_n554), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n630), .A2(new_n602), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n521), .A2(new_n719), .A3(new_n527), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n532), .A2(KEYINPUT30), .A3(new_n719), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n557), .B1(new_n631), .B2(new_n630), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n585), .A2(new_n615), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n327), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n532), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n725), .B1(new_n728), .B2(KEYINPUT92), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT92), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n532), .B2(new_n727), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n724), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n717), .B1(new_n732), .B2(new_n694), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n654), .A2(new_n546), .A3(new_n535), .A4(new_n694), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n528), .A2(KEYINPUT92), .A3(new_n327), .A4(new_n726), .ZN(new_n735));
  INV_X1    g0535(.A(new_n725), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n735), .A2(new_n731), .A3(new_n736), .ZN(new_n737));
  OAI211_X1 g0537(.A(KEYINPUT31), .B(new_n686), .C1(new_n737), .C2(new_n724), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n733), .A2(new_n734), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G330), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n716), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n708), .B1(new_n742), .B2(G1), .ZN(G364));
  NOR2_X1   g0543(.A1(new_n298), .A2(G20), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n208), .B1(new_n744), .B2(G45), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n703), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n692), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(G330), .B2(new_n690), .ZN(new_n749));
  INV_X1    g0549(.A(new_n747), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n218), .B1(G20), .B2(new_n324), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n209), .A2(new_n327), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n754), .A2(G190), .A3(G200), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n371), .A2(new_n376), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n755), .A2(G311), .B1(new_n758), .B2(G326), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G179), .A2(G200), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G190), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n759), .B1(new_n549), .B2(new_n763), .ZN(new_n764));
  XOR2_X1   g0564(.A(new_n764), .B(KEYINPUT94), .Z(new_n765));
  NOR3_X1   g0565(.A1(new_n754), .A2(new_n371), .A3(G200), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n270), .B1(new_n766), .B2(G322), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n209), .A2(G179), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n756), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n760), .A2(G20), .A3(new_n371), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n770), .A2(G303), .B1(new_n772), .B2(G329), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n376), .A2(G190), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n753), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(KEYINPUT33), .B(G317), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n768), .A2(new_n774), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n776), .A2(new_n777), .B1(new_n779), .B2(G283), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n765), .A2(new_n767), .A3(new_n773), .A4(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n755), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n782), .A2(new_n232), .B1(new_n778), .B2(new_n234), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n401), .B(new_n783), .C1(G68), .C2(new_n776), .ZN(new_n784));
  XOR2_X1   g0584(.A(KEYINPUT93), .B(KEYINPUT32), .Z(new_n785));
  NAND3_X1  g0585(.A1(new_n772), .A2(new_n785), .A3(G159), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n785), .B1(new_n772), .B2(G159), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(G97), .B2(new_n762), .ZN(new_n788));
  OAI22_X1  g0588(.A1(new_n757), .A2(new_n202), .B1(new_n769), .B2(new_n229), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(G58), .B2(new_n766), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n784), .A2(new_n786), .A3(new_n788), .A4(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n752), .B1(new_n781), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(G13), .A2(G33), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(G20), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n751), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n213), .A2(new_n401), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n797), .A2(G355), .B1(new_n505), .B2(new_n213), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n213), .A2(new_n485), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n799), .B1(G45), .B2(new_n223), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n255), .A2(new_n263), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n798), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n750), .B(new_n792), .C1(new_n796), .C2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n795), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n803), .B1(new_n690), .B2(new_n804), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n749), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(G396));
  NOR2_X1   g0607(.A1(new_n343), .A2(new_n686), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n686), .B1(new_n340), .B2(new_n342), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n347), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n808), .B1(new_n343), .B2(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n715), .B(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n747), .B1(new_n812), .B2(new_n740), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n740), .B2(new_n812), .ZN(new_n814));
  AOI22_X1  g0614(.A1(G137), .A2(new_n758), .B1(new_n776), .B2(G150), .ZN(new_n815));
  INV_X1    g0615(.A(G143), .ZN(new_n816));
  INV_X1    g0616(.A(new_n766), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n815), .B1(new_n782), .B2(new_n409), .C1(new_n816), .C2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT34), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n818), .A2(new_n819), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n779), .A2(G68), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n772), .A2(G132), .ZN(new_n823));
  OAI211_X1 g0623(.A(new_n822), .B(new_n823), .C1(new_n202), .C2(new_n769), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n485), .B1(new_n763), .B2(new_n220), .ZN(new_n825));
  NOR4_X1   g0625(.A1(new_n820), .A2(new_n821), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(G303), .ZN(new_n827));
  INV_X1    g0627(.A(G283), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n757), .A2(new_n827), .B1(new_n775), .B2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(G116), .B2(new_n755), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n830), .B(KEYINPUT95), .Z(new_n831));
  AOI22_X1  g0631(.A1(new_n766), .A2(G294), .B1(G87), .B2(new_n779), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n234), .B2(new_n769), .ZN(new_n833));
  INV_X1    g0633(.A(G311), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n401), .B1(new_n834), .B2(new_n771), .C1(new_n763), .C2(new_n492), .ZN(new_n835));
  NOR3_X1   g0635(.A1(new_n831), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n751), .B1(new_n826), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n751), .A2(new_n793), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n750), .B1(new_n232), .B2(new_n838), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n837), .B(new_n839), .C1(new_n811), .C2(new_n794), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n814), .A2(new_n840), .ZN(G384));
  INV_X1    g0641(.A(KEYINPUT96), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n311), .A2(new_n307), .A3(new_n312), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n309), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n308), .A2(new_n686), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n309), .A2(KEYINPUT96), .A3(new_n843), .ZN(new_n847));
  NOR3_X1   g0647(.A1(new_n313), .A2(new_n289), .A3(new_n845), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n850), .A2(new_n739), .A3(new_n811), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT99), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT98), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n473), .A2(new_n480), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT37), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n470), .A2(new_n471), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n440), .B1(new_n856), .B2(new_n421), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n855), .B1(new_n857), .B2(new_n684), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n853), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n438), .A2(new_n441), .ZN(new_n860));
  INV_X1    g0660(.A(new_n684), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT37), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n862), .A2(KEYINPUT98), .A3(new_n473), .A4(new_n480), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n295), .B1(new_n434), .B2(new_n437), .ZN(new_n864));
  OAI211_X1 g0664(.A(KEYINPUT97), .B(new_n414), .C1(new_n465), .C2(new_n467), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(new_n420), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n436), .A2(KEYINPUT97), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n441), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n459), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n861), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n870), .A2(new_n871), .A3(new_n480), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n859), .A2(new_n863), .B1(new_n872), .B2(KEYINPUT37), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n871), .B1(new_n676), .B2(new_n674), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT38), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  OR2_X1    g0676(.A1(new_n866), .A2(new_n867), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n351), .B1(new_n470), .B2(new_n471), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n440), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n480), .B1(new_n879), .B2(new_n684), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n879), .A2(new_n476), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT37), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n455), .A2(new_n477), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT98), .B1(new_n883), .B2(new_n862), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n854), .A2(new_n858), .A3(new_n853), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n483), .A2(new_n861), .A3(new_n869), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT38), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n852), .B1(new_n876), .B2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n875), .B1(new_n873), .B2(new_n874), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n886), .A2(KEYINPUT38), .A3(new_n887), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n890), .A2(new_n891), .A3(KEYINPUT99), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n851), .B1(new_n889), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(KEYINPUT100), .B1(new_n893), .B2(KEYINPUT40), .ZN(new_n894));
  INV_X1    g0694(.A(new_n851), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n890), .A2(new_n891), .A3(KEYINPUT99), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT99), .B1(new_n890), .B2(new_n891), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT100), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT40), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n898), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n894), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n860), .A2(new_n861), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(new_n473), .A3(new_n480), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n859), .A2(new_n863), .B1(KEYINPUT37), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n903), .B1(new_n676), .B2(new_n674), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n875), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n891), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n895), .A2(KEYINPUT40), .A3(new_n908), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n902), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n484), .A2(new_n739), .ZN(new_n911));
  OAI21_X1  g0711(.A(G330), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n912), .A2(KEYINPUT101), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n910), .A2(new_n911), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n912), .B2(KEYINPUT101), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n676), .A2(new_n861), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n890), .A2(new_n891), .A3(KEYINPUT39), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT39), .B1(new_n907), .B2(new_n891), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n309), .A2(new_n686), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n846), .A2(new_n849), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n715), .A2(new_n811), .ZN(new_n923));
  INV_X1    g0723(.A(new_n808), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n897), .B2(new_n896), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n921), .A2(new_n926), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n484), .B(new_n714), .C1(new_n715), .C2(KEYINPUT29), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n679), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n927), .B(new_n929), .ZN(new_n930));
  NOR3_X1   g0730(.A1(new_n913), .A2(new_n915), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n744), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n931), .B1(G1), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n930), .B1(new_n913), .B2(new_n915), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n934), .A2(KEYINPUT102), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(KEYINPUT102), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n933), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n641), .A2(KEYINPUT35), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n641), .A2(KEYINPUT35), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n938), .A2(G116), .A3(new_n219), .A4(new_n939), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n940), .B(KEYINPUT36), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n411), .A2(G77), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n251), .B1(new_n223), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n943), .A2(G1), .A3(new_n298), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n937), .A2(new_n941), .A3(new_n944), .ZN(G367));
  NAND2_X1  g0745(.A1(new_n659), .A2(new_n686), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n646), .B(new_n648), .C1(new_n644), .C2(new_n694), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n948), .A2(new_n699), .A3(new_n700), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n949), .A2(KEYINPUT42), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT103), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n947), .A2(new_n575), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n686), .B1(new_n952), .B2(new_n646), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n949), .B2(KEYINPUT42), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n499), .A2(new_n686), .ZN(new_n956));
  MUX2_X1   g0756(.A(new_n657), .B(new_n665), .S(new_n956), .Z(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT43), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT104), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT43), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n951), .A2(new_n962), .A3(new_n954), .A4(new_n957), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n955), .A2(KEYINPUT104), .A3(new_n958), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n961), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT105), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n961), .A2(new_n963), .A3(KEYINPUT105), .A4(new_n964), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n948), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n969), .B1(new_n697), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT106), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n972), .A2(KEYINPUT44), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n972), .A2(KEYINPUT44), .ZN(new_n974));
  OR4_X1    g0774(.A1(new_n701), .A2(new_n973), .A3(new_n948), .A4(new_n974), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n972), .B(KEYINPUT44), .C1(new_n701), .C2(new_n948), .ZN(new_n976));
  AND3_X1   g0776(.A1(new_n701), .A2(KEYINPUT45), .A3(new_n948), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT45), .B1(new_n701), .B2(new_n948), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n975), .B(new_n976), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(KEYINPUT107), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(new_n697), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n699), .A2(new_n700), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n696), .B2(new_n700), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(new_n691), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n742), .B1(new_n981), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n703), .B(KEYINPUT41), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n745), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n697), .A2(new_n970), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n967), .A2(new_n989), .A3(new_n968), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n971), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  AND2_X1   g0791(.A1(new_n957), .A2(new_n795), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n799), .A2(new_n246), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n993), .B(new_n796), .C1(new_n212), .C2(new_n330), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n425), .B1(new_n834), .B2(new_n757), .C1(new_n782), .C2(new_n828), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n817), .A2(new_n827), .B1(new_n492), .B2(new_n778), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n770), .A2(KEYINPUT46), .A3(G116), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT46), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n769), .B2(new_n505), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n997), .B(new_n999), .C1(new_n234), .C2(new_n763), .ZN(new_n1000));
  INV_X1    g0800(.A(G317), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n775), .A2(new_n549), .B1(new_n771), .B2(new_n1001), .ZN(new_n1002));
  NOR4_X1   g0802(.A1(new_n995), .A2(new_n996), .A3(new_n1000), .A4(new_n1002), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n817), .A2(new_n352), .B1(new_n221), .B2(new_n763), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n1004), .A2(KEYINPUT108), .B1(new_n816), .B2(new_n757), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(KEYINPUT108), .B2(new_n1004), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT109), .Z(new_n1007));
  AOI22_X1  g0807(.A1(new_n779), .A2(G77), .B1(new_n772), .B2(G137), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n220), .B2(new_n769), .C1(new_n782), .C2(new_n202), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n401), .B(new_n1009), .C1(G159), .C2(new_n776), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1003), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT110), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT47), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n747), .B(new_n994), .C1(new_n1013), .C2(new_n752), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n991), .B1(new_n992), .B2(new_n1014), .ZN(G387));
  NAND2_X1  g0815(.A1(new_n741), .A2(new_n984), .ZN(new_n1016));
  AND2_X1   g0816(.A1(new_n1016), .A2(KEYINPUT111), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n984), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n742), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1016), .A2(KEYINPUT111), .ZN(new_n1021));
  NOR4_X1   g0821(.A1(new_n1017), .A2(new_n1020), .A3(new_n1021), .A4(new_n704), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  OR2_X1    g0823(.A1(new_n696), .A2(new_n804), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n705), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n797), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(G107), .B2(new_n212), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n243), .A2(G45), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n799), .ZN(new_n1029));
  AOI211_X1 g0829(.A(G45), .B(new_n1025), .C1(G68), .C2(G77), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n331), .A2(G50), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT50), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1029), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1027), .B1(new_n1028), .B2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n796), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n747), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n817), .A2(new_n202), .B1(new_n352), .B2(new_n771), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G68), .B2(new_n755), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n758), .A2(G159), .B1(new_n779), .B2(G97), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n331), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G77), .A2(new_n770), .B1(new_n776), .B2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n763), .A2(new_n330), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1042), .A2(new_n425), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .A4(new_n1043), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n779), .A2(G116), .B1(new_n772), .B2(G326), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n763), .A2(new_n828), .B1(new_n769), .B2(new_n549), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G322), .A2(new_n758), .B1(new_n776), .B2(G311), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n782), .B2(new_n827), .C1(new_n1001), .C2(new_n817), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT48), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1046), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n1049), .B2(new_n1048), .ZN(new_n1051));
  INV_X1    g0851(.A(KEYINPUT49), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n425), .B(new_n1045), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1044), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1036), .B1(new_n1055), .B2(new_n751), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1018), .A2(new_n746), .B1(new_n1024), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1023), .A2(new_n1057), .ZN(G393));
  XOR2_X1   g0858(.A(new_n979), .B(new_n697), .Z(new_n1059));
  NAND2_X1  g0859(.A1(new_n1019), .A2(new_n1059), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1060), .B(new_n703), .C1(new_n1019), .C2(new_n981), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1059), .A2(new_n745), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n796), .B1(new_n492), .B2(new_n212), .C1(new_n1029), .C2(new_n250), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n1063), .A2(new_n747), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n270), .B1(new_n779), .B2(G107), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1065), .B1(new_n827), .B2(new_n775), .C1(new_n782), .C2(new_n549), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(G116), .B2(new_n762), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n766), .A2(G311), .B1(new_n758), .B2(G317), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT52), .Z(new_n1069));
  AOI22_X1  g0869(.A1(new_n770), .A2(G283), .B1(new_n772), .B2(G322), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT112), .Z(new_n1071));
  NAND3_X1  g0871(.A1(new_n1067), .A2(new_n1069), .A3(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n766), .A2(G159), .B1(new_n758), .B2(G150), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT51), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n775), .A2(new_n202), .B1(new_n771), .B2(new_n816), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n1040), .B2(new_n755), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n762), .A2(G77), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n769), .A2(new_n221), .B1(new_n778), .B2(new_n229), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1078), .A2(new_n425), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1072), .B1(new_n1074), .B2(new_n1080), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT113), .Z(new_n1082));
  OAI221_X1 g0882(.A(new_n1064), .B1(new_n948), .B2(new_n804), .C1(new_n1082), .C2(new_n752), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1061), .A2(new_n1062), .A3(new_n1083), .ZN(G390));
  NAND2_X1  g0884(.A1(new_n810), .A2(new_n343), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n694), .B(new_n1085), .C1(new_n711), .C2(new_n713), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n922), .B1(new_n1086), .B2(new_n924), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n920), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n908), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(KEYINPUT114), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT114), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n920), .B1(new_n907), .B2(new_n891), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n662), .A2(new_n658), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n709), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n713), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n686), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n808), .B1(new_n1096), .B2(new_n1085), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1091), .B(new_n1092), .C1(new_n1097), .C2(new_n922), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1090), .A2(new_n1098), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n925), .A2(new_n920), .B1(new_n918), .B2(new_n917), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n739), .A2(G330), .A3(new_n811), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1101), .A2(new_n922), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1102), .A2(KEYINPUT115), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n1099), .A2(new_n1100), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1103), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n746), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n838), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n747), .B1(new_n1040), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n769), .A2(new_n352), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT53), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n766), .A2(G132), .B1(new_n758), .B2(G128), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1110), .B(new_n1111), .C1(new_n202), .C2(new_n778), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(KEYINPUT54), .B(G143), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n401), .B1(new_n755), .B2(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n776), .A2(G137), .B1(new_n772), .B2(G125), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1115), .B(new_n1116), .C1(new_n409), .C2(new_n763), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n758), .A2(G283), .B1(G294), .B2(new_n772), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n1118), .B1(new_n234), .B2(new_n775), .C1(new_n782), .C2(new_n492), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n766), .A2(G116), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n270), .B1(new_n770), .B2(G87), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1120), .A2(new_n1121), .A3(new_n822), .A4(new_n1077), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n1112), .A2(new_n1117), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1108), .B1(new_n1123), .B2(new_n751), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n919), .B2(new_n794), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1106), .A2(new_n1125), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1126), .A2(KEYINPUT117), .ZN(new_n1127));
  INV_X1    g0927(.A(KEYINPUT117), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n1106), .B2(new_n1125), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n484), .A2(G330), .A3(new_n739), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n928), .A2(new_n679), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1102), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT116), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1101), .A2(new_n1134), .A3(new_n922), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1134), .B1(new_n1101), .B2(new_n922), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1133), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n923), .A2(new_n924), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1101), .A2(new_n922), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1133), .A2(new_n1097), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1132), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n704), .B1(new_n1130), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1143), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n1127), .A2(new_n1129), .B1(new_n1146), .B2(new_n1148), .ZN(G378));
  INV_X1    g0949(.A(new_n1132), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n355), .A2(new_n861), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n394), .B(new_n1152), .Z(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n909), .A2(G330), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1156), .B1(new_n902), .B2(new_n1158), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1157), .B(new_n1155), .C1(new_n894), .C2(new_n901), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n927), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n893), .A2(KEYINPUT100), .A3(KEYINPUT40), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n899), .B1(new_n898), .B2(new_n900), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1158), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n1155), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n927), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n902), .A2(new_n1158), .A3(new_n1156), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1165), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1151), .A2(new_n1161), .A3(new_n1168), .A4(KEYINPUT57), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n927), .A2(KEYINPUT119), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1170), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1165), .A2(new_n1167), .A3(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(new_n1171), .A2(new_n1173), .B1(new_n1150), .B2(new_n1147), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n703), .B(new_n1169), .C1(new_n1174), .C2(KEYINPUT57), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n747), .B1(G50), .B2(new_n1107), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT118), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n770), .A2(G77), .B1(new_n772), .B2(G283), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n220), .B2(new_n778), .C1(new_n817), .C2(new_n234), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G116), .A2(new_n758), .B1(new_n776), .B2(G97), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n330), .B2(new_n782), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n763), .A2(new_n221), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n425), .A2(new_n262), .ZN(new_n1183));
  NOR4_X1   g0983(.A1(new_n1179), .A2(new_n1181), .A3(new_n1182), .A4(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(G50), .B1(new_n268), .B2(new_n262), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n1184), .A2(KEYINPUT58), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n766), .A2(G128), .B1(new_n758), .B2(G125), .ZN(new_n1187));
  INV_X1    g0987(.A(G137), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1187), .B1(new_n1188), .B2(new_n782), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G132), .A2(new_n776), .B1(new_n770), .B2(new_n1114), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n352), .B2(new_n763), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1193), .A2(KEYINPUT59), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n268), .B(new_n262), .C1(new_n778), .C2(new_n409), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G124), .B2(new_n772), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT59), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1196), .B1(new_n1192), .B2(new_n1197), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1186), .B1(KEYINPUT58), .B2(new_n1184), .C1(new_n1194), .C2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1177), .B1(new_n1199), .B2(new_n751), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n1155), .B2(new_n794), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1202), .B1(new_n1203), .B2(new_n746), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1175), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(G375));
  NAND2_X1  g1006(.A1(new_n1141), .A2(KEYINPUT116), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1102), .B1(new_n1207), .B2(new_n1135), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1139), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1132), .B(new_n1142), .C1(new_n1208), .C2(new_n1209), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1144), .A2(new_n986), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n922), .A2(new_n793), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n1212), .B(KEYINPUT120), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n270), .B1(new_n779), .B2(G77), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1214), .B1(new_n492), .B2(new_n769), .C1(new_n505), .C2(new_n775), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n782), .A2(new_n234), .B1(new_n771), .B2(new_n827), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n817), .A2(new_n828), .B1(new_n757), .B2(new_n549), .ZN(new_n1217));
  NOR4_X1   g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1042), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n770), .A2(G159), .B1(new_n772), .B2(G128), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(new_n220), .B2(new_n778), .C1(new_n817), .C2(new_n1188), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G132), .A2(new_n758), .B1(new_n776), .B2(new_n1114), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n352), .B2(new_n782), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n485), .B1(new_n763), .B2(new_n202), .ZN(new_n1223));
  NOR3_X1   g1023(.A1(new_n1220), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n751), .B1(new_n1218), .B2(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1225), .B(new_n747), .C1(G68), .C2(new_n1107), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1213), .A2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1142), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1227), .B1(new_n1228), .B2(new_n746), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1211), .A2(new_n1229), .ZN(G381));
  NAND3_X1  g1030(.A1(new_n1023), .A2(new_n806), .A3(new_n1057), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1231), .A2(G384), .ZN(new_n1232));
  XOR2_X1   g1032(.A(new_n1232), .B(KEYINPUT121), .Z(new_n1233));
  NOR2_X1   g1033(.A1(new_n1014), .A2(new_n992), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n991), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(G390), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1233), .A2(G381), .A3(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1126), .B1(new_n1145), .B2(new_n1147), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(new_n1205), .A3(new_n1240), .ZN(G407));
  NAND4_X1  g1041(.A1(new_n1205), .A2(G213), .A3(new_n685), .A4(new_n1240), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(G407), .A2(G213), .A3(new_n1242), .ZN(G409));
  INV_X1    g1043(.A(KEYINPUT123), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT122), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT60), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1246), .B1(new_n1228), .B2(new_n1150), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1210), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1245), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(KEYINPUT122), .B(new_n1210), .C1(new_n1143), .C2(new_n1246), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n704), .B1(new_n1248), .B2(KEYINPUT60), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1252), .A2(G384), .A3(new_n1229), .ZN(new_n1253));
  AOI21_X1  g1053(.A(G384), .B1(new_n1252), .B2(new_n1229), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1244), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1252), .A2(new_n1229), .ZN(new_n1256));
  INV_X1    g1056(.A(G384), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1252), .A2(G384), .A3(new_n1229), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(KEYINPUT123), .A3(new_n1259), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n685), .A2(G213), .A3(G2897), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1255), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT124), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1261), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1265), .A2(KEYINPUT125), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT125), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1267), .B(new_n1264), .C1(new_n1253), .C2(new_n1254), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n1262), .A2(new_n1263), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1175), .A2(G378), .A3(new_n1204), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1203), .A2(new_n986), .A3(new_n1151), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1161), .A2(new_n1168), .A3(new_n746), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n1201), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1240), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1270), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n685), .A2(G213), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  AND2_X1   g1077(.A1(new_n1255), .A2(new_n1260), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1278), .A2(KEYINPUT124), .A3(new_n1261), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1269), .A2(new_n1277), .A3(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1275), .A2(new_n1276), .A3(new_n1278), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(KEYINPUT62), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT61), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT62), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1275), .A2(new_n1284), .A3(new_n1276), .A4(new_n1278), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1280), .A2(new_n1282), .A3(new_n1283), .A4(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT126), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(G393), .A2(G396), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1231), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(G387), .A2(G390), .ZN(new_n1291));
  AND3_X1   g1091(.A1(new_n1288), .A2(new_n1290), .A3(new_n1291), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1290), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1286), .A2(new_n1295), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1275), .A2(KEYINPUT63), .A3(new_n1278), .A4(new_n1276), .ZN(new_n1297));
  AND2_X1   g1097(.A1(new_n1297), .A2(new_n1294), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT63), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1281), .A2(new_n1299), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1298), .A2(new_n1283), .A3(new_n1280), .A4(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1296), .A2(new_n1301), .ZN(G405));
  INV_X1    g1102(.A(new_n1270), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1240), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1304), .B1(new_n1175), .B2(new_n1204), .ZN(new_n1305));
  OAI21_X1  g1105(.A(KEYINPUT127), .B1(new_n1303), .B2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT127), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1307), .B(new_n1270), .C1(new_n1205), .C2(new_n1304), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1306), .A2(new_n1308), .A3(new_n1278), .ZN(new_n1309));
  OAI221_X1 g1109(.A(new_n1270), .B1(new_n1254), .B2(new_n1253), .C1(new_n1205), .C2(new_n1304), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n1295), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1309), .A2(new_n1310), .A3(new_n1294), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(G402));
endmodule


