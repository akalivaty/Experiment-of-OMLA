//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n570, new_n571, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT67), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n452), .B(new_n453), .Z(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n456), .A2(G567), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n454), .A2(G2106), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n459), .B1(new_n460), .B2(KEYINPUT69), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n461), .B1(KEYINPUT69), .B2(new_n460), .ZN(G319));
  OR2_X1    g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI22_X1  g040(.A1(new_n465), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(new_n471), .A3(G101), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT70), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n465), .A2(new_n467), .ZN(new_n476));
  INV_X1    g051(.A(G137), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n468), .A2(new_n478), .ZN(G160));
  AND2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n467), .B1(new_n463), .B2(new_n464), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n467), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  OAI211_X1 g065(.A(G138), .B(new_n467), .C1(new_n480), .C2(new_n481), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n493), .A2(new_n467), .A3(G138), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT72), .B1(new_n482), .B2(new_n494), .ZN(new_n495));
  AND3_X1   g070(.A1(new_n493), .A2(new_n467), .A3(G138), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT72), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n465), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n492), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n500), .A2(KEYINPUT71), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(KEYINPUT71), .ZN(new_n502));
  OAI21_X1  g077(.A(G2105), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n503), .A2(new_n505), .B1(new_n485), .B2(G126), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n499), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT73), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n499), .A2(KEYINPUT73), .A3(new_n506), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(G543), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n513), .B1(new_n514), .B2(KEYINPUT75), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(KEYINPUT5), .A3(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT74), .B(G651), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n518), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G88), .ZN(new_n525));
  OAI21_X1  g100(.A(G543), .B1(new_n521), .B2(new_n522), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(G50), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(new_n519), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n525), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(G166));
  NAND2_X1  g107(.A1(new_n527), .A2(G51), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n524), .A2(G89), .ZN(new_n534));
  AND2_X1   g109(.A1(G63), .A2(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n518), .A2(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n533), .A2(new_n534), .A3(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  NAND2_X1  g116(.A1(new_n524), .A2(G90), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n527), .A2(G52), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n519), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  NAND2_X1  g122(.A1(new_n524), .A2(G81), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n527), .A2(G43), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  OR2_X1    g125(.A1(new_n550), .A2(new_n519), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n548), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  AND2_X1   g134(.A1(new_n515), .A2(new_n517), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n524), .A2(G91), .B1(G651), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n527), .B2(G53), .ZN(new_n565));
  INV_X1    g140(.A(G53), .ZN(new_n566));
  NOR3_X1   g141(.A1(new_n526), .A2(KEYINPUT9), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n563), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT76), .ZN(G299));
  OR2_X1    g144(.A1(new_n531), .A2(KEYINPUT77), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n531), .A2(KEYINPUT77), .ZN(new_n571));
  AND2_X1   g146(.A1(new_n570), .A2(new_n571), .ZN(G303));
  NAND2_X1  g147(.A1(new_n527), .A2(G49), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n524), .A2(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n560), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n519), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(G86), .ZN(new_n582));
  INV_X1    g157(.A(G48), .ZN(new_n583));
  OAI221_X1 g158(.A(new_n581), .B1(new_n523), .B2(new_n582), .C1(new_n583), .C2(new_n526), .ZN(G305));
  NAND2_X1  g159(.A1(new_n524), .A2(G85), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n527), .A2(G47), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OAI211_X1 g162(.A(new_n585), .B(new_n586), .C1(new_n519), .C2(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  OAI211_X1 g164(.A(G92), .B(new_n518), .C1(new_n521), .C2(new_n522), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n590), .B(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(G651), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n560), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n593), .B1(new_n596), .B2(KEYINPUT78), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(KEYINPUT78), .B2(new_n596), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n527), .A2(G54), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n592), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n589), .B1(new_n601), .B2(G868), .ZN(G284));
  OAI21_X1  g177(.A(new_n589), .B1(new_n601), .B2(G868), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT76), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n568), .B(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n604), .B1(new_n606), .B2(G868), .ZN(G297));
  OAI21_X1  g182(.A(new_n604), .B1(new_n606), .B2(G868), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n601), .B1(new_n609), .B2(G860), .ZN(G148));
  NAND2_X1  g185(.A1(new_n601), .A2(new_n609), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n485), .A2(G123), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n467), .A2(G111), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  INV_X1    g192(.A(G135), .ZN(new_n618));
  OAI221_X1 g193(.A(new_n615), .B1(new_n616), .B2(new_n617), .C1(new_n618), .C2(new_n476), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT79), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2096), .Z(new_n621));
  NAND2_X1  g196(.A1(new_n465), .A2(new_n470), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(KEYINPUT13), .B(G2100), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n621), .A2(new_n625), .ZN(G156));
  XOR2_X1   g201(.A(KEYINPUT15), .B(G2435), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2438), .ZN(new_n628));
  XOR2_X1   g203(.A(G2427), .B(G2430), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT80), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n628), .A2(new_n630), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n631), .A2(KEYINPUT14), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2451), .B(G2454), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n633), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G14), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n638), .A2(new_n639), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n641), .A2(new_n642), .ZN(G401));
  XOR2_X1   g218(.A(G2067), .B(G2678), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT82), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2072), .B(G2078), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT81), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n645), .B1(KEYINPUT83), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(KEYINPUT83), .B2(new_n647), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n647), .B(KEYINPUT17), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n650), .A2(new_n645), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2084), .B(G2090), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n649), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  OR3_X1    g228(.A1(new_n650), .A2(new_n645), .A3(new_n652), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n644), .A2(new_n652), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n647), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT18), .Z(new_n657));
  NAND3_X1  g232(.A1(new_n653), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2100), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT84), .B(G2096), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  AND2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT20), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n664), .A2(new_n665), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n663), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n663), .B2(new_n669), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT85), .Z(new_n673));
  XOR2_X1   g248(.A(G1981), .B(G1986), .Z(new_n674));
  XNOR2_X1  g249(.A(G1991), .B(G1996), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n673), .B(new_n678), .ZN(G229));
  INV_X1    g254(.A(G16), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(G23), .ZN(new_n681));
  INV_X1    g256(.A(G288), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n681), .B1(new_n682), .B2(new_n680), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT89), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT33), .B(G1976), .Z(new_n685));
  OR2_X1    g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT88), .B(KEYINPUT34), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT87), .B(G16), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n689), .A2(G22), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(G166), .B2(new_n689), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(G1971), .ZN(new_n692));
  MUX2_X1   g267(.A(G6), .B(G305), .S(G16), .Z(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT32), .B(G1981), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n684), .A2(new_n685), .ZN(new_n697));
  NAND4_X1  g272(.A1(new_n686), .A2(new_n687), .A3(new_n696), .A4(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G24), .B(G290), .S(new_n689), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(G1986), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n485), .A2(G119), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n467), .A2(G107), .ZN(new_n702));
  OAI21_X1  g277(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n703));
  INV_X1    g278(.A(G131), .ZN(new_n704));
  OAI221_X1 g279(.A(new_n701), .B1(new_n702), .B2(new_n703), .C1(new_n704), .C2(new_n476), .ZN(new_n705));
  MUX2_X1   g280(.A(G25), .B(new_n705), .S(G29), .Z(new_n706));
  XOR2_X1   g281(.A(KEYINPUT35), .B(G1991), .Z(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(KEYINPUT86), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n706), .B(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n700), .A2(new_n709), .ZN(new_n710));
  AND3_X1   g285(.A1(new_n698), .A2(KEYINPUT90), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(KEYINPUT90), .B1(new_n698), .B2(new_n710), .ZN(new_n712));
  AND3_X1   g287(.A1(new_n686), .A2(new_n697), .A3(new_n696), .ZN(new_n713));
  OAI22_X1  g288(.A1(new_n711), .A2(new_n712), .B1(new_n687), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(KEYINPUT91), .A2(KEYINPUT36), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT92), .Z(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n714), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n485), .A2(G128), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n467), .A2(G116), .ZN(new_n720));
  OAI21_X1  g295(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n721));
  INV_X1    g296(.A(G140), .ZN(new_n722));
  OAI221_X1 g297(.A(new_n719), .B1(new_n720), .B2(new_n721), .C1(new_n722), .C2(new_n476), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G29), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT94), .Z(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G26), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT28), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G2067), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n689), .A2(G19), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(new_n553), .B2(new_n689), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(G1341), .Z(new_n734));
  NAND2_X1  g309(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n680), .A2(G4), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n601), .B2(new_n680), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT93), .B(G1348), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n737), .B(new_n738), .Z(new_n739));
  NOR2_X1   g314(.A1(G168), .A2(new_n680), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n680), .B2(G21), .ZN(new_n741));
  INV_X1    g316(.A(G1966), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT31), .B(G11), .Z(new_n744));
  NOR2_X1   g319(.A1(new_n620), .A2(new_n726), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT100), .B(G28), .ZN(new_n746));
  AOI21_X1  g321(.A(G29), .B1(new_n746), .B2(KEYINPUT30), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(KEYINPUT101), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n747), .A2(KEYINPUT101), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n746), .A2(KEYINPUT30), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n744), .B(new_n745), .C1(new_n748), .C2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G34), .ZN(new_n753));
  AND2_X1   g328(.A1(new_n753), .A2(KEYINPUT24), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(KEYINPUT24), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n726), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G160), .B2(new_n726), .ZN(new_n757));
  INV_X1    g332(.A(G2084), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n743), .A2(new_n752), .A3(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(G171), .A2(new_n680), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G5), .B2(new_n680), .ZN(new_n762));
  INV_X1    g337(.A(G1961), .ZN(new_n763));
  OAI22_X1  g338(.A1(new_n762), .A2(new_n763), .B1(new_n741), .B2(new_n742), .ZN(new_n764));
  NOR4_X1   g339(.A1(new_n735), .A2(new_n739), .A3(new_n760), .A4(new_n764), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n762), .A2(new_n763), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n726), .A2(G27), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT102), .Z(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G164), .B2(new_n726), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G2078), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n726), .A2(G35), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G162), .B2(new_n726), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT29), .Z(new_n773));
  INV_X1    g348(.A(G2090), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  NOR4_X1   g351(.A1(new_n766), .A2(new_n770), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n726), .A2(G33), .ZN(new_n778));
  INV_X1    g353(.A(G127), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n482), .A2(new_n779), .ZN(new_n780));
  AND2_X1   g355(.A1(G115), .A2(G2104), .ZN(new_n781));
  OAI21_X1  g356(.A(G2105), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT95), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI211_X1 g359(.A(KEYINPUT95), .B(G2105), .C1(new_n780), .C2(new_n781), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT25), .ZN(new_n786));
  NAND2_X1  g361(.A1(G103), .A2(G2104), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(G2105), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n467), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n483), .A2(G139), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n784), .A2(new_n785), .A3(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT96), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n778), .B1(new_n793), .B2(G29), .ZN(new_n794));
  INV_X1    g369(.A(G2072), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT26), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n470), .A2(G105), .ZN(new_n799));
  INV_X1    g374(.A(G141), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n476), .B2(new_n800), .ZN(new_n801));
  AOI211_X1 g376(.A(new_n798), .B(new_n801), .C1(G129), .C2(new_n485), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT98), .ZN(new_n803));
  OR3_X1    g378(.A1(new_n803), .A2(KEYINPUT99), .A3(new_n726), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(new_n726), .ZN(new_n805));
  OAI21_X1  g380(.A(KEYINPUT99), .B1(G29), .B2(G32), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT27), .B(G1996), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n765), .A2(new_n777), .A3(new_n796), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n688), .A2(G20), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT23), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n606), .B2(new_n680), .ZN(new_n813));
  INV_X1    g388(.A(G1956), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n794), .A2(new_n795), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT97), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(KEYINPUT103), .B1(new_n810), .B2(new_n818), .ZN(new_n819));
  AND3_X1   g394(.A1(new_n809), .A2(new_n777), .A3(new_n796), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT103), .ZN(new_n821));
  INV_X1    g396(.A(new_n818), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n820), .A2(new_n821), .A3(new_n822), .A4(new_n765), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n714), .A2(new_n717), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n718), .A2(new_n824), .A3(new_n825), .ZN(G150));
  INV_X1    g401(.A(G150), .ZN(G311));
  NOR2_X1   g402(.A1(new_n600), .A2(new_n609), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n518), .A2(G67), .ZN(new_n831));
  AND2_X1   g406(.A1(G80), .A2(G543), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n580), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT105), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n834), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT106), .B(G55), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n527), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n524), .A2(G93), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n835), .A2(new_n836), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n552), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n830), .B(new_n841), .Z(new_n842));
  AND2_X1   g417(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n842), .A2(KEYINPUT39), .ZN(new_n844));
  NOR3_X1   g419(.A1(new_n843), .A2(new_n844), .A3(G860), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n840), .A2(G860), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT37), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n845), .A2(new_n847), .ZN(G145));
  XNOR2_X1  g423(.A(new_n620), .B(G162), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G160), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n485), .A2(G130), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n467), .A2(G118), .ZN(new_n852));
  OAI21_X1  g427(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n853));
  INV_X1    g428(.A(G142), .ZN(new_n854));
  OAI221_X1 g429(.A(new_n851), .B1(new_n852), .B2(new_n853), .C1(new_n854), .C2(new_n476), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT107), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n623), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n705), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT108), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n793), .A2(new_n802), .ZN(new_n860));
  INV_X1    g435(.A(new_n803), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n861), .B2(new_n793), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n507), .B(new_n723), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n864), .A2(KEYINPUT108), .A3(new_n858), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n850), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n866), .B(new_n850), .C1(new_n859), .C2(new_n864), .ZN(new_n868));
  INV_X1    g443(.A(G37), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT40), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(G395));
  XNOR2_X1  g448(.A(new_n841), .B(new_n611), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n606), .A2(new_n600), .ZN(new_n875));
  NAND2_X1  g450(.A1(G299), .A2(new_n601), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT41), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n875), .A2(new_n876), .A3(KEYINPUT41), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n878), .B1(new_n883), .B2(new_n874), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  XOR2_X1   g461(.A(G288), .B(KEYINPUT109), .Z(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(G305), .ZN(new_n888));
  XNOR2_X1  g463(.A(G290), .B(new_n531), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(new_n890));
  NOR2_X1   g465(.A1(new_n890), .A2(KEYINPUT110), .ZN(new_n891));
  OAI211_X1 g466(.A(KEYINPUT42), .B(new_n878), .C1(new_n883), .C2(new_n874), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n886), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n891), .B1(new_n886), .B2(new_n892), .ZN(new_n894));
  OAI21_X1  g469(.A(G868), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(G868), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n840), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(G295));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n897), .ZN(G331));
  XNOR2_X1  g474(.A(KEYINPUT111), .B(KEYINPUT44), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n901));
  XNOR2_X1  g476(.A(G301), .B(G286), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n841), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n841), .A2(new_n902), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n904), .A2(new_n877), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n905), .A2(KEYINPUT112), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(KEYINPUT112), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n904), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n907), .B1(new_n911), .B2(new_n882), .ZN(new_n912));
  OR2_X1    g487(.A1(new_n912), .A2(new_n890), .ZN(new_n913));
  AOI21_X1  g488(.A(G37), .B1(new_n912), .B2(new_n890), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n901), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n890), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n904), .A2(new_n877), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n917), .B1(new_n909), .B2(new_n908), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n880), .A2(new_n881), .B1(new_n904), .B2(new_n905), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n903), .B1(new_n908), .B2(new_n909), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n890), .B(new_n906), .C1(new_n883), .C2(new_n921), .ZN(new_n922));
  AND4_X1   g497(.A1(new_n901), .A2(new_n920), .A3(new_n922), .A4(new_n869), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n900), .B1(new_n915), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n913), .A2(new_n901), .A3(new_n914), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n920), .A2(new_n869), .A3(new_n922), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n925), .B(KEYINPUT44), .C1(new_n926), .C2(new_n901), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n924), .A2(new_n927), .ZN(G397));
  XNOR2_X1  g503(.A(KEYINPUT113), .B(G1384), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n929), .B1(new_n499), .B2(new_n506), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n930), .A2(KEYINPUT45), .ZN(new_n931));
  INV_X1    g506(.A(G40), .ZN(new_n932));
  NOR3_X1   g507(.A1(new_n468), .A2(new_n478), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n934), .A2(G1996), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n936), .A2(new_n803), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n937), .A2(KEYINPUT114), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(KEYINPUT114), .ZN(new_n939));
  INV_X1    g514(.A(new_n934), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n723), .B(new_n730), .ZN(new_n941));
  INV_X1    g516(.A(G1996), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n941), .B1(new_n942), .B2(new_n802), .ZN(new_n943));
  AOI22_X1  g518(.A1(new_n938), .A2(new_n939), .B1(new_n940), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n707), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n705), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n705), .A2(new_n945), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n940), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(G290), .B(G1986), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n949), .B1(new_n940), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT61), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n568), .B(KEYINPUT57), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT50), .ZN(new_n955));
  INV_X1    g530(.A(G1384), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n499), .A2(KEYINPUT73), .A3(new_n506), .ZN(new_n957));
  AOI21_X1  g532(.A(KEYINPUT73), .B1(new_n499), .B2(new_n506), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n955), .B(new_n956), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT116), .ZN(new_n960));
  AOI21_X1  g535(.A(G1384), .B1(new_n499), .B2(new_n506), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n933), .B(new_n960), .C1(new_n961), .C2(new_n955), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n507), .A2(new_n956), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT50), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n960), .B1(new_n965), .B2(new_n933), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n814), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT120), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n933), .B1(new_n961), .B2(new_n955), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT116), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n970), .A2(new_n959), .A3(new_n962), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT120), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n972), .A3(new_n814), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n968), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AOI22_X1  g552(.A1(new_n483), .A2(G137), .B1(new_n474), .B2(new_n472), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n978), .B(G40), .C1(new_n467), .C2(new_n466), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n979), .B1(KEYINPUT45), .B2(new_n930), .ZN(new_n980));
  XNOR2_X1  g555(.A(KEYINPUT56), .B(G2072), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n977), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n954), .B1(new_n974), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n982), .ZN(new_n984));
  AOI211_X1 g559(.A(new_n984), .B(new_n953), .C1(new_n968), .C2(new_n973), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n952), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n979), .B1(new_n955), .B2(new_n961), .ZN(new_n987));
  AOI21_X1  g562(.A(G1384), .B1(new_n509), .B2(new_n510), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n987), .B1(new_n988), .B2(new_n955), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n738), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n933), .A2(new_n961), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(G2067), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n990), .A2(KEYINPUT60), .A3(new_n993), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n601), .A2(KEYINPUT122), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n992), .B1(new_n989), .B2(new_n738), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n601), .A2(KEYINPUT122), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n998), .A2(new_n995), .A3(KEYINPUT60), .A4(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n990), .A2(new_n993), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT60), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n997), .A2(new_n1000), .A3(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(KEYINPUT121), .B(G1996), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n977), .A2(new_n980), .A3(new_n1006), .ZN(new_n1007));
  XOR2_X1   g582(.A(KEYINPUT58), .B(G1341), .Z(new_n1008));
  NAND2_X1  g583(.A1(new_n991), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT59), .B1(new_n1010), .B2(new_n553), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT59), .ZN(new_n1012));
  AOI211_X1 g587(.A(new_n1012), .B(new_n552), .C1(new_n1007), .C2(new_n1009), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1004), .A2(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n971), .A2(new_n972), .A3(new_n814), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n972), .B1(new_n971), .B2(new_n814), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n982), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n953), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n974), .A2(new_n954), .A3(new_n982), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(KEYINPUT61), .A3(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n986), .A2(new_n1015), .A3(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n998), .A2(new_n600), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1020), .B1(new_n983), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n570), .A2(G8), .A3(new_n571), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G8), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n971), .A2(new_n1030), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n970), .A2(KEYINPUT117), .A3(new_n959), .A4(new_n962), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(new_n774), .A3(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n980), .B1(new_n988), .B2(KEYINPUT45), .ZN(new_n1034));
  INV_X1    g609(.A(G1971), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1029), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1033), .A2(KEYINPUT118), .A3(new_n1036), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1028), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g616(.A(KEYINPUT45), .B(new_n956), .C1(new_n957), .C2(new_n958), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n979), .B1(new_n964), .B2(new_n976), .ZN(new_n1043));
  INV_X1    g618(.A(G2078), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT123), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1042), .A2(new_n1043), .A3(KEYINPUT123), .A4(new_n1044), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(KEYINPUT53), .A3(new_n1048), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1044), .B(new_n980), .C1(new_n988), .C2(KEYINPUT45), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n1051));
  XNOR2_X1  g626(.A(KEYINPUT124), .B(G1961), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1050), .A2(new_n1051), .B1(new_n989), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1049), .A2(new_n1053), .A3(G301), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n931), .A2(new_n1051), .A3(G2078), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n980), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT54), .B(new_n1054), .C1(new_n1057), .C2(G301), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(new_n742), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n758), .B(new_n987), .C1(new_n988), .C2(new_n955), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(new_n1061), .A3(G168), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT51), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1063), .A2(new_n1029), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(G168), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT51), .B1(new_n1062), .B2(G8), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1058), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT115), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n774), .B(new_n987), .C1(new_n988), .C2(new_n955), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1036), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1072), .ZN(new_n1074));
  AOI21_X1  g649(.A(G1971), .B1(new_n977), .B2(new_n980), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT115), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1028), .A2(G8), .A3(new_n1073), .A4(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(G305), .A2(G1981), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n524), .A2(G86), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n527), .A2(G48), .ZN(new_n1080));
  INV_X1    g655(.A(G1981), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .A4(new_n581), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1078), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT49), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1078), .A2(KEYINPUT49), .A3(new_n1082), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n991), .A2(G8), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1085), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G1976), .ZN(new_n1090));
  NOR2_X1   g665(.A1(G288), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT52), .B1(new_n1091), .B2(new_n1087), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT52), .B1(G288), .B2(new_n1090), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1088), .B(new_n1093), .C1(new_n1090), .C2(G288), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1089), .A2(new_n1092), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1077), .A2(new_n1096), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1041), .A2(new_n1070), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1025), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(G171), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT125), .ZN(new_n1102));
  AOI21_X1  g677(.A(G301), .B1(new_n1049), .B2(new_n1053), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT125), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1057), .A2(G301), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1102), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n1107), .A2(KEYINPUT126), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT126), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1099), .A2(new_n1111), .ZN(new_n1112));
  AOI211_X1 g687(.A(new_n1029), .B(G286), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT63), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  AND2_X1   g690(.A1(new_n1062), .A2(G8), .ZN(new_n1116));
  OAI221_X1 g691(.A(KEYINPUT62), .B1(new_n1065), .B2(new_n1066), .C1(new_n1116), .C2(KEYINPUT51), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1118), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(new_n1103), .B(KEYINPUT125), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1115), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1041), .A2(new_n1097), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT119), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1076), .A2(G8), .A3(new_n1073), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1026), .B(KEYINPUT55), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1125), .B1(new_n1128), .B2(new_n1096), .ZN(new_n1129));
  AOI211_X1 g704(.A(KEYINPUT119), .B(new_n1095), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1077), .B(new_n1113), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(KEYINPUT63), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1077), .A2(new_n1095), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1089), .A2(new_n1090), .A3(new_n682), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1087), .B1(new_n1134), .B2(new_n1082), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1124), .A2(new_n1132), .A3(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n951), .B1(new_n1112), .B2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n934), .B1(new_n802), .B2(new_n941), .ZN(new_n1139));
  OR2_X1    g714(.A1(new_n936), .A2(KEYINPUT46), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n936), .A2(KEYINPUT46), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1142), .B(KEYINPUT47), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n944), .A2(new_n947), .ZN(new_n1144));
  OR2_X1    g719(.A1(new_n723), .A2(G2067), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n934), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n949), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n934), .A2(G1986), .A3(G290), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n1148), .B(KEYINPUT48), .Z(new_n1149));
  AOI211_X1 g724(.A(new_n1143), .B(new_n1146), .C1(new_n1147), .C2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1138), .A2(new_n1150), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g726(.A1(new_n915), .A2(new_n923), .ZN(new_n1153));
  OAI21_X1  g727(.A(G319), .B1(new_n641), .B2(new_n642), .ZN(new_n1154));
  NOR3_X1   g728(.A1(G227), .A2(G229), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n1156));
  XNOR2_X1  g730(.A(new_n1155), .B(new_n1156), .ZN(new_n1157));
  OAI21_X1  g731(.A(new_n1157), .B1(new_n867), .B2(new_n870), .ZN(new_n1158));
  NOR2_X1   g732(.A1(new_n1153), .A2(new_n1158), .ZN(G308));
  OAI221_X1 g733(.A(new_n1157), .B1(new_n867), .B2(new_n870), .C1(new_n915), .C2(new_n923), .ZN(G225));
endmodule


