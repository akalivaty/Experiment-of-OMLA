//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n437, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n563, new_n564, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n584, new_n585, new_n586, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n648, new_n651, new_n653, new_n654,
    new_n655, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1260, new_n1261, new_n1262, new_n1263,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1272, new_n1273, new_n1274;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(new_n437));
  INV_X1    g012(.A(new_n437), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g020(.A(KEYINPUT67), .B(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n462), .B1(new_n463), .B2(G125), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AND3_X1   g041(.A1(new_n465), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(KEYINPUT68), .B1(new_n465), .B2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(G101), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(G137), .A3(new_n465), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT69), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n469), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n466), .B1(new_n472), .B2(new_n474), .ZN(G160));
  OR2_X1    g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n476), .A2(KEYINPUT70), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT70), .ZN(new_n479));
  AND2_X1   g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NOR2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(G2105), .B1(new_n478), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n465), .B1(new_n478), .B2(new_n482), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  OR2_X1    g061(.A1(G100), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n484), .A2(new_n486), .A3(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n492));
  OAI211_X1 g067(.A(G126), .B(G2105), .C1(new_n480), .C2(new_n481), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(KEYINPUT71), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n463), .A2(new_n465), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n463), .A2(new_n499), .A3(new_n465), .A4(new_n496), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n494), .B1(new_n498), .B2(new_n500), .ZN(G164));
  OR2_X1    g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n502), .A2(new_n503), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n505), .B1(new_n502), .B2(new_n503), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n508), .A2(G88), .B1(new_n509), .B2(G50), .ZN(new_n510));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G62), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n511), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G651), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n510), .A2(new_n517), .ZN(G166));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT7), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n519), .A2(KEYINPUT7), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n508), .A2(G89), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n523), .B1(new_n512), .B2(new_n513), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n506), .A2(KEYINPUT72), .A3(new_n507), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n524), .A2(new_n525), .A3(G63), .A4(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  AND2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  OAI21_X1  g105(.A(G543), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT73), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT6), .B(G651), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n533), .A2(new_n534), .A3(G543), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n528), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n527), .A2(new_n536), .ZN(G168));
  NAND3_X1  g112(.A1(new_n524), .A2(new_n525), .A3(G64), .ZN(new_n538));
  NAND2_X1  g113(.A1(G77), .A2(G543), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(KEYINPUT74), .ZN(new_n542));
  INV_X1    g117(.A(G651), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(new_n538), .B2(new_n539), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT74), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n532), .A2(new_n535), .ZN(new_n547));
  XNOR2_X1  g122(.A(KEYINPUT75), .B(G90), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n547), .A2(G52), .B1(new_n508), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n542), .A2(new_n546), .A3(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  NAND3_X1  g126(.A1(new_n524), .A2(new_n525), .A3(G56), .ZN(new_n552));
  INV_X1    g127(.A(G68), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n553), .B2(new_n505), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G651), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n506), .A2(new_n507), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n556), .A2(new_n533), .A3(G81), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n557), .B1(new_n547), .B2(G43), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n566), .A2(G65), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(G65), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n556), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(G78), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n570), .B2(new_n505), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G651), .ZN(new_n572));
  INV_X1    g147(.A(G53), .ZN(new_n573));
  OR3_X1    g148(.A1(new_n531), .A2(KEYINPUT9), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT9), .B1(new_n531), .B2(new_n573), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n556), .A2(new_n533), .ZN(new_n577));
  INV_X1    g152(.A(G91), .ZN(new_n578));
  OAI21_X1  g153(.A(KEYINPUT76), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  NOR3_X1   g155(.A1(new_n577), .A2(KEYINPUT76), .A3(new_n578), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n572), .B(new_n576), .C1(new_n580), .C2(new_n581), .ZN(G299));
  INV_X1    g157(.A(G168), .ZN(G286));
  NAND2_X1  g158(.A1(new_n510), .A2(new_n517), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(KEYINPUT78), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(KEYINPUT78), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(G303));
  INV_X1    g162(.A(G74), .ZN(new_n588));
  NOR3_X1   g163(.A1(new_n512), .A2(new_n513), .A3(new_n523), .ZN(new_n589));
  AOI21_X1  g164(.A(KEYINPUT72), .B1(new_n506), .B2(new_n507), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n591), .A2(new_n592), .A3(G651), .ZN(new_n593));
  AOI21_X1  g168(.A(G74), .B1(new_n524), .B2(new_n525), .ZN(new_n594));
  OAI21_X1  g169(.A(KEYINPUT79), .B1(new_n594), .B2(new_n543), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G87), .ZN(new_n597));
  INV_X1    g172(.A(G49), .ZN(new_n598));
  OAI22_X1  g173(.A1(new_n577), .A2(new_n597), .B1(new_n598), .B2(new_n531), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n596), .A2(new_n600), .ZN(G288));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n602));
  INV_X1    g177(.A(G61), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n506), .B2(new_n507), .ZN(new_n604));
  NAND2_X1  g179(.A1(G73), .A2(G543), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(KEYINPUT80), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT80), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n607), .A2(G73), .A3(G543), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n602), .B(G651), .C1(new_n604), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n508), .A2(G86), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n509), .A2(G48), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n606), .B(new_n608), .C1(new_n514), .C2(new_n603), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n602), .B1(new_n614), .B2(G651), .ZN(new_n615));
  OAI21_X1  g190(.A(KEYINPUT82), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(G651), .B1(new_n604), .B2(new_n609), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(KEYINPUT81), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT82), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n508), .A2(G86), .B1(new_n509), .B2(G48), .ZN(new_n620));
  NAND4_X1  g195(.A1(new_n618), .A2(new_n619), .A3(new_n620), .A4(new_n610), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(G305));
  AOI22_X1  g198(.A1(new_n547), .A2(G47), .B1(G85), .B2(new_n508), .ZN(new_n624));
  INV_X1    g199(.A(KEYINPUT83), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n524), .A2(new_n525), .A3(G60), .ZN(new_n626));
  NAND2_X1  g201(.A1(G72), .A2(G543), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n625), .B1(new_n628), .B2(G651), .ZN(new_n629));
  AOI211_X1 g204(.A(KEYINPUT83), .B(new_n543), .C1(new_n626), .C2(new_n627), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n624), .B1(new_n629), .B2(new_n630), .ZN(G290));
  INV_X1    g206(.A(G868), .ZN(new_n632));
  OR3_X1    g207(.A1(G171), .A2(KEYINPUT84), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(KEYINPUT84), .B1(G171), .B2(new_n632), .ZN(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT85), .B(KEYINPUT10), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(G92), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n636), .B1(new_n577), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n508), .A2(G92), .A3(new_n635), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n547), .A2(G54), .ZN(new_n641));
  AND2_X1   g216(.A1(new_n556), .A2(G66), .ZN(new_n642));
  AND2_X1   g217(.A1(G79), .A2(G543), .ZN(new_n643));
  OAI21_X1  g218(.A(G651), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AND3_X1   g219(.A1(new_n640), .A2(new_n641), .A3(new_n644), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n633), .B(new_n634), .C1(G868), .C2(new_n645), .ZN(G284));
  OAI211_X1 g221(.A(new_n633), .B(new_n634), .C1(G868), .C2(new_n645), .ZN(G321));
  NAND2_X1  g222(.A1(G299), .A2(new_n632), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n648), .B1(new_n632), .B2(G168), .ZN(G297));
  OAI21_X1  g224(.A(new_n648), .B1(new_n632), .B2(G168), .ZN(G280));
  INV_X1    g225(.A(G559), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n645), .B1(new_n651), .B2(G860), .ZN(G148));
  NOR2_X1   g227(.A1(new_n559), .A2(G868), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n645), .A2(new_n651), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT86), .Z(new_n655));
  AOI21_X1  g230(.A(new_n653), .B1(new_n655), .B2(G868), .ZN(G323));
  XNOR2_X1  g231(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g232(.A(new_n463), .B1(new_n467), .B2(new_n468), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT12), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT13), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n660), .A2(G2100), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n483), .A2(G135), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n485), .A2(G123), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n465), .A2(G111), .ZN(new_n664));
  OAI21_X1  g239(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n662), .B(new_n663), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(G2096), .Z(new_n667));
  NAND2_X1  g242(.A1(new_n660), .A2(G2100), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n661), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT87), .ZN(G156));
  INV_X1    g245(.A(G14), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT15), .B(G2435), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT88), .B(G2438), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2427), .B(G2430), .Z(new_n675));
  OR2_X1    g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n675), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n676), .A2(KEYINPUT14), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2451), .B(G2454), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT16), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G2443), .B(G2446), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n682), .ZN(new_n684));
  INV_X1    g259(.A(new_n680), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n678), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n678), .A2(new_n685), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n684), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1341), .B(G1348), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n671), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n683), .A2(new_n688), .ZN(new_n693));
  AOI21_X1  g268(.A(KEYINPUT89), .B1(new_n693), .B2(new_n690), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT89), .ZN(new_n695));
  AOI211_X1 g270(.A(new_n695), .B(new_n691), .C1(new_n683), .C2(new_n688), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n692), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G401));
  XNOR2_X1  g273(.A(G2067), .B(G2678), .ZN(new_n699));
  XNOR2_X1  g274(.A(G2072), .B(G2078), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XOR2_X1   g276(.A(G2084), .B(G2090), .Z(new_n702));
  OR3_X1    g277(.A1(new_n701), .A2(KEYINPUT90), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(KEYINPUT90), .B1(new_n701), .B2(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(new_n699), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n700), .B(KEYINPUT17), .Z(new_n706));
  OAI211_X1 g281(.A(new_n703), .B(new_n704), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n702), .A2(new_n699), .A3(new_n700), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT18), .Z(new_n709));
  NAND3_X1  g284(.A1(new_n706), .A2(new_n702), .A3(new_n705), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n707), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(G2096), .B(G2100), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(G227));
  XNOR2_X1  g288(.A(G1981), .B(G1986), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(G1971), .B(G1976), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT19), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  XOR2_X1   g293(.A(G1956), .B(G2474), .Z(new_n719));
  XOR2_X1   g294(.A(G1961), .B(G1966), .Z(new_n720));
  AND2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT20), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n719), .A2(new_n720), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n718), .A2(new_n724), .ZN(new_n725));
  OR3_X1    g300(.A1(new_n718), .A2(new_n721), .A3(new_n724), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n723), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT20), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n722), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n726), .A2(new_n725), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(new_n728), .ZN(new_n735));
  XOR2_X1   g310(.A(G1991), .B(G1996), .Z(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n730), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n737), .B1(new_n730), .B2(new_n735), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n715), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n727), .A2(new_n729), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n734), .A2(new_n728), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n736), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n744), .A2(new_n714), .A3(new_n738), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n741), .A2(new_n745), .ZN(G229));
  OAI21_X1  g321(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n747));
  INV_X1    g322(.A(G107), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(G2105), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT92), .ZN(new_n750));
  OR2_X1    g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n751), .A2(new_n752), .B1(new_n483), .B2(G131), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT91), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n485), .A2(new_n754), .A3(G119), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n754), .B1(new_n485), .B2(G119), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n753), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  MUX2_X1   g333(.A(G25), .B(new_n758), .S(G29), .Z(new_n759));
  XOR2_X1   g334(.A(KEYINPUT35), .B(G1991), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G16), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(G24), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n547), .A2(G47), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n508), .A2(G85), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n628), .A2(G651), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(KEYINPUT83), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n628), .A2(new_n625), .A3(G651), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n766), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n763), .B1(new_n770), .B2(new_n762), .ZN(new_n771));
  OR2_X1    g346(.A1(new_n771), .A2(G1986), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(G1986), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n761), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n762), .A2(G22), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G166), .B2(new_n762), .ZN(new_n776));
  INV_X1    g351(.A(G1971), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n776), .B(new_n777), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n762), .A2(G23), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G288), .B2(G16), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT33), .B(G1976), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT94), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n780), .A2(new_n782), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n762), .A2(G6), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(new_n622), .B2(new_n762), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT32), .B(G1981), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT93), .ZN(new_n789));
  INV_X1    g364(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n787), .A2(new_n790), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n784), .A2(new_n785), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT34), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n774), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n794), .A2(KEYINPUT95), .A3(new_n795), .ZN(new_n797));
  INV_X1    g372(.A(KEYINPUT95), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n793), .B2(KEYINPUT34), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n796), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(KEYINPUT36), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT36), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n802), .B(new_n796), .C1(new_n797), .C2(new_n799), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(G105), .B1(new_n467), .B2(new_n468), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(KEYINPUT99), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT99), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n807), .B(G105), .C1(new_n467), .C2(new_n468), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n485), .A2(G129), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n483), .A2(G141), .ZN(new_n811));
  NAND3_X1  g386(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(KEYINPUT26), .Z(new_n813));
  NAND4_X1  g388(.A1(new_n809), .A2(new_n810), .A3(new_n811), .A4(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(G29), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(new_n816), .B2(G32), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT27), .B(G1996), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT100), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT101), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n816), .A2(G26), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(KEYINPUT28), .Z(new_n825));
  OAI21_X1  g400(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n826));
  INV_X1    g401(.A(G116), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(G2105), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n485), .B2(G128), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n483), .A2(G140), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n825), .B1(new_n831), .B2(G29), .ZN(new_n832));
  INV_X1    g407(.A(G2067), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n762), .A2(G20), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT23), .Z(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(G299), .B2(G16), .ZN(new_n837));
  INV_X1    g412(.A(G1956), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(G34), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n840), .A2(KEYINPUT24), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(KEYINPUT24), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n816), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(G160), .B2(new_n816), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G2084), .ZN(new_n845));
  NOR4_X1   g420(.A1(new_n823), .A2(new_n834), .A3(new_n839), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n762), .A2(G19), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT96), .Z(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n559), .B2(G16), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(G1341), .Z(new_n850));
  NAND2_X1  g425(.A1(new_n762), .A2(G21), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(G168), .B2(new_n762), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n852), .A2(G1966), .ZN(new_n853));
  XNOR2_X1  g428(.A(KEYINPUT31), .B(G11), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT30), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n816), .B1(new_n855), .B2(G28), .ZN(new_n856));
  AND2_X1   g431(.A1(new_n856), .A2(KEYINPUT102), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(G28), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n856), .B2(KEYINPUT102), .ZN(new_n859));
  OAI221_X1 g434(.A(new_n854), .B1(new_n857), .B2(new_n859), .C1(new_n666), .C2(new_n816), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n853), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(G29), .A2(G33), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(KEYINPUT97), .Z(new_n863));
  NAND3_X1  g438(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT98), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT25), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n483), .A2(G139), .ZN(new_n867));
  AOI22_X1  g442(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n868), .A2(new_n465), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n863), .B1(new_n870), .B2(new_n816), .ZN(new_n871));
  INV_X1    g446(.A(G2072), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(G27), .A2(G29), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(G164), .B2(G29), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n875), .A2(G2078), .ZN(new_n876));
  AOI22_X1  g451(.A1(new_n852), .A2(G1966), .B1(G2078), .B2(new_n875), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n861), .A2(new_n873), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  AOI211_X1 g453(.A(new_n850), .B(new_n878), .C1(new_n822), .C2(new_n821), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n816), .A2(G35), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT103), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n881), .B1(new_n489), .B2(G29), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT29), .ZN(new_n883));
  INV_X1    g458(.A(G2090), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n762), .A2(G5), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n886), .B1(G171), .B2(new_n762), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n887), .A2(G1961), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(G1961), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n885), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n645), .A2(G16), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n891), .B1(G4), .B2(G16), .ZN(new_n892));
  INV_X1    g467(.A(G1348), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(new_n872), .B2(new_n871), .ZN(new_n895));
  OAI22_X1  g470(.A1(new_n818), .A2(new_n820), .B1(new_n893), .B2(new_n892), .ZN(new_n896));
  AOI211_X1 g471(.A(new_n895), .B(new_n896), .C1(new_n884), .C2(new_n883), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n846), .A2(new_n879), .A3(new_n890), .A4(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT104), .B1(new_n804), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n901));
  AOI211_X1 g476(.A(new_n901), .B(new_n898), .C1(new_n801), .C2(new_n803), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n900), .A2(new_n902), .ZN(G311));
  NAND2_X1  g478(.A1(new_n804), .A2(new_n899), .ZN(G150));
  NAND2_X1  g479(.A1(new_n645), .A2(G559), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n905), .B(KEYINPUT38), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n556), .A2(new_n533), .A3(G93), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n907), .B1(new_n547), .B2(G55), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n524), .A2(new_n525), .A3(G67), .ZN(new_n909));
  NAND2_X1  g484(.A1(G80), .A2(G543), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(G651), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n559), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n555), .A2(new_n558), .A3(new_n908), .A4(new_n912), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n906), .B(new_n917), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n918), .A2(KEYINPUT39), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(KEYINPUT39), .ZN(new_n920));
  NOR3_X1   g495(.A1(new_n919), .A2(new_n920), .A3(G860), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n913), .A2(G860), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT37), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n921), .A2(new_n923), .ZN(G145));
  NAND2_X1  g499(.A1(new_n498), .A2(new_n500), .ZN(new_n925));
  INV_X1    g500(.A(new_n494), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n831), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(G164), .A2(new_n830), .A3(new_n829), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n928), .A2(new_n814), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n814), .B1(new_n928), .B2(new_n929), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n930), .A2(new_n931), .A3(new_n870), .ZN(new_n932));
  INV_X1    g507(.A(new_n870), .ZN(new_n933));
  INV_X1    g508(.A(new_n929), .ZN(new_n934));
  AOI21_X1  g509(.A(G164), .B1(new_n830), .B2(new_n829), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n815), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n928), .A2(new_n814), .A3(new_n929), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n932), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n483), .A2(G142), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n940), .B(KEYINPUT105), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n485), .A2(G130), .ZN(new_n942));
  OR2_X1    g517(.A1(G106), .A2(G2105), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n943), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n758), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n659), .ZN(new_n950));
  OAI211_X1 g525(.A(KEYINPUT106), .B(new_n753), .C1(new_n756), .C2(new_n757), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n950), .B1(new_n949), .B2(new_n951), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n947), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT108), .ZN(new_n956));
  INV_X1    g531(.A(new_n951), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n485), .A2(G119), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT91), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n755), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT106), .B1(new_n960), .B2(new_n753), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n659), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n962), .A2(new_n946), .A3(new_n952), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n939), .A2(new_n955), .A3(new_n956), .A4(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(G160), .B(new_n489), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n965), .B(new_n666), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n870), .B1(new_n930), .B2(new_n931), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n936), .A2(new_n933), .A3(new_n937), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n962), .A2(new_n946), .A3(new_n952), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n946), .B1(new_n962), .B2(new_n952), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n964), .A2(new_n966), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n939), .A2(new_n955), .A3(new_n963), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT108), .ZN(new_n975));
  AOI21_X1  g550(.A(G37), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT107), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n939), .A2(new_n955), .A3(KEYINPUT107), .A4(new_n963), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n979), .A3(new_n972), .ZN(new_n980));
  INV_X1    g555(.A(new_n966), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n976), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g559(.A1(new_n913), .A2(new_n632), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n654), .B(KEYINPUT86), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(new_n917), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT41), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n640), .A2(new_n641), .A3(new_n644), .ZN(new_n989));
  AND2_X1   g564(.A1(G299), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g565(.A1(G299), .A2(new_n989), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n581), .ZN(new_n993));
  AOI22_X1  g568(.A1(new_n993), .A2(new_n579), .B1(G651), .B2(new_n571), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n645), .A2(new_n576), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(G299), .A2(new_n989), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n995), .A2(KEYINPUT41), .A3(new_n996), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n992), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n987), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n990), .A2(new_n991), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n999), .B(new_n1000), .C1(new_n1002), .C2(new_n987), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1003), .B1(new_n1000), .B2(new_n999), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n770), .A2(new_n622), .ZN(new_n1005));
  NAND3_X1  g580(.A1(G290), .A2(new_n616), .A3(new_n621), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n584), .B1(new_n596), .B2(new_n600), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1008), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n596), .A2(new_n584), .A3(new_n600), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1012));
  AOI221_X4 g587(.A(new_n599), .B1(new_n510), .B2(new_n517), .C1(new_n593), .C2(new_n595), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1013), .A2(new_n1008), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1014), .A2(new_n1006), .A3(new_n1005), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT110), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1012), .A2(KEYINPUT110), .A3(new_n1015), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(KEYINPUT42), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1021), .B1(KEYINPUT42), .B2(new_n1016), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1004), .B(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n985), .B1(new_n1023), .B2(new_n632), .ZN(G295));
  OAI21_X1  g599(.A(new_n985), .B1(new_n1023), .B2(new_n632), .ZN(G331));
  INV_X1    g600(.A(KEYINPUT43), .ZN(new_n1026));
  AND4_X1   g601(.A1(new_n555), .A2(new_n558), .A3(new_n908), .A4(new_n912), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n555), .A2(new_n558), .B1(new_n908), .B2(new_n912), .ZN(new_n1028));
  NOR3_X1   g603(.A1(new_n527), .A2(KEYINPUT111), .A3(new_n536), .ZN(new_n1029));
  NOR3_X1   g604(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  OR3_X1    g605(.A1(new_n527), .A2(KEYINPUT111), .A3(new_n536), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1031), .B1(new_n914), .B2(new_n915), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT111), .B1(new_n527), .B2(new_n536), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT112), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n547), .A2(G52), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n508), .A2(new_n548), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1035), .B(new_n1036), .C1(new_n544), .C2(new_n545), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n544), .A2(new_n545), .ZN(new_n1038));
  OAI211_X1 g613(.A(new_n1033), .B(new_n1034), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1034), .B1(G301), .B2(new_n1033), .ZN(new_n1041));
  OAI22_X1  g616(.A1(new_n1030), .A2(new_n1032), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1029), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1033), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT112), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n914), .A2(new_n1031), .A3(new_n915), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1043), .A2(new_n1045), .A3(new_n1039), .A4(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1042), .A2(new_n1001), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT113), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT113), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1042), .A2(new_n1050), .A3(new_n1001), .A4(new_n1047), .ZN(new_n1051));
  AND4_X1   g626(.A1(new_n1045), .A2(new_n1043), .A3(new_n1039), .A4(new_n1046), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1046), .A2(new_n1043), .B1(new_n1045), .B2(new_n1039), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n998), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1049), .A2(new_n1051), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(G37), .B1(new_n1055), .B2(new_n1020), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1014), .A2(new_n1006), .A3(new_n1005), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1005), .A2(new_n1006), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1057), .A2(new_n1058), .A3(new_n1017), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT110), .B1(new_n1012), .B2(new_n1015), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1061), .A2(new_n1049), .A3(new_n1051), .A4(new_n1054), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1026), .B1(new_n1056), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1054), .A2(new_n1048), .ZN(new_n1064));
  AOI21_X1  g639(.A(G37), .B1(new_n1064), .B2(new_n1020), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1065), .A2(new_n1062), .A3(new_n1026), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n1063), .A2(new_n1066), .A3(KEYINPUT44), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1065), .A2(new_n1062), .A3(KEYINPUT114), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT43), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT114), .B1(new_n1065), .B2(new_n1062), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1068), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1065), .A2(new_n1062), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT114), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1075), .A2(KEYINPUT115), .A3(KEYINPUT43), .A4(new_n1069), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1056), .A2(new_n1026), .A3(new_n1062), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1072), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1067), .B1(new_n1078), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g654(.A1(G160), .A2(G40), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT116), .B(KEYINPUT45), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(G164), .B2(G1384), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G1986), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n770), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1086), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n770), .A2(new_n1085), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(KEYINPUT117), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(G1996), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n814), .B(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(new_n831), .B(new_n833), .ZN(new_n1094));
  INV_X1    g669(.A(new_n760), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n758), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n960), .A2(new_n760), .A3(new_n753), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1093), .A2(new_n1094), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  AOI22_X1  g673(.A1(new_n1088), .A2(new_n1091), .B1(new_n1083), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(G8), .ZN(new_n1100));
  INV_X1    g675(.A(G40), .ZN(new_n1101));
  AOI211_X1 g676(.A(new_n1101), .B(new_n466), .C1(new_n472), .C2(new_n474), .ZN(new_n1102));
  NOR2_X1   g677(.A1(G164), .A2(G1384), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1100), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n618), .A2(new_n610), .A3(new_n620), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1106), .A2(G1981), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT49), .ZN(new_n1108));
  NOR3_X1   g683(.A1(new_n613), .A2(new_n615), .A3(G1981), .ZN(new_n1109));
  OR3_X1    g684(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1108), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1110), .A2(new_n1104), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(G1976), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1112), .A2(new_n1113), .A3(new_n596), .A4(new_n600), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1109), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1105), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1117), .B(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(G2084), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT50), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1103), .A2(new_n1121), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1122), .A2(new_n1102), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1119), .A2(new_n1120), .A3(new_n1123), .ZN(new_n1124));
  OR3_X1    g699(.A1(G164), .A2(G1384), .A3(new_n1081), .ZN(new_n1125));
  OAI211_X1 g700(.A(new_n1125), .B(new_n1102), .C1(KEYINPUT45), .C2(new_n1103), .ZN(new_n1126));
  INV_X1    g701(.A(G1966), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g703(.A(new_n1100), .B(G286), .C1(new_n1124), .C2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(G288), .A2(new_n1113), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT52), .B1(new_n1105), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT52), .B1(G288), .B2(new_n1113), .ZN(new_n1132));
  OAI211_X1 g707(.A(new_n1104), .B(new_n1132), .C1(new_n1113), .C2(G288), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1131), .A2(new_n1112), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1119), .A2(new_n1123), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1103), .A2(KEYINPUT45), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1136), .A2(new_n1102), .A3(new_n1082), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  OAI22_X1  g713(.A1(new_n1135), .A2(G2090), .B1(G1971), .B2(new_n1138), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1139), .A2(G8), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n585), .A2(new_n586), .A3(G8), .ZN(new_n1141));
  XNOR2_X1  g716(.A(new_n1141), .B(KEYINPUT55), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1129), .B(new_n1134), .C1(new_n1140), .C2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1116), .B1(new_n1144), .B2(KEYINPUT63), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1139), .A2(G8), .A3(new_n1143), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1122), .A2(new_n1102), .A3(new_n1117), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1148), .A2(new_n884), .B1(new_n1137), .B2(new_n777), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1142), .B1(new_n1149), .B2(new_n1100), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1146), .A2(new_n1134), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1124), .A2(G168), .A3(new_n1128), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(G8), .ZN(new_n1153));
  AOI21_X1  g728(.A(G168), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT51), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT51), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1152), .A2(new_n1156), .A3(G8), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1151), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n1160));
  OR3_X1    g735(.A1(new_n1126), .A2(new_n1160), .A3(G2078), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1160), .B1(new_n1126), .B2(G2078), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1161), .A2(KEYINPUT53), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT53), .ZN(new_n1164));
  INV_X1    g739(.A(G2078), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1138), .A2(new_n1165), .ZN(new_n1166));
  XOR2_X1   g741(.A(KEYINPUT125), .B(G1961), .Z(new_n1167));
  AOI22_X1  g742(.A1(new_n1164), .A2(new_n1166), .B1(new_n1135), .B2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(G301), .B1(new_n1163), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1138), .A2(KEYINPUT53), .A3(new_n1165), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1164), .B1(new_n1137), .B2(G2078), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1122), .A2(new_n1102), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1172), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1167), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1170), .B(new_n1171), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1177), .A2(G171), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1159), .B1(new_n1169), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1159), .B1(new_n1177), .B2(G171), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1163), .A2(new_n1168), .A3(G301), .ZN(new_n1181));
  AOI21_X1  g756(.A(KEYINPUT126), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1180), .A2(new_n1181), .A3(KEYINPUT126), .ZN(new_n1183));
  OAI211_X1 g758(.A(new_n1158), .B(new_n1179), .C1(new_n1182), .C2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(G1348), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1186), .A2(G2067), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n645), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT119), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT57), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n994), .A2(new_n1189), .A3(new_n1190), .A4(new_n576), .ZN(new_n1191));
  NAND2_X1  g766(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1193));
  NAND3_X1  g768(.A1(G299), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1191), .A2(new_n1194), .ZN(new_n1195));
  AND2_X1   g770(.A1(new_n1147), .A2(new_n838), .ZN(new_n1196));
  XNOR2_X1  g771(.A(KEYINPUT56), .B(G2072), .ZN(new_n1197));
  XOR2_X1   g772(.A(new_n1197), .B(KEYINPUT120), .Z(new_n1198));
  INV_X1    g773(.A(new_n1198), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1137), .A2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1195), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1188), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1147), .A2(new_n838), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1195), .ZN(new_n1204));
  OAI211_X1 g779(.A(new_n1203), .B(new_n1204), .C1(new_n1137), .C2(new_n1199), .ZN(new_n1205));
  AND2_X1   g780(.A1(new_n1202), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g781(.A1(new_n1201), .A2(new_n1205), .A3(KEYINPUT61), .ZN(new_n1207));
  XOR2_X1   g782(.A(KEYINPUT58), .B(G1341), .Z(new_n1208));
  NAND2_X1  g783(.A1(new_n1186), .A2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g784(.A(new_n1209), .B1(new_n1137), .B2(G1996), .ZN(new_n1210));
  INV_X1    g785(.A(KEYINPUT121), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT59), .ZN(new_n1213));
  NOR2_X1   g788(.A1(new_n1213), .A2(KEYINPUT122), .ZN(new_n1214));
  OAI211_X1 g789(.A(new_n1209), .B(KEYINPUT121), .C1(G1996), .C2(new_n1137), .ZN(new_n1215));
  NAND4_X1  g790(.A1(new_n1212), .A2(new_n560), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  INV_X1    g791(.A(KEYINPUT60), .ZN(new_n1217));
  NAND2_X1  g792(.A1(new_n645), .A2(new_n1217), .ZN(new_n1218));
  OR3_X1    g793(.A1(new_n1185), .A2(new_n1187), .A3(new_n1218), .ZN(new_n1219));
  NAND3_X1  g794(.A1(new_n1207), .A2(new_n1216), .A3(new_n1219), .ZN(new_n1220));
  OAI221_X1 g795(.A(new_n989), .B1(G2067), .B2(new_n1186), .C1(new_n1175), .C2(G1348), .ZN(new_n1221));
  AOI21_X1  g796(.A(new_n1217), .B1(new_n1221), .B2(new_n1188), .ZN(new_n1222));
  XOR2_X1   g797(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1223));
  AOI21_X1  g798(.A(new_n559), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1223), .B1(new_n1224), .B2(new_n1215), .ZN(new_n1225));
  NOR3_X1   g800(.A1(new_n1220), .A2(new_n1222), .A3(new_n1225), .ZN(new_n1226));
  AOI21_X1  g801(.A(KEYINPUT61), .B1(new_n1201), .B2(new_n1205), .ZN(new_n1227));
  INV_X1    g802(.A(KEYINPUT123), .ZN(new_n1228));
  XNOR2_X1  g803(.A(new_n1227), .B(new_n1228), .ZN(new_n1229));
  AOI21_X1  g804(.A(new_n1206), .B1(new_n1226), .B2(new_n1229), .ZN(new_n1230));
  OAI21_X1  g805(.A(new_n1145), .B1(new_n1184), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1134), .A2(new_n1150), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1233), .A2(KEYINPUT62), .ZN(new_n1234));
  INV_X1    g809(.A(KEYINPUT62), .ZN(new_n1235));
  NAND3_X1  g810(.A1(new_n1155), .A2(new_n1235), .A3(new_n1157), .ZN(new_n1236));
  NAND3_X1  g811(.A1(new_n1234), .A2(new_n1169), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g812(.A(KEYINPUT63), .ZN(new_n1238));
  AOI22_X1  g813(.A1(new_n1140), .A2(new_n1143), .B1(new_n1129), .B2(new_n1238), .ZN(new_n1239));
  AOI21_X1  g814(.A(new_n1232), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g815(.A(new_n1099), .B1(new_n1231), .B2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g816(.A(new_n1084), .B1(new_n815), .B2(new_n1094), .ZN(new_n1242));
  INV_X1    g817(.A(KEYINPUT46), .ZN(new_n1243));
  NAND2_X1  g818(.A1(new_n1083), .A2(new_n1092), .ZN(new_n1244));
  AOI21_X1  g819(.A(new_n1242), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1245));
  OAI21_X1  g820(.A(new_n1245), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1246));
  XNOR2_X1  g821(.A(new_n1246), .B(KEYINPUT47), .ZN(new_n1247));
  NOR2_X1   g822(.A1(new_n1084), .A2(new_n1090), .ZN(new_n1248));
  OR2_X1    g823(.A1(new_n1248), .A2(KEYINPUT48), .ZN(new_n1249));
  NAND2_X1  g824(.A1(new_n1098), .A2(new_n1083), .ZN(new_n1250));
  NAND2_X1  g825(.A1(new_n1248), .A2(KEYINPUT48), .ZN(new_n1251));
  NAND3_X1  g826(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g827(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1253));
  OAI22_X1  g828(.A1(new_n1253), .A2(new_n1097), .B1(G2067), .B2(new_n831), .ZN(new_n1254));
  NAND2_X1  g829(.A1(new_n1254), .A2(new_n1083), .ZN(new_n1255));
  NAND3_X1  g830(.A1(new_n1247), .A2(new_n1252), .A3(new_n1255), .ZN(new_n1256));
  INV_X1    g831(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g832(.A1(new_n1241), .A2(new_n1257), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g833(.A1(new_n1056), .A2(new_n1062), .ZN(new_n1260));
  NAND2_X1  g834(.A1(new_n1260), .A2(KEYINPUT43), .ZN(new_n1261));
  INV_X1    g835(.A(new_n1066), .ZN(new_n1262));
  NAND2_X1  g836(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  OR2_X1    g837(.A1(G227), .A2(new_n460), .ZN(new_n1264));
  AOI21_X1  g838(.A(new_n1264), .B1(new_n741), .B2(new_n745), .ZN(new_n1265));
  NAND2_X1  g839(.A1(new_n697), .A2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g840(.A(new_n1266), .B1(new_n976), .B2(new_n982), .ZN(new_n1267));
  AOI21_X1  g841(.A(KEYINPUT127), .B1(new_n1263), .B2(new_n1267), .ZN(new_n1268));
  OAI211_X1 g842(.A(new_n1267), .B(KEYINPUT127), .C1(new_n1063), .C2(new_n1066), .ZN(new_n1269));
  INV_X1    g843(.A(new_n1269), .ZN(new_n1270));
  NOR2_X1   g844(.A1(new_n1268), .A2(new_n1270), .ZN(G308));
  OAI21_X1  g845(.A(new_n1267), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1272));
  INV_X1    g846(.A(KEYINPUT127), .ZN(new_n1273));
  NAND2_X1  g847(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g848(.A1(new_n1274), .A2(new_n1269), .ZN(G225));
endmodule


