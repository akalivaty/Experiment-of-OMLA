//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 0 1 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998;
  INV_X1    g000(.A(KEYINPUT10), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT64), .B1(new_n188), .B2(G143), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n188), .A2(G143), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(KEYINPUT1), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(new_n196), .A3(new_n195), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n191), .A2(G146), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT1), .ZN(new_n199));
  OAI21_X1  g013(.A(G128), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n191), .A2(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n195), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n187), .B1(new_n197), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G104), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT79), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT79), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G104), .ZN(new_n208));
  AOI21_X1  g022(.A(G107), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G104), .ZN(new_n211));
  OAI21_X1  g025(.A(G101), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT79), .B(G104), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT3), .B1(new_n213), .B2(G107), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(new_n210), .A3(G104), .ZN(new_n216));
  AOI21_X1  g030(.A(KEYINPUT80), .B1(new_n213), .B2(G107), .ZN(new_n217));
  AND4_X1   g031(.A1(KEYINPUT80), .A2(new_n206), .A3(new_n208), .A4(G107), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n214), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n204), .B(new_n212), .C1(new_n219), .C2(G101), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT82), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n206), .A2(new_n208), .A3(G107), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT80), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n213), .A2(KEYINPUT80), .A3(G107), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G101), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n227), .A2(new_n228), .A3(new_n214), .A4(new_n216), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n229), .A2(KEYINPUT82), .A3(new_n212), .A4(new_n204), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n222), .A2(new_n230), .ZN(new_n231));
  AND2_X1   g045(.A1(KEYINPUT81), .A2(G101), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n217), .A2(new_n218), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n216), .B1(new_n209), .B2(new_n215), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(KEYINPUT4), .A3(new_n229), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n198), .B1(new_n189), .B2(new_n192), .ZN(new_n237));
  NAND2_X1  g051(.A1(KEYINPUT0), .A2(G128), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n237), .A2(new_n239), .B1(new_n241), .B2(new_n202), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n219), .A2(KEYINPUT81), .A3(new_n243), .A4(G101), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n236), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G134), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n246), .A2(G137), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(G137), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n247), .B1(KEYINPUT11), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(KEYINPUT65), .A2(G137), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(KEYINPUT65), .A2(G137), .ZN(new_n252));
  NAND2_X1  g066(.A1(KEYINPUT11), .A2(G134), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(G131), .B1(new_n249), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G137), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT11), .B1(new_n256), .B2(G134), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n257), .B1(new_n246), .B2(G137), .ZN(new_n258));
  OR2_X1    g072(.A1(KEYINPUT65), .A2(G137), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n259), .A2(KEYINPUT11), .A3(G134), .A4(new_n250), .ZN(new_n260));
  INV_X1    g074(.A(G131), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n237), .B(new_n196), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n229), .A2(new_n212), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n187), .ZN(new_n267));
  NAND4_X1  g081(.A1(new_n231), .A2(new_n245), .A3(new_n264), .A4(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(G110), .B(G140), .ZN(new_n269));
  INV_X1    g083(.A(G227), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(G953), .ZN(new_n271));
  XOR2_X1   g085(.A(new_n269), .B(new_n271), .Z(new_n272));
  NAND2_X1  g086(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT83), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n231), .A2(new_n245), .A3(new_n267), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n263), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT83), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n268), .A2(new_n277), .A3(new_n272), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n274), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n229), .A2(new_n212), .A3(new_n265), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n197), .A2(new_n203), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n281), .B1(new_n229), .B2(new_n212), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n263), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT12), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI211_X1 g099(.A(KEYINPUT12), .B(new_n263), .C1(new_n280), .C2(new_n282), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(new_n268), .ZN(new_n288));
  INV_X1    g102(.A(new_n272), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n279), .A2(G469), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G469), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n287), .A2(new_n268), .A3(new_n272), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n272), .B1(new_n276), .B2(new_n268), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n292), .B(new_n293), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n292), .A2(new_n293), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n291), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT84), .ZN(new_n300));
  INV_X1    g114(.A(G221), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT9), .B(G234), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n301), .B1(new_n303), .B2(new_n293), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n299), .A2(new_n300), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n300), .B1(new_n299), .B2(new_n305), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G237), .ZN(new_n309));
  INV_X1    g123(.A(G953), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(new_n310), .A3(G214), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n311), .B(G143), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(new_n261), .ZN(new_n313));
  INV_X1    g127(.A(G125), .ZN(new_n314));
  NOR3_X1   g128(.A1(new_n314), .A2(KEYINPUT16), .A3(G140), .ZN(new_n315));
  INV_X1    g129(.A(G140), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n316), .B1(new_n317), .B2(new_n314), .ZN(new_n318));
  NAND3_X1  g132(.A1(KEYINPUT77), .A2(G125), .A3(G140), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n315), .B1(new_n320), .B2(KEYINPUT16), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G146), .ZN(new_n322));
  XNOR2_X1  g136(.A(G125), .B(G140), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n323), .A2(KEYINPUT19), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n324), .B1(KEYINPUT19), .B2(new_n320), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n313), .B(new_n322), .C1(G146), .C2(new_n325), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n312), .A2(new_n261), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(KEYINPUT18), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n188), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(new_n320), .B2(new_n188), .ZN(new_n330));
  INV_X1    g144(.A(new_n312), .ZN(new_n331));
  NAND2_X1  g145(.A1(KEYINPUT18), .A2(G131), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n332), .B(KEYINPUT88), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n328), .B(new_n330), .C1(new_n331), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n326), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(G113), .B(G122), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT89), .B(G104), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n336), .B(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n321), .B(new_n188), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n327), .A2(KEYINPUT17), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n340), .B(new_n341), .C1(new_n313), .C2(KEYINPUT17), .ZN(new_n342));
  INV_X1    g156(.A(new_n338), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(new_n334), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT20), .ZN(new_n346));
  INV_X1    g160(.A(G475), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .A4(new_n293), .ZN(new_n348));
  AOI211_X1 g162(.A(G475), .B(G902), .C1(new_n339), .C2(new_n344), .ZN(new_n349));
  XOR2_X1   g163(.A(KEYINPUT87), .B(KEYINPUT20), .Z(new_n350));
  OAI21_X1  g164(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n344), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n343), .B1(new_n342), .B2(new_n334), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n293), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT90), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(KEYINPUT90), .B(new_n293), .C1(new_n352), .C2(new_n353), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(G475), .A3(new_n357), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n194), .A2(G143), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n191), .A2(G128), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(new_n246), .ZN(new_n362));
  INV_X1    g176(.A(G122), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G116), .ZN(new_n364));
  INV_X1    g178(.A(G116), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G122), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n364), .A2(new_n366), .A3(new_n210), .ZN(new_n367));
  AOI21_X1  g181(.A(KEYINPUT14), .B1(new_n363), .B2(G116), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n368), .B1(new_n365), .B2(G122), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n366), .A2(KEYINPUT14), .ZN(new_n370));
  OAI21_X1  g184(.A(G107), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n362), .A2(new_n367), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n360), .B1(KEYINPUT13), .B2(new_n359), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n191), .A2(G128), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT13), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(KEYINPUT91), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT91), .B1(new_n374), .B2(new_n375), .ZN(new_n378));
  OAI21_X1  g192(.A(G134), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n364), .A2(new_n366), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G107), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n381), .A2(new_n367), .B1(new_n361), .B2(new_n246), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n379), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n372), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT74), .B(G217), .ZN(new_n385));
  OR3_X1    g199(.A1(new_n302), .A2(new_n385), .A3(G953), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n384), .B(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n293), .ZN(new_n388));
  INV_X1    g202(.A(G478), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n389), .A2(KEYINPUT15), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n388), .B(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(G952), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n393), .A2(G953), .ZN(new_n394));
  NAND2_X1  g208(.A1(G234), .A2(G237), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  XOR2_X1   g210(.A(KEYINPUT21), .B(G898), .Z(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(G902), .A3(G953), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AND4_X1   g213(.A1(new_n351), .A2(new_n358), .A3(new_n392), .A4(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(G214), .B1(G237), .B2(G902), .ZN(new_n401));
  XNOR2_X1  g215(.A(G110), .B(G122), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G119), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT66), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT66), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G119), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(new_n407), .A3(G116), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n365), .A2(G119), .ZN(new_n409));
  INV_X1    g223(.A(G113), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT2), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT2), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G113), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n408), .A2(new_n409), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT67), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n414), .B1(new_n408), .B2(new_n409), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n408), .A2(new_n409), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT67), .ZN(new_n420));
  INV_X1    g234(.A(new_n414), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n236), .A2(new_n244), .A3(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT85), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n236), .A2(new_n424), .A3(KEYINPUT85), .A4(new_n244), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n229), .A2(new_n212), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n408), .A2(KEYINPUT5), .A3(new_n409), .ZN(new_n430));
  OAI21_X1  g244(.A(G113), .B1(new_n408), .B2(KEYINPUT5), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n415), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n428), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n403), .B1(new_n427), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n425), .A2(new_n426), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n436), .A2(new_n428), .A3(new_n433), .A4(new_n402), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n435), .A2(KEYINPUT6), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n439), .B(new_n403), .C1(new_n427), .C2(new_n434), .ZN(new_n440));
  MUX2_X1   g254(.A(new_n242), .B(new_n281), .S(new_n314), .Z(new_n441));
  NAND2_X1  g255(.A1(new_n310), .A2(G224), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n441), .B(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n438), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G210), .B1(G237), .B2(G902), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT86), .B1(new_n310), .B2(G224), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n442), .A2(KEYINPUT7), .ZN(new_n447));
  OR3_X1    g261(.A1(new_n441), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n447), .B1(new_n441), .B2(new_n446), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n429), .B(new_n432), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n402), .B(KEYINPUT8), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(G902), .B1(new_n453), .B2(new_n437), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n444), .A2(new_n445), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n445), .B1(new_n444), .B2(new_n454), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n400), .B(new_n401), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(KEYINPUT92), .B1(new_n308), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n299), .A2(new_n305), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT84), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n299), .A2(new_n300), .A3(new_n305), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT92), .ZN(new_n463));
  INV_X1    g277(.A(new_n457), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  XNOR2_X1  g279(.A(KEYINPUT22), .B(G137), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n310), .A2(G221), .A3(G234), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n466), .B(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n322), .A2(new_n329), .ZN(new_n470));
  OR2_X1    g284(.A1(new_n194), .A2(KEYINPUT23), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n194), .A2(KEYINPUT23), .A3(G119), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(KEYINPUT66), .B(G119), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n194), .A2(KEYINPUT23), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G110), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(KEYINPUT78), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n474), .A2(new_n475), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n479), .A2(new_n477), .A3(new_n471), .A4(new_n472), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT78), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AND2_X1   g296(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  XOR2_X1   g297(.A(KEYINPUT24), .B(G110), .Z(new_n484));
  OR3_X1    g298(.A1(new_n404), .A2(KEYINPUT75), .A3(G128), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT75), .B1(new_n404), .B2(G128), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n405), .A2(new_n407), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n485), .B(new_n486), .C1(new_n487), .C2(new_n194), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT76), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n474), .A2(G128), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT76), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n486), .A4(new_n485), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n484), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n470), .B1(new_n483), .B2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n321), .B(G146), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n489), .A2(new_n492), .A3(new_n484), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n476), .A2(new_n477), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n469), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n478), .A2(new_n482), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n329), .B(new_n322), .C1(new_n501), .C2(new_n493), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n503), .A3(new_n468), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n385), .B1(G234), .B2(new_n293), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n506), .A2(G902), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT25), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n502), .A2(new_n503), .A3(new_n468), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n468), .B1(new_n502), .B2(new_n503), .ZN(new_n511));
  OAI211_X1 g325(.A(new_n509), .B(new_n293), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n506), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n509), .B1(new_n505), .B2(new_n293), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n508), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n309), .A2(new_n310), .A3(G210), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(KEYINPUT27), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT26), .B(G101), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n517), .B(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT68), .ZN(new_n520));
  AOI21_X1  g334(.A(G134), .B1(new_n259), .B2(new_n250), .ZN(new_n521));
  OAI21_X1  g335(.A(G131), .B1(new_n521), .B2(new_n247), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n522), .A2(new_n262), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n523), .A2(new_n281), .B1(new_n263), .B2(new_n242), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n419), .A2(new_n421), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(KEYINPUT67), .A3(new_n415), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n422), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n520), .B1(new_n524), .B2(new_n527), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n258), .A2(new_n261), .A3(new_n260), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n261), .B1(new_n258), .B2(new_n260), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n242), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n281), .A2(new_n262), .A3(new_n522), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n527), .A2(new_n520), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  OAI211_X1 g348(.A(KEYINPUT69), .B(new_n519), .C1(new_n528), .C2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n532), .A2(new_n531), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT30), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT30), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n532), .A2(new_n531), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n527), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n535), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n519), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT68), .B1(new_n536), .B2(new_n424), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n543), .B1(new_n544), .B2(new_n533), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(KEYINPUT69), .ZN(new_n546));
  OAI21_X1  g360(.A(KEYINPUT31), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n544), .A2(new_n533), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n536), .A2(new_n424), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(KEYINPUT28), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT71), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n536), .B(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT28), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n553), .A3(new_n527), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n550), .A2(new_n554), .A3(new_n543), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n547), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n540), .B1(new_n545), .B2(KEYINPUT69), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n519), .B1(new_n528), .B2(new_n534), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT69), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT70), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT31), .ZN(new_n562));
  NAND4_X1  g376(.A1(new_n557), .A2(new_n560), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n557), .A2(new_n560), .A3(new_n562), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT70), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n556), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(G472), .A2(G902), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT72), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT32), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n565), .A2(new_n563), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n557), .A2(new_n560), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n550), .A2(new_n554), .ZN(new_n573));
  AOI22_X1  g387(.A1(KEYINPUT31), .A2(new_n572), .B1(new_n573), .B2(new_n543), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT32), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n576), .A3(new_n568), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n570), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n543), .B1(new_n550), .B2(new_n554), .ZN(new_n579));
  AOI21_X1  g393(.A(G902), .B1(new_n579), .B2(KEYINPUT29), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT73), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n541), .A2(new_n548), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n543), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT29), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI22_X1  g399(.A1(new_n580), .A2(new_n581), .B1(new_n579), .B2(new_n585), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n580), .A2(new_n581), .ZN(new_n587));
  OAI21_X1  g401(.A(G472), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n515), .B1(new_n578), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n458), .A2(new_n465), .A3(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(G101), .ZN(G3));
  NAND2_X1  g405(.A1(new_n575), .A2(new_n568), .ZN(new_n592));
  INV_X1    g406(.A(G472), .ZN(new_n593));
  AOI21_X1  g407(.A(G902), .B1(new_n571), .B2(new_n574), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(new_n515), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n462), .ZN(new_n597));
  XOR2_X1   g411(.A(new_n597), .B(KEYINPUT93), .Z(new_n598));
  OAI211_X1 g412(.A(new_n399), .B(new_n401), .C1(new_n455), .C2(new_n456), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n387), .A2(new_n389), .A3(new_n293), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n387), .A2(KEYINPUT33), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n387), .A2(KEYINPUT33), .ZN(new_n603));
  AOI21_X1  g417(.A(G902), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n600), .B1(new_n604), .B2(new_n389), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n358), .A2(new_n351), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n599), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n598), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT94), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT95), .ZN(new_n612));
  XNOR2_X1  g426(.A(KEYINPUT34), .B(G104), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT96), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n612), .B(new_n614), .ZN(G6));
  INV_X1    g429(.A(new_n401), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n444), .A2(new_n454), .ZN(new_n617));
  INV_X1    g431(.A(new_n445), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n444), .A2(new_n445), .A3(new_n454), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n616), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT97), .ZN(new_n622));
  OR2_X1    g436(.A1(new_n358), .A2(new_n622), .ZN(new_n623));
  OR2_X1    g437(.A1(new_n349), .A2(new_n350), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n349), .A2(new_n350), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n392), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n358), .A2(new_n622), .ZN(new_n627));
  AND3_X1   g441(.A1(new_n623), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT98), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n621), .A2(new_n628), .A3(new_n629), .A4(new_n399), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n623), .A2(new_n626), .A3(new_n627), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT98), .B1(new_n599), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n598), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g448(.A(KEYINPUT35), .B(G107), .Z(new_n635));
  XNOR2_X1  g449(.A(new_n634), .B(new_n635), .ZN(G9));
  NAND2_X1  g450(.A1(new_n502), .A2(new_n503), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n468), .A2(KEYINPUT36), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n507), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n640), .B1(new_n513), .B2(new_n514), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI211_X1 g457(.A(KEYINPUT99), .B(new_n640), .C1(new_n513), .C2(new_n514), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n595), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n458), .A2(new_n465), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT37), .B(G110), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G12));
  AOI21_X1  g464(.A(new_n576), .B1(new_n575), .B2(new_n568), .ZN(new_n651));
  AOI211_X1 g465(.A(KEYINPUT32), .B(new_n569), .C1(new_n571), .C2(new_n574), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n588), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OR2_X1    g467(.A1(new_n398), .A2(G900), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n396), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n631), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n645), .B(new_n401), .C1(new_n456), .C2(new_n455), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n462), .A2(new_n653), .A3(new_n657), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n655), .B(KEYINPUT39), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n462), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n619), .A2(new_n620), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT38), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n519), .B1(new_n548), .B2(new_n549), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n557), .B2(new_n560), .ZN(new_n669));
  OAI21_X1  g483(.A(G472), .B1(new_n669), .B2(G902), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(new_n651), .B2(new_n652), .ZN(new_n671));
  INV_X1    g485(.A(new_n607), .ZN(new_n672));
  NOR4_X1   g486(.A1(new_n645), .A2(new_n672), .A3(new_n392), .A4(new_n616), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n667), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n662), .B1(new_n462), .B2(new_n663), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n665), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n191), .ZN(G45));
  NOR2_X1   g491(.A1(new_n608), .A2(new_n656), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n462), .A2(new_n653), .A3(new_n659), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G146), .ZN(G48));
  INV_X1    g494(.A(new_n515), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n293), .B1(new_n294), .B2(new_n295), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(G469), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(new_n305), .A3(new_n296), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n653), .A2(new_n609), .A3(new_n681), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT41), .B(G113), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G15));
  NAND3_X1  g502(.A1(new_n633), .A2(new_n589), .A3(new_n685), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G116), .ZN(G18));
  OAI21_X1  g504(.A(new_n401), .B1(new_n455), .B2(new_n456), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(new_n684), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n653), .A2(new_n692), .A3(new_n400), .A4(new_n645), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G119), .ZN(G21));
  AOI21_X1  g508(.A(new_n392), .B1(new_n358), .B2(new_n351), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n401), .B(new_n695), .C1(new_n455), .C2(new_n456), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n683), .A2(new_n305), .A3(new_n296), .A4(new_n399), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g512(.A(KEYINPUT100), .B1(new_n594), .B2(new_n593), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT100), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n700), .B(G472), .C1(new_n566), .C2(G902), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n698), .A2(new_n702), .A3(new_n592), .A4(new_n681), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G122), .ZN(G24));
  NOR2_X1   g518(.A1(new_n566), .A2(new_n569), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n705), .B1(new_n699), .B2(new_n701), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n706), .A2(new_n645), .A3(new_n678), .A4(new_n692), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G125), .ZN(G27));
  NAND3_X1  g522(.A1(new_n619), .A2(new_n401), .A3(new_n620), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT102), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n279), .A2(KEYINPUT101), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT101), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n274), .A2(new_n713), .A3(new_n276), .A4(new_n278), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n712), .A2(new_n290), .A3(new_n714), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n296), .B(new_n298), .C1(new_n715), .C2(new_n292), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n619), .A2(KEYINPUT102), .A3(new_n401), .A4(new_n620), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n711), .A2(new_n305), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n678), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(KEYINPUT42), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n719), .A2(new_n589), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n653), .A2(new_n681), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n723), .A2(new_n718), .A3(new_n720), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT42), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n722), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT103), .B(G131), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G33));
  NAND3_X1  g542(.A1(new_n719), .A2(new_n589), .A3(new_n657), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G134), .ZN(G36));
  NOR2_X1   g544(.A1(new_n607), .A2(new_n605), .ZN(new_n731));
  XOR2_X1   g545(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n607), .A2(new_n605), .A3(new_n736), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n734), .A2(new_n646), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n595), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n711), .A2(new_n717), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT106), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n711), .A2(new_n744), .A3(new_n717), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n738), .A2(KEYINPUT44), .A3(new_n595), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n741), .A2(new_n743), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n296), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n279), .A2(new_n290), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n292), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n712), .A2(KEYINPUT45), .A3(new_n290), .A4(new_n714), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n297), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n748), .B1(new_n753), .B2(KEYINPUT46), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n751), .A2(new_n752), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n298), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n304), .B1(new_n754), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT104), .B1(new_n759), .B2(new_n663), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n759), .A2(KEYINPUT104), .A3(new_n663), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n747), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n256), .ZN(G39));
  OR2_X1    g578(.A1(new_n759), .A2(KEYINPUT47), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n759), .A2(KEYINPUT47), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR4_X1   g581(.A1(new_n742), .A2(new_n653), .A3(new_n720), .A4(new_n681), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G140), .ZN(G42));
  NOR3_X1   g584(.A1(new_n734), .A2(new_n396), .A3(new_n737), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n706), .A2(new_n681), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n692), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n683), .A2(new_n296), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n742), .A2(new_n304), .A3(new_n775), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n671), .A2(new_n396), .A3(new_n515), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n774), .B(new_n394), .C1(new_n608), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n776), .A2(new_n771), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n780), .A2(KEYINPUT115), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(KEYINPUT115), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n589), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n783), .A2(KEYINPUT48), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(KEYINPUT48), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n779), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n743), .A2(new_n745), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n775), .A2(new_n305), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n787), .B(new_n773), .C1(new_n767), .C2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(KEYINPUT51), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n666), .A2(KEYINPUT38), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n666), .A2(KEYINPUT38), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n793), .A2(new_n616), .A3(new_n794), .A4(new_n685), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT114), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n797));
  OR3_X1    g611(.A1(new_n796), .A2(new_n797), .A3(new_n772), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n797), .B1(new_n796), .B2(new_n772), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AOI211_X1 g614(.A(new_n705), .B(new_n646), .C1(new_n699), .C2(new_n701), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n801), .B1(new_n781), .B2(new_n782), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n776), .A2(new_n672), .A3(new_n605), .A4(new_n777), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n800), .A2(new_n789), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n786), .B1(new_n792), .B2(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n804), .A2(new_n792), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n596), .A2(new_n462), .A3(new_n609), .ZN(new_n808));
  OR2_X1    g622(.A1(new_n607), .A2(new_n392), .ZN(new_n809));
  OR3_X1    g623(.A1(new_n599), .A2(KEYINPUT107), .A3(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(KEYINPUT107), .B1(new_n599), .B2(new_n809), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n810), .A2(new_n596), .A3(new_n462), .A4(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n590), .A2(new_n648), .A3(new_n808), .A4(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n624), .A2(new_n625), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n392), .A2(new_n655), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n627), .A2(new_n623), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n711), .A2(new_n717), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT108), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n646), .B1(new_n578), .B2(new_n588), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT108), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n711), .A2(new_n820), .A3(new_n816), .A4(new_n717), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n818), .A2(new_n462), .A3(new_n819), .A4(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n719), .A2(new_n678), .A3(new_n801), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(new_n729), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n813), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n689), .A2(new_n686), .A3(new_n693), .A4(new_n703), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n726), .A2(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n707), .A2(new_n660), .A3(new_n679), .ZN(new_n828));
  INV_X1    g642(.A(new_n696), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n655), .B(KEYINPUT109), .ZN(new_n830));
  OR3_X1    g644(.A1(new_n641), .A2(new_n304), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n671), .A2(new_n829), .A3(new_n716), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT110), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n831), .B1(new_n578), .B2(new_n670), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n836), .A2(KEYINPUT110), .A3(new_n829), .A4(new_n716), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT52), .B1(new_n828), .B2(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n828), .A2(new_n838), .A3(KEYINPUT52), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n825), .B(new_n827), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT112), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n844), .B1(new_n726), .B2(new_n826), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n719), .A2(new_n589), .A3(new_n678), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n723), .A2(new_n718), .ZN(new_n847));
  AOI22_X1  g661(.A1(new_n846), .A2(KEYINPUT42), .B1(new_n847), .B2(new_n721), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n633), .A2(new_n589), .A3(new_n685), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n686), .A2(new_n703), .A3(new_n693), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n848), .A2(new_n851), .A3(KEYINPUT112), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n845), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n828), .A2(new_n838), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT52), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n828), .A2(new_n838), .A3(KEYINPUT52), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n853), .A2(new_n858), .A3(KEYINPUT53), .A4(new_n825), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n843), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT113), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n843), .A2(new_n859), .A3(KEYINPUT113), .A4(new_n860), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT111), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n843), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n841), .A2(KEYINPUT111), .A3(new_n842), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n858), .A2(KEYINPUT53), .A3(new_n827), .A4(new_n825), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT54), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n807), .A2(new_n865), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n393), .A2(new_n310), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n775), .B(KEYINPUT49), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n731), .A2(new_n305), .A3(new_n401), .A4(new_n681), .ZN(new_n876));
  OR4_X1    g690(.A1(new_n667), .A2(new_n671), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n874), .A2(new_n877), .ZN(G75));
  INV_X1    g692(.A(KEYINPUT56), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n843), .A2(new_n859), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(G902), .ZN(new_n881));
  INV_X1    g695(.A(G210), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n438), .A2(new_n440), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(new_n443), .ZN(new_n885));
  XOR2_X1   g699(.A(new_n885), .B(KEYINPUT55), .Z(new_n886));
  AND2_X1   g700(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n883), .A2(new_n886), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n310), .A2(G952), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(G51));
  NAND4_X1  g704(.A1(new_n880), .A2(G902), .A3(new_n752), .A4(new_n751), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT117), .ZN(new_n892));
  INV_X1    g706(.A(new_n861), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n860), .B1(new_n843), .B2(new_n859), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n297), .B(KEYINPUT57), .Z(new_n896));
  OAI22_X1  g710(.A1(new_n895), .A2(new_n896), .B1(new_n295), .B2(new_n294), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n889), .B1(new_n892), .B2(new_n897), .ZN(G54));
  INV_X1    g712(.A(KEYINPUT58), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n881), .A2(new_n899), .A3(new_n347), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n900), .A2(new_n345), .ZN(new_n901));
  INV_X1    g715(.A(new_n889), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n902), .B1(new_n900), .B2(new_n345), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n901), .A2(new_n903), .ZN(G60));
  NAND2_X1  g718(.A1(G478), .A2(G902), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT59), .ZN(new_n906));
  INV_X1    g720(.A(new_n603), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n906), .B1(new_n907), .B2(new_n601), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n902), .B1(new_n895), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n865), .A2(new_n871), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n906), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n907), .A2(new_n601), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(G63));
  NAND2_X1  g727(.A1(G217), .A2(G902), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT118), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT60), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n880), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n505), .B(KEYINPUT119), .Z(new_n918));
  AOI21_X1  g732(.A(new_n889), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n639), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n919), .B1(new_n920), .B2(new_n917), .ZN(new_n921));
  XOR2_X1   g735(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n922), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n919), .B(new_n924), .C1(new_n920), .C2(new_n917), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n923), .A2(new_n925), .ZN(G66));
  NOR2_X1   g740(.A1(new_n813), .A2(new_n826), .ZN(new_n927));
  AND2_X1   g741(.A1(G224), .A2(G953), .ZN(new_n928));
  AOI22_X1  g742(.A1(new_n927), .A2(new_n310), .B1(new_n397), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n884), .B1(G898), .B2(new_n310), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(G69));
  INV_X1    g745(.A(G900), .ZN(new_n932));
  OAI21_X1  g746(.A(G953), .B1(new_n270), .B2(new_n932), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT124), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT127), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n537), .A2(new_n539), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT121), .Z(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(new_n325), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n707), .A2(new_n660), .A3(new_n679), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(KEYINPUT125), .B1(new_n941), .B2(new_n763), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n828), .A2(new_n940), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n939), .A2(KEYINPUT122), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n741), .A2(new_n746), .ZN(new_n946));
  INV_X1    g760(.A(new_n762), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n787), .B(new_n946), .C1(new_n947), .C2(new_n760), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT125), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n945), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n942), .A2(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n589), .B(new_n829), .C1(new_n947), .C2(new_n760), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n952), .A2(new_n769), .A3(new_n848), .A4(new_n729), .ZN(new_n953));
  INV_X1    g767(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g768(.A(G953), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n310), .A2(G900), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n935), .B(new_n938), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n938), .ZN(new_n958));
  INV_X1    g772(.A(new_n676), .ZN(new_n959));
  AOI21_X1  g773(.A(KEYINPUT62), .B1(new_n945), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n961));
  AOI211_X1 g775(.A(new_n961), .B(new_n676), .C1(new_n943), .C2(new_n944), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n769), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n809), .A2(new_n608), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n589), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n462), .A2(new_n663), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n965), .A2(new_n966), .A3(new_n742), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n763), .A2(KEYINPUT123), .A3(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT123), .ZN(new_n969));
  INV_X1    g783(.A(new_n967), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n969), .B1(new_n948), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n968), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n963), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n958), .B1(new_n973), .B2(G953), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n957), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n956), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n953), .B1(new_n942), .B2(new_n950), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n976), .B1(new_n977), .B2(G953), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n935), .B1(new_n978), .B2(new_n938), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n934), .B1(new_n975), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n938), .ZN(new_n981));
  INV_X1    g795(.A(new_n934), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n981), .A2(new_n974), .A3(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT126), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n981), .A2(new_n974), .A3(KEYINPUT126), .A4(new_n982), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n980), .A2(new_n985), .A3(new_n986), .ZN(G72));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT63), .Z(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n990), .B1(new_n973), .B2(new_n927), .ZN(new_n991));
  INV_X1    g805(.A(new_n582), .ZN(new_n992));
  NOR3_X1   g806(.A1(new_n991), .A2(new_n543), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n990), .B1(new_n977), .B2(new_n927), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n992), .A2(new_n543), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n902), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(new_n990), .B1(new_n572), .B2(new_n583), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n870), .A2(new_n997), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n993), .A2(new_n996), .A3(new_n998), .ZN(G57));
endmodule


