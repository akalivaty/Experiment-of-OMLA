

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U322 ( .A(n348), .B(G148GAT), .ZN(n349) );
  XNOR2_X1 U323 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U324 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n408) );
  XNOR2_X1 U325 ( .A(n409), .B(n408), .ZN(n526) );
  NOR2_X1 U326 ( .A1(n515), .A2(n424), .ZN(n565) );
  XOR2_X1 U327 ( .A(n459), .B(KEYINPUT28), .Z(n530) );
  XNOR2_X1 U328 ( .A(n443), .B(KEYINPUT58), .ZN(n444) );
  XNOR2_X1 U329 ( .A(n445), .B(n444), .ZN(G1351GAT) );
  XOR2_X1 U330 ( .A(KEYINPUT67), .B(G162GAT), .Z(n291) );
  XNOR2_X1 U331 ( .A(G190GAT), .B(G134GAT), .ZN(n290) );
  XNOR2_X1 U332 ( .A(n291), .B(n290), .ZN(n301) );
  XOR2_X1 U333 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n299) );
  INV_X1 U334 ( .A(KEYINPUT7), .ZN(n295) );
  XOR2_X1 U335 ( .A(KEYINPUT8), .B(G50GAT), .Z(n293) );
  XNOR2_X1 U336 ( .A(G43GAT), .B(G36GAT), .ZN(n292) );
  XNOR2_X1 U337 ( .A(n293), .B(n292), .ZN(n294) );
  XNOR2_X1 U338 ( .A(n295), .B(n294), .ZN(n367) );
  XOR2_X1 U339 ( .A(G92GAT), .B(KEYINPUT75), .Z(n297) );
  XNOR2_X1 U340 ( .A(G99GAT), .B(G85GAT), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n297), .B(n296), .ZN(n347) );
  XNOR2_X1 U342 ( .A(n367), .B(n347), .ZN(n298) );
  XNOR2_X1 U343 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U344 ( .A(n301), .B(n300), .ZN(n309) );
  NAND2_X1 U345 ( .A1(G232GAT), .A2(G233GAT), .ZN(n307) );
  XOR2_X1 U346 ( .A(KEYINPUT10), .B(KEYINPUT66), .Z(n303) );
  XNOR2_X1 U347 ( .A(G29GAT), .B(KEYINPUT80), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n303), .B(n302), .ZN(n305) );
  XOR2_X1 U349 ( .A(G106GAT), .B(G218GAT), .Z(n304) );
  XNOR2_X1 U350 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U351 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U352 ( .A(n309), .B(n308), .ZN(n556) );
  XOR2_X1 U353 ( .A(KEYINPUT2), .B(G162GAT), .Z(n311) );
  XNOR2_X1 U354 ( .A(G155GAT), .B(G148GAT), .ZN(n310) );
  XNOR2_X1 U355 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U356 ( .A(KEYINPUT3), .B(n312), .Z(n333) );
  XOR2_X1 U357 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n314) );
  XNOR2_X1 U358 ( .A(G50GAT), .B(KEYINPUT23), .ZN(n313) );
  XNOR2_X1 U359 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U360 ( .A(n333), .B(n315), .ZN(n325) );
  XOR2_X1 U361 ( .A(G22GAT), .B(KEYINPUT89), .Z(n317) );
  NAND2_X1 U362 ( .A1(G228GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U363 ( .A(n317), .B(n316), .ZN(n320) );
  XOR2_X1 U364 ( .A(G211GAT), .B(KEYINPUT21), .Z(n319) );
  XNOR2_X1 U365 ( .A(G197GAT), .B(G218GAT), .ZN(n318) );
  XNOR2_X1 U366 ( .A(n319), .B(n318), .ZN(n413) );
  XOR2_X1 U367 ( .A(n320), .B(n413), .Z(n323) );
  XNOR2_X1 U368 ( .A(G106GAT), .B(G78GAT), .ZN(n321) );
  XNOR2_X1 U369 ( .A(n321), .B(G204GAT), .ZN(n358) );
  XNOR2_X1 U370 ( .A(G141GAT), .B(n358), .ZN(n322) );
  XNOR2_X1 U371 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U372 ( .A(n325), .B(n324), .ZN(n459) );
  XOR2_X1 U373 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n327) );
  XNOR2_X1 U374 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n326) );
  XNOR2_X1 U375 ( .A(n327), .B(n326), .ZN(n342) );
  XOR2_X1 U376 ( .A(G120GAT), .B(G57GAT), .Z(n343) );
  XOR2_X1 U377 ( .A(KEYINPUT90), .B(KEYINPUT5), .Z(n329) );
  XNOR2_X1 U378 ( .A(G85GAT), .B(KEYINPUT4), .ZN(n328) );
  XNOR2_X1 U379 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U380 ( .A(n343), .B(n330), .Z(n332) );
  NAND2_X1 U381 ( .A1(G225GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U382 ( .A(n332), .B(n331), .ZN(n334) );
  XOR2_X1 U383 ( .A(n334), .B(n333), .Z(n340) );
  XOR2_X1 U384 ( .A(G1GAT), .B(G113GAT), .Z(n336) );
  XNOR2_X1 U385 ( .A(G29GAT), .B(G141GAT), .ZN(n335) );
  XNOR2_X1 U386 ( .A(n336), .B(n335), .ZN(n368) );
  XOR2_X1 U387 ( .A(G127GAT), .B(KEYINPUT85), .Z(n338) );
  XNOR2_X1 U388 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n337) );
  XNOR2_X1 U389 ( .A(n338), .B(n337), .ZN(n428) );
  XNOR2_X1 U390 ( .A(n368), .B(n428), .ZN(n339) );
  XNOR2_X1 U391 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U392 ( .A(n342), .B(n341), .ZN(n466) );
  XNOR2_X1 U393 ( .A(KEYINPUT93), .B(n466), .ZN(n515) );
  XOR2_X1 U394 ( .A(KEYINPUT32), .B(KEYINPUT76), .Z(n345) );
  XOR2_X1 U395 ( .A(G176GAT), .B(G64GAT), .Z(n416) );
  XNOR2_X1 U396 ( .A(n343), .B(n416), .ZN(n344) );
  XNOR2_X1 U397 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U398 ( .A(n346), .B(KEYINPUT31), .Z(n352) );
  XOR2_X1 U399 ( .A(n347), .B(KEYINPUT78), .Z(n350) );
  NAND2_X1 U400 ( .A1(G230GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U401 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U402 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n354) );
  XNOR2_X1 U403 ( .A(KEYINPUT77), .B(KEYINPUT74), .ZN(n353) );
  XNOR2_X1 U404 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U405 ( .A(n356), .B(n355), .ZN(n360) );
  XNOR2_X1 U406 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n357) );
  XNOR2_X1 U407 ( .A(n357), .B(KEYINPUT72), .ZN(n384) );
  XOR2_X1 U408 ( .A(n358), .B(n384), .Z(n359) );
  XNOR2_X1 U409 ( .A(n360), .B(n359), .ZN(n570) );
  OR2_X1 U410 ( .A1(n570), .A2(KEYINPUT65), .ZN(n362) );
  NAND2_X1 U411 ( .A1(n570), .A2(KEYINPUT65), .ZN(n361) );
  NAND2_X1 U412 ( .A1(n362), .A2(n361), .ZN(n363) );
  XNOR2_X1 U413 ( .A(n363), .B(KEYINPUT41), .ZN(n502) );
  XOR2_X1 U414 ( .A(KEYINPUT70), .B(KEYINPUT68), .Z(n365) );
  XNOR2_X1 U415 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n364) );
  XNOR2_X1 U416 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U417 ( .A(n367), .B(n366), .ZN(n375) );
  XOR2_X1 U418 ( .A(G22GAT), .B(G15GAT), .Z(n381) );
  XOR2_X1 U419 ( .A(n368), .B(n381), .Z(n370) );
  NAND2_X1 U420 ( .A1(G229GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U421 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U422 ( .A(n371), .B(KEYINPUT69), .Z(n373) );
  XOR2_X1 U423 ( .A(G169GAT), .B(G8GAT), .Z(n418) );
  XNOR2_X1 U424 ( .A(G197GAT), .B(n418), .ZN(n372) );
  XNOR2_X1 U425 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U426 ( .A(n375), .B(n374), .Z(n566) );
  NOR2_X1 U427 ( .A1(n502), .A2(n566), .ZN(n377) );
  INV_X1 U428 ( .A(KEYINPUT46), .ZN(n376) );
  XNOR2_X1 U429 ( .A(n377), .B(n376), .ZN(n399) );
  INV_X1 U430 ( .A(n556), .ZN(n397) );
  XOR2_X1 U431 ( .A(G57GAT), .B(G211GAT), .Z(n379) );
  XNOR2_X1 U432 ( .A(G127GAT), .B(G78GAT), .ZN(n378) );
  XNOR2_X1 U433 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U434 ( .A(n380), .B(G155GAT), .Z(n383) );
  XNOR2_X1 U435 ( .A(n381), .B(G183GAT), .ZN(n382) );
  XNOR2_X1 U436 ( .A(n383), .B(n382), .ZN(n388) );
  XOR2_X1 U437 ( .A(n384), .B(KEYINPUT81), .Z(n386) );
  NAND2_X1 U438 ( .A1(G231GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U439 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U440 ( .A(n388), .B(n387), .Z(n396) );
  XOR2_X1 U441 ( .A(KEYINPUT15), .B(G64GAT), .Z(n390) );
  XNOR2_X1 U442 ( .A(G8GAT), .B(G1GAT), .ZN(n389) );
  XNOR2_X1 U443 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U444 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n392) );
  XNOR2_X1 U445 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n391) );
  XNOR2_X1 U446 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U447 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U448 ( .A(n396), .B(n395), .ZN(n538) );
  NOR2_X1 U449 ( .A1(n397), .A2(n538), .ZN(n398) );
  NAND2_X1 U450 ( .A1(n399), .A2(n398), .ZN(n401) );
  XOR2_X1 U451 ( .A(KEYINPUT113), .B(KEYINPUT47), .Z(n400) );
  XNOR2_X1 U452 ( .A(n401), .B(n400), .ZN(n407) );
  XNOR2_X1 U453 ( .A(n566), .B(KEYINPUT71), .ZN(n531) );
  XNOR2_X1 U454 ( .A(n397), .B(KEYINPUT36), .ZN(n577) );
  NAND2_X1 U455 ( .A1(n577), .A2(n538), .ZN(n402) );
  XOR2_X1 U456 ( .A(KEYINPUT114), .B(n402), .Z(n403) );
  XNOR2_X1 U457 ( .A(KEYINPUT45), .B(n403), .ZN(n404) );
  NAND2_X1 U458 ( .A1(n570), .A2(n404), .ZN(n405) );
  NOR2_X1 U459 ( .A1(n531), .A2(n405), .ZN(n406) );
  NOR2_X1 U460 ( .A1(n407), .A2(n406), .ZN(n409) );
  XOR2_X1 U461 ( .A(KEYINPUT18), .B(G190GAT), .Z(n411) );
  XNOR2_X1 U462 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n410) );
  XNOR2_X1 U463 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U464 ( .A(KEYINPUT17), .B(n412), .Z(n429) );
  XNOR2_X1 U465 ( .A(n429), .B(n413), .ZN(n422) );
  XOR2_X1 U466 ( .A(G92GAT), .B(G204GAT), .Z(n415) );
  NAND2_X1 U467 ( .A1(G226GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U468 ( .A(n415), .B(n414), .ZN(n417) );
  XOR2_X1 U469 ( .A(n417), .B(n416), .Z(n420) );
  XNOR2_X1 U470 ( .A(G36GAT), .B(n418), .ZN(n419) );
  XNOR2_X1 U471 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U472 ( .A(n422), .B(n421), .ZN(n453) );
  NOR2_X1 U473 ( .A1(n526), .A2(n453), .ZN(n423) );
  XOR2_X1 U474 ( .A(KEYINPUT54), .B(n423), .Z(n424) );
  NAND2_X1 U475 ( .A1(n459), .A2(n565), .ZN(n425) );
  XNOR2_X1 U476 ( .A(n425), .B(KEYINPUT55), .ZN(n442) );
  XOR2_X1 U477 ( .A(G120GAT), .B(G176GAT), .Z(n427) );
  XNOR2_X1 U478 ( .A(G169GAT), .B(KEYINPUT87), .ZN(n426) );
  XNOR2_X1 U479 ( .A(n427), .B(n426), .ZN(n433) );
  XOR2_X1 U480 ( .A(G71GAT), .B(n428), .Z(n431) );
  XNOR2_X1 U481 ( .A(G113GAT), .B(n429), .ZN(n430) );
  XNOR2_X1 U482 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U483 ( .A(n433), .B(n432), .ZN(n441) );
  NAND2_X1 U484 ( .A1(G227GAT), .A2(G233GAT), .ZN(n439) );
  XOR2_X1 U485 ( .A(KEYINPUT88), .B(KEYINPUT20), .Z(n435) );
  XNOR2_X1 U486 ( .A(G15GAT), .B(KEYINPUT86), .ZN(n434) );
  XNOR2_X1 U487 ( .A(n435), .B(n434), .ZN(n437) );
  XOR2_X1 U488 ( .A(G43GAT), .B(G99GAT), .Z(n436) );
  XNOR2_X1 U489 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U490 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X2 U491 ( .A(n441), .B(n440), .ZN(n527) );
  NAND2_X1 U492 ( .A1(n442), .A2(n527), .ZN(n562) );
  NOR2_X1 U493 ( .A1(n556), .A2(n562), .ZN(n445) );
  INV_X1 U494 ( .A(G190GAT), .ZN(n443) );
  INV_X1 U495 ( .A(n531), .ZN(n446) );
  NOR2_X1 U496 ( .A1(n446), .A2(n562), .ZN(n449) );
  XNOR2_X1 U497 ( .A(KEYINPUT123), .B(KEYINPUT124), .ZN(n447) );
  XNOR2_X1 U498 ( .A(n447), .B(G169GAT), .ZN(n448) );
  XNOR2_X1 U499 ( .A(n449), .B(n448), .ZN(G1348GAT) );
  XOR2_X1 U500 ( .A(KEYINPUT99), .B(KEYINPUT34), .Z(n474) );
  NAND2_X1 U501 ( .A1(n570), .A2(n531), .ZN(n450) );
  XOR2_X1 U502 ( .A(KEYINPUT79), .B(n450), .Z(n486) );
  XOR2_X1 U503 ( .A(KEYINPUT84), .B(KEYINPUT16), .Z(n452) );
  NAND2_X1 U504 ( .A1(n538), .A2(n556), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(n472) );
  INV_X1 U506 ( .A(n453), .ZN(n518) );
  XNOR2_X1 U507 ( .A(n518), .B(KEYINPUT27), .ZN(n462) );
  NAND2_X1 U508 ( .A1(n515), .A2(n462), .ZN(n525) );
  NOR2_X1 U509 ( .A1(n530), .A2(n525), .ZN(n454) );
  XOR2_X1 U510 ( .A(KEYINPUT94), .B(n454), .Z(n455) );
  NOR2_X1 U511 ( .A1(n527), .A2(n455), .ZN(n470) );
  NAND2_X1 U512 ( .A1(n527), .A2(n518), .ZN(n456) );
  NAND2_X1 U513 ( .A1(n456), .A2(n459), .ZN(n457) );
  XNOR2_X1 U514 ( .A(n457), .B(KEYINPUT96), .ZN(n458) );
  XNOR2_X1 U515 ( .A(n458), .B(KEYINPUT25), .ZN(n464) );
  NOR2_X1 U516 ( .A1(n459), .A2(n527), .ZN(n461) );
  XNOR2_X1 U517 ( .A(KEYINPUT95), .B(KEYINPUT26), .ZN(n460) );
  XOR2_X1 U518 ( .A(n461), .B(n460), .Z(n564) );
  AND2_X1 U519 ( .A1(n462), .A2(n564), .ZN(n463) );
  NOR2_X1 U520 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U521 ( .A(n465), .B(KEYINPUT97), .ZN(n467) );
  NAND2_X1 U522 ( .A1(n467), .A2(n466), .ZN(n468) );
  XOR2_X1 U523 ( .A(KEYINPUT98), .B(n468), .Z(n469) );
  NOR2_X1 U524 ( .A1(n470), .A2(n469), .ZN(n484) );
  INV_X1 U525 ( .A(n484), .ZN(n471) );
  NAND2_X1 U526 ( .A1(n472), .A2(n471), .ZN(n503) );
  NOR2_X1 U527 ( .A1(n486), .A2(n503), .ZN(n479) );
  NAND2_X1 U528 ( .A1(n479), .A2(n515), .ZN(n473) );
  XNOR2_X1 U529 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U530 ( .A(G1GAT), .B(n475), .ZN(G1324GAT) );
  NAND2_X1 U531 ( .A1(n518), .A2(n479), .ZN(n476) );
  XNOR2_X1 U532 ( .A(n476), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U533 ( .A(G15GAT), .B(KEYINPUT35), .Z(n478) );
  NAND2_X1 U534 ( .A1(n479), .A2(n527), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n481) );
  NAND2_X1 U537 ( .A1(n479), .A2(n530), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U539 ( .A(G22GAT), .B(n482), .ZN(G1327GAT) );
  XOR2_X1 U540 ( .A(G29GAT), .B(KEYINPUT39), .Z(n490) );
  INV_X1 U541 ( .A(n538), .ZN(n574) );
  NAND2_X1 U542 ( .A1(n574), .A2(n577), .ZN(n483) );
  NOR2_X1 U543 ( .A1(n484), .A2(n483), .ZN(n485) );
  XNOR2_X1 U544 ( .A(KEYINPUT37), .B(n485), .ZN(n514) );
  NOR2_X1 U545 ( .A1(n514), .A2(n486), .ZN(n488) );
  XOR2_X1 U546 ( .A(KEYINPUT103), .B(KEYINPUT38), .Z(n487) );
  XNOR2_X1 U547 ( .A(n488), .B(n487), .ZN(n499) );
  NAND2_X1 U548 ( .A1(n515), .A2(n499), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U550 ( .A(n491), .B(KEYINPUT105), .Z(n493) );
  XNOR2_X1 U551 ( .A(KEYINPUT102), .B(KEYINPUT104), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  NAND2_X1 U553 ( .A1(n499), .A2(n518), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n494), .B(G36GAT), .ZN(G1329GAT) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(KEYINPUT106), .ZN(n498) );
  XOR2_X1 U556 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n496) );
  NAND2_X1 U557 ( .A1(n499), .A2(n527), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(G1330GAT) );
  NAND2_X1 U560 ( .A1(n499), .A2(n530), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n500), .B(KEYINPUT108), .ZN(n501) );
  XNOR2_X1 U562 ( .A(G50GAT), .B(n501), .ZN(G1331GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT109), .B(KEYINPUT42), .Z(n505) );
  INV_X1 U564 ( .A(n502), .ZN(n548) );
  NAND2_X1 U565 ( .A1(n566), .A2(n548), .ZN(n513) );
  NOR2_X1 U566 ( .A1(n513), .A2(n503), .ZN(n509) );
  NAND2_X1 U567 ( .A1(n509), .A2(n515), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NAND2_X1 U570 ( .A1(n518), .A2(n509), .ZN(n507) );
  XNOR2_X1 U571 ( .A(n507), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U572 ( .A1(n527), .A2(n509), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n508), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U575 ( .A1(n509), .A2(n530), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U577 ( .A(G78GAT), .B(n512), .ZN(G1335GAT) );
  XOR2_X1 U578 ( .A(G85GAT), .B(KEYINPUT111), .Z(n517) );
  NOR2_X1 U579 ( .A1(n514), .A2(n513), .ZN(n522) );
  NAND2_X1 U580 ( .A1(n522), .A2(n515), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(G1336GAT) );
  NAND2_X1 U582 ( .A1(n518), .A2(n522), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n519), .B(KEYINPUT112), .ZN(n520) );
  XNOR2_X1 U584 ( .A(G92GAT), .B(n520), .ZN(G1337GAT) );
  NAND2_X1 U585 ( .A1(n527), .A2(n522), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n521), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U587 ( .A1(n522), .A2(n530), .ZN(n523) );
  XNOR2_X1 U588 ( .A(n523), .B(KEYINPUT44), .ZN(n524) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  XNOR2_X1 U590 ( .A(G113GAT), .B(KEYINPUT116), .ZN(n533) );
  NOR2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n546) );
  NAND2_X1 U592 ( .A1(n546), .A2(n527), .ZN(n528) );
  XOR2_X1 U593 ( .A(KEYINPUT115), .B(n528), .Z(n529) );
  NOR2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n543) );
  NAND2_X1 U595 ( .A1(n531), .A2(n543), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT117), .Z(n535) );
  NAND2_X1 U598 ( .A1(n543), .A2(n548), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(n537) );
  XOR2_X1 U600 ( .A(KEYINPUT49), .B(KEYINPUT118), .Z(n536) );
  XNOR2_X1 U601 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(KEYINPUT120), .ZN(n542) );
  XOR2_X1 U603 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n540) );
  NAND2_X1 U604 ( .A1(n543), .A2(n538), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n542), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U607 ( .A(G134GAT), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U608 ( .A1(n543), .A2(n397), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  NAND2_X1 U610 ( .A1(n546), .A2(n564), .ZN(n555) );
  NOR2_X1 U611 ( .A1(n566), .A2(n555), .ZN(n547) );
  XOR2_X1 U612 ( .A(G141GAT), .B(n547), .Z(G1344GAT) );
  NOR2_X1 U613 ( .A1(n502), .A2(n555), .ZN(n553) );
  XOR2_X1 U614 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n550) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(KEYINPUT121), .B(n551), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  NOR2_X1 U619 ( .A1(n574), .A2(n555), .ZN(n554) );
  XOR2_X1 U620 ( .A(G155GAT), .B(n554), .Z(G1346GAT) );
  NOR2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U622 ( .A(G162GAT), .B(n557), .Z(G1347GAT) );
  NOR2_X1 U623 ( .A1(n562), .A2(n502), .ZN(n561) );
  XOR2_X1 U624 ( .A(KEYINPUT57), .B(KEYINPUT125), .Z(n559) );
  XNOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1349GAT) );
  NOR2_X1 U628 ( .A1(n574), .A2(n562), .ZN(n563) );
  XOR2_X1 U629 ( .A(G183GAT), .B(n563), .Z(G1350GAT) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n576) );
  NOR2_X1 U631 ( .A1(n566), .A2(n576), .ZN(n568) );
  XNOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  NOR2_X1 U635 ( .A1(n570), .A2(n576), .ZN(n572) );
  XNOR2_X1 U636 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G204GAT), .B(n573), .ZN(G1353GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n576), .ZN(n575) );
  XOR2_X1 U640 ( .A(G211GAT), .B(n575), .Z(G1354GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n580) );
  INV_X1 U642 ( .A(n576), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

