//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 1 0 0 0 0 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT70), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT11), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G137), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT11), .A3(G134), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(G137), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G131), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n191), .A2(new_n193), .A3(new_n197), .A4(new_n194), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n199));
  AND2_X1   g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n198), .A2(new_n199), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n196), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g018(.A(new_n198), .B(new_n199), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT67), .A3(new_n196), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT0), .A2(G128), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n208), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n208), .A2(new_n210), .ZN(new_n213));
  XOR2_X1   g027(.A(KEYINPUT0), .B(G128), .Z(new_n214));
  OAI21_X1  g028(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n204), .A2(new_n206), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT1), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n208), .A2(new_n210), .A3(new_n217), .A4(G128), .ZN(new_n218));
  INV_X1    g032(.A(G128), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G128), .ZN(new_n222));
  AOI22_X1  g036(.A1(new_n220), .A2(new_n222), .B1(new_n208), .B2(KEYINPUT1), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n218), .B1(new_n223), .B2(new_n213), .ZN(new_n224));
  INV_X1    g038(.A(new_n194), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n190), .A2(G137), .ZN(new_n226));
  OAI21_X1  g040(.A(G131), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n205), .A2(new_n224), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n216), .A2(KEYINPUT30), .A3(new_n228), .ZN(new_n229));
  XOR2_X1   g043(.A(KEYINPUT2), .B(G113), .Z(new_n230));
  XNOR2_X1  g044(.A(G116), .B(G119), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(KEYINPUT66), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT2), .B(G113), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT66), .ZN(new_n234));
  INV_X1    g048(.A(G116), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n235), .A2(G119), .ZN(new_n236));
  AND2_X1   g050(.A1(new_n235), .A2(G119), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n233), .B(new_n234), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n232), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n202), .A2(new_n215), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n228), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT30), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n240), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n229), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(G237), .A2(G953), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G210), .ZN(new_n247));
  XOR2_X1   g061(.A(new_n247), .B(KEYINPUT27), .Z(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(G101), .ZN(new_n249));
  XOR2_X1   g063(.A(new_n248), .B(new_n249), .Z(new_n250));
  AND2_X1   g064(.A1(new_n224), .A2(new_n227), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n239), .B1(new_n251), .B2(new_n205), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT68), .B1(new_n216), .B2(new_n252), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n216), .A2(new_n252), .A3(KEYINPUT68), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n245), .B(new_n250), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT31), .ZN(new_n256));
  INV_X1    g070(.A(new_n253), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n216), .A2(new_n252), .A3(KEYINPUT68), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT31), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n259), .A2(new_n260), .A3(new_n250), .A4(new_n245), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n256), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n242), .ZN(new_n263));
  OAI22_X1  g077(.A1(new_n254), .A2(new_n253), .B1(new_n240), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(KEYINPUT28), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n216), .A2(new_n228), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT69), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n216), .A2(KEYINPUT69), .A3(new_n228), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n240), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT28), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n250), .B1(new_n265), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n188), .B1(new_n262), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT32), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT32), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n276), .B(new_n188), .C1(new_n262), .C2(new_n273), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n265), .A2(new_n272), .A3(new_n250), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT29), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n259), .A2(new_n245), .ZN(new_n281));
  INV_X1    g095(.A(new_n250), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n279), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n266), .A2(new_n239), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(new_n254), .B2(new_n253), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT28), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n282), .A2(new_n280), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n287), .A2(new_n272), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT71), .ZN(new_n290));
  INV_X1    g104(.A(G902), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n287), .A2(new_n272), .A3(new_n292), .A4(new_n288), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n284), .A2(new_n290), .A3(new_n291), .A4(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G472), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n278), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(G110), .B(G140), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n297), .B(KEYINPUT77), .ZN(new_n298));
  INV_X1    g112(.A(G953), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G227), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n298), .B(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G104), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT3), .B1(new_n302), .B2(G107), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT3), .ZN(new_n304));
  INV_X1    g118(.A(G107), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(G104), .ZN(new_n306));
  INV_X1    g120(.A(G101), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n302), .A2(G107), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n303), .A2(new_n306), .A3(new_n307), .A4(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n302), .A2(G107), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n305), .A2(G104), .ZN(new_n311));
  OAI21_X1  g125(.A(G101), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n313), .A2(G128), .B1(new_n208), .B2(new_n210), .ZN(new_n314));
  INV_X1    g128(.A(new_n218), .ZN(new_n315));
  OAI211_X1 g129(.A(new_n309), .B(new_n312), .C1(new_n314), .C2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n309), .A2(new_n312), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n316), .B1(new_n224), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(KEYINPUT12), .A3(new_n202), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n204), .A2(new_n206), .A3(new_n319), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT12), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n321), .A2(KEYINPUT80), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT80), .B1(new_n321), .B2(new_n322), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n320), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT78), .B(KEYINPUT10), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n316), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT79), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n327), .B(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n204), .A2(new_n206), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n303), .A2(new_n306), .A3(new_n308), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT4), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n332), .A3(G101), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n331), .A2(G101), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n309), .A2(KEYINPUT4), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n215), .B(new_n333), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n318), .A2(KEYINPUT10), .A3(new_n224), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n329), .A2(new_n330), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n301), .B1(new_n325), .B2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n327), .B(KEYINPUT79), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n204), .A2(new_n206), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n342), .A2(new_n343), .A3(new_n338), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n330), .B1(new_n329), .B2(new_n339), .ZN(new_n345));
  INV_X1    g159(.A(new_n301), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n344), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n291), .B1(new_n341), .B2(new_n347), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n344), .A2(new_n346), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n325), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n343), .B1(new_n342), .B2(new_n338), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n301), .B1(new_n351), .B2(new_n340), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(G902), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  XOR2_X1   g168(.A(KEYINPUT81), .B(G469), .Z(new_n355));
  AOI22_X1  g169(.A1(new_n348), .A2(G469), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT91), .B1(new_n235), .B2(G122), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT91), .ZN(new_n358));
  INV_X1    g172(.A(G122), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(G116), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n235), .A2(G122), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n305), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(KEYINPUT14), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n361), .B(new_n362), .C1(KEYINPUT14), .C2(new_n305), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n220), .A2(new_n222), .A3(G143), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n209), .A2(G128), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n190), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n190), .B1(new_n367), .B2(new_n368), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n365), .B(new_n366), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT13), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n368), .A2(new_n373), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n367), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n374), .B1(new_n376), .B2(KEYINPUT92), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT92), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n367), .A2(new_n378), .A3(new_n375), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n190), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n361), .A2(new_n305), .A3(new_n362), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n369), .B1(new_n381), .B2(new_n363), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n372), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(KEYINPUT9), .B(G234), .ZN(new_n384));
  INV_X1    g198(.A(G217), .ZN(new_n385));
  NOR3_X1   g199(.A1(new_n384), .A2(new_n385), .A3(G953), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n372), .B(new_n386), .C1(new_n380), .C2(new_n382), .ZN(new_n389));
  AOI21_X1  g203(.A(G902), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G478), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n392), .A2(KEYINPUT15), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT93), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n390), .B(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n394), .B1(new_n396), .B2(new_n393), .ZN(new_n397));
  INV_X1    g211(.A(G237), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(new_n299), .A3(G214), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n209), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n246), .A2(G143), .A3(G214), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G131), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT86), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT17), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT86), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n402), .A2(new_n406), .A3(G131), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n400), .A2(new_n197), .A3(new_n401), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n404), .A2(new_n405), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G140), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G125), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n411), .A2(KEYINPUT16), .ZN(new_n412));
  INV_X1    g226(.A(G125), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G140), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n411), .A2(new_n414), .A3(KEYINPUT16), .ZN(new_n415));
  AOI21_X1  g229(.A(G146), .B1(new_n412), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n412), .A2(G146), .A3(new_n415), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n406), .B1(new_n402), .B2(G131), .ZN(new_n421));
  AOI211_X1 g235(.A(KEYINPUT86), .B(new_n197), .C1(new_n400), .C2(new_n401), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT17), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n409), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n411), .A2(new_n414), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(KEYINPUT85), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n411), .A2(new_n414), .A3(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(G146), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n425), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n207), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(KEYINPUT18), .A2(G131), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n400), .A2(new_n401), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n402), .A2(KEYINPUT18), .A3(G131), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  XNOR2_X1  g250(.A(G113), .B(G122), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT88), .B(G104), .ZN(new_n438));
  XNOR2_X1  g252(.A(new_n437), .B(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n424), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n436), .ZN(new_n441));
  INV_X1    g255(.A(new_n418), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n421), .A2(new_n422), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n442), .B1(new_n443), .B2(new_n408), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n426), .A2(KEYINPUT19), .A3(new_n428), .ZN(new_n445));
  OR2_X1    g259(.A1(new_n425), .A2(KEYINPUT19), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n207), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT87), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n445), .A2(KEYINPUT87), .A3(new_n207), .A4(new_n446), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n441), .B1(new_n444), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n440), .B1(new_n452), .B2(new_n439), .ZN(new_n453));
  NOR2_X1   g267(.A1(G475), .A2(G902), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n454), .A2(KEYINPUT89), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n454), .A2(KEYINPUT89), .ZN(new_n456));
  NOR3_X1   g270(.A1(new_n455), .A2(new_n456), .A3(KEYINPUT20), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT90), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n453), .A2(new_n454), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT20), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n453), .A2(KEYINPUT90), .A3(new_n457), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(new_n440), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n439), .B1(new_n424), .B2(new_n436), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n291), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G475), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n299), .A2(G952), .ZN(new_n469));
  INV_X1    g283(.A(G234), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n469), .B1(new_n470), .B2(new_n398), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(G902), .B(G953), .C1(new_n470), .C2(new_n398), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n473), .B(KEYINPUT94), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT21), .B(G898), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n397), .A2(new_n464), .A3(new_n468), .A4(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(G221), .B1(new_n384), .B2(G902), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(G214), .B1(G237), .B2(G902), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n239), .B(new_n333), .C1(new_n334), .C2(new_n335), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n230), .A2(new_n231), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n483), .A2(new_n309), .A3(new_n312), .ZN(new_n484));
  OR2_X1    g298(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n485));
  NAND2_X1  g299(.A1(KEYINPUT82), .A2(KEYINPUT5), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n236), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT83), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(new_n486), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n231), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT83), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n236), .A2(new_n485), .A3(new_n491), .A4(new_n486), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n488), .A2(G113), .A3(new_n490), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n484), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(G110), .B(G122), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n482), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  OAI211_X1 g310(.A(G125), .B(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n299), .A2(G224), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n498), .A2(KEYINPUT7), .ZN(new_n499));
  OAI221_X1 g313(.A(new_n497), .B1(KEYINPUT84), .B2(new_n499), .C1(new_n224), .C2(G125), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n499), .B1(new_n497), .B2(KEYINPUT84), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n497), .B1(new_n224), .B2(G125), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n496), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  XOR2_X1   g318(.A(new_n495), .B(KEYINPUT8), .Z(new_n505));
  NAND2_X1  g319(.A1(new_n493), .A2(new_n483), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(new_n317), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n231), .A2(KEYINPUT5), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n488), .A2(G113), .A3(new_n492), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n484), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n505), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(G902), .B1(new_n504), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n482), .A2(new_n494), .ZN(new_n514));
  INV_X1    g328(.A(new_n495), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(KEYINPUT6), .A3(new_n496), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT6), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n514), .A2(new_n518), .A3(new_n515), .ZN(new_n519));
  XOR2_X1   g333(.A(new_n502), .B(new_n498), .Z(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(G210), .B1(G237), .B2(G902), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n513), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n522), .B1(new_n513), .B2(new_n521), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n481), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR4_X1   g339(.A1(new_n356), .A2(new_n478), .A3(new_n480), .A4(new_n525), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT22), .B(G137), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n299), .A2(G221), .A3(G234), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XOR2_X1   g343(.A(new_n529), .B(KEYINPUT73), .Z(new_n530));
  NAND2_X1  g344(.A1(new_n418), .A2(new_n431), .ZN(new_n531));
  AOI21_X1  g345(.A(KEYINPUT23), .B1(new_n219), .B2(G119), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n219), .A2(G119), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT65), .B(G128), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(KEYINPUT23), .A3(G119), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT72), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT72), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n536), .A2(new_n539), .A3(KEYINPUT23), .A4(G119), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n535), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G110), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n536), .A2(G119), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n544), .B1(G119), .B2(new_n219), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT24), .B(G110), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n531), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n538), .A2(new_n540), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n542), .B1(new_n549), .B2(new_n534), .ZN(new_n550));
  OAI22_X1  g364(.A1(new_n442), .A2(new_n416), .B1(new_n545), .B2(new_n546), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n530), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g367(.A1(new_n541), .A2(new_n542), .B1(new_n545), .B2(new_n546), .ZN(new_n554));
  OAI221_X1 g368(.A(new_n529), .B1(new_n550), .B2(new_n551), .C1(new_n554), .C2(new_n531), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n385), .B1(G234), .B2(new_n291), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(G902), .ZN(new_n558));
  XOR2_X1   g372(.A(KEYINPUT74), .B(KEYINPUT75), .Z(new_n559));
  XNOR2_X1  g373(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n556), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT76), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n553), .A2(new_n555), .A3(new_n291), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT25), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n553), .A2(new_n555), .A3(KEYINPUT25), .A4(new_n291), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n568), .A2(new_n557), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n563), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n296), .A2(new_n526), .A3(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(G101), .ZN(G3));
  INV_X1    g386(.A(KEYINPUT95), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n525), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n522), .ZN(new_n575));
  AND3_X1   g389(.A1(new_n517), .A2(new_n519), .A3(new_n520), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n496), .A2(new_n500), .A3(new_n503), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n291), .B1(new_n577), .B2(new_n511), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n575), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n513), .A2(new_n521), .A3(new_n522), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(KEYINPUT95), .A3(new_n481), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n574), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n391), .A2(new_n395), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n390), .A2(KEYINPUT93), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n392), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT33), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n388), .A2(new_n587), .A3(new_n389), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n587), .B1(new_n388), .B2(new_n389), .ZN(new_n589));
  OAI211_X1 g403(.A(G478), .B(new_n291), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  AOI22_X1  g404(.A1(new_n464), .A2(new_n468), .B1(new_n586), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n583), .A2(new_n477), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT96), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT96), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n583), .A2(new_n594), .A3(new_n477), .A4(new_n591), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n291), .B1(new_n262), .B2(new_n273), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(G472), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n598), .A2(new_n274), .ZN(new_n599));
  OR2_X1    g413(.A1(new_n563), .A2(new_n569), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n600), .A2(new_n356), .A3(new_n480), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n596), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT97), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT34), .B(G104), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G6));
  NOR2_X1   g419(.A1(new_n461), .A2(KEYINPUT20), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT20), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n607), .B1(new_n453), .B2(new_n454), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n468), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n397), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n583), .A2(new_n477), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(new_n599), .A3(new_n601), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G107), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT98), .B(KEYINPUT35), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G9));
  NOR2_X1   g430(.A1(new_n548), .A2(new_n552), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n530), .A2(KEYINPUT36), .ZN(new_n618));
  XOR2_X1   g432(.A(new_n617), .B(new_n618), .Z(new_n619));
  AOI22_X1  g433(.A1(new_n568), .A2(new_n557), .B1(new_n619), .B2(new_n560), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n478), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n356), .A2(new_n480), .ZN(new_n622));
  INV_X1    g436(.A(new_n525), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n599), .A2(new_n621), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT37), .B(G110), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G12));
  INV_X1    g440(.A(new_n620), .ZN(new_n627));
  INV_X1    g441(.A(G900), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n474), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n471), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n468), .B(new_n630), .C1(new_n606), .C2(new_n608), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n397), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n583), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n348), .A2(G469), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n354), .A2(new_n355), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n479), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT99), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n638), .A2(new_n296), .A3(new_n639), .ZN(new_n640));
  AOI22_X1  g454(.A1(new_n275), .A2(new_n277), .B1(new_n294), .B2(G472), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n620), .B1(new_n574), .B2(new_n582), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n642), .A2(new_n479), .A3(new_n636), .A4(new_n632), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT99), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G128), .ZN(G30));
  XOR2_X1   g460(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n630), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n622), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT40), .ZN(new_n650));
  AOI21_X1  g464(.A(G902), .B1(new_n281), .B2(new_n250), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n651), .B1(new_n250), .B2(new_n286), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(G472), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n278), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n620), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n464), .A2(new_n468), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(new_n397), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n581), .B(KEYINPUT38), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n657), .A2(new_n481), .A3(new_n658), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n650), .A2(new_n655), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT101), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G143), .ZN(G45));
  AOI21_X1  g476(.A(new_n637), .B1(new_n278), .B2(new_n295), .ZN(new_n663));
  INV_X1    g477(.A(new_n630), .ZN(new_n664));
  AOI221_X4 g478(.A(new_n664), .B1(new_n586), .B2(new_n590), .C1(new_n464), .C2(new_n468), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n642), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G146), .ZN(G48));
  AOI21_X1  g482(.A(new_n600), .B1(new_n278), .B2(new_n295), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n352), .B1(new_n325), .B2(new_n349), .ZN(new_n671));
  OAI21_X1  g485(.A(G469), .B1(new_n671), .B2(G902), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n635), .A2(new_n672), .A3(new_n479), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n596), .ZN(new_n675));
  XNOR2_X1  g489(.A(KEYINPUT41), .B(G113), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G15));
  NAND2_X1  g491(.A1(new_n674), .A2(new_n612), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G116), .ZN(G18));
  AOI21_X1  g493(.A(new_n673), .B1(new_n574), .B2(new_n582), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n296), .A2(new_n680), .A3(new_n681), .A4(new_n621), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n635), .A2(new_n672), .A3(new_n479), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n621), .A2(new_n683), .A3(new_n583), .ZN(new_n684));
  OAI21_X1  g498(.A(KEYINPUT102), .B1(new_n641), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G119), .ZN(G21));
  XOR2_X1   g501(.A(new_n188), .B(KEYINPUT103), .Z(new_n688));
  AOI21_X1  g502(.A(new_n250), .B1(new_n287), .B2(new_n272), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n688), .B1(new_n262), .B2(new_n689), .ZN(new_n690));
  AND2_X1   g504(.A1(new_n256), .A2(new_n261), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n265), .A2(new_n272), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n282), .ZN(new_n693));
  AOI21_X1  g507(.A(G902), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT104), .B(G472), .Z(new_n695));
  OAI211_X1 g509(.A(new_n570), .B(new_n690), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n695), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n597), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(KEYINPUT105), .A3(new_n570), .A4(new_n690), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n657), .A2(new_n583), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n703), .A2(new_n476), .A3(new_n673), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  AND4_X1   g520(.A1(new_n627), .A2(new_n700), .A3(new_n665), .A4(new_n690), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n680), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G125), .ZN(G27));
  INV_X1    g523(.A(new_n581), .ZN(new_n710));
  INV_X1    g524(.A(new_n481), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n480), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n710), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n341), .A2(new_n347), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n714), .A2(new_n715), .A3(G469), .A4(new_n291), .ZN(new_n716));
  INV_X1    g530(.A(G469), .ZN(new_n717));
  INV_X1    g531(.A(new_n320), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n321), .A2(new_n322), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT80), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n321), .A2(KEYINPUT80), .A3(new_n322), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n718), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n346), .B1(new_n723), .B2(new_n344), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n349), .A2(new_n351), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n717), .B1(new_n726), .B2(new_n291), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n716), .B1(new_n727), .B2(new_n715), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n713), .B1(new_n728), .B2(new_n635), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n296), .A2(new_n729), .A3(new_n570), .A4(new_n665), .ZN(new_n730));
  NOR2_X1   g544(.A1(KEYINPUT107), .A2(KEYINPUT42), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n731), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n669), .A2(new_n665), .A3(new_n729), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G131), .ZN(G33));
  NAND4_X1  g550(.A1(new_n296), .A2(new_n729), .A3(new_n570), .A4(new_n632), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G134), .ZN(G36));
  OR2_X1    g552(.A1(new_n714), .A2(KEYINPUT45), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n714), .A2(KEYINPUT45), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(G469), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(G469), .A2(G902), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT46), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n741), .A2(KEYINPUT46), .A3(new_n742), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n635), .A3(new_n746), .ZN(new_n747));
  AND2_X1   g561(.A1(new_n747), .A2(new_n479), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n648), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT108), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n748), .A2(new_n751), .A3(new_n648), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT43), .B1(new_n656), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n586), .A2(new_n590), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n656), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n755), .B(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n599), .A2(new_n620), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n759), .A3(KEYINPUT44), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n581), .A2(new_n711), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT44), .B1(new_n758), .B2(new_n759), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n753), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G137), .ZN(G39));
  AND4_X1   g580(.A1(new_n641), .A2(new_n600), .A3(new_n665), .A4(new_n761), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n748), .A2(KEYINPUT47), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n748), .A2(KEYINPUT47), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT110), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n748), .B(KEYINPUT47), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT110), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n773), .A3(new_n767), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G140), .ZN(G42));
  XOR2_X1   g590(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n777));
  AOI22_X1  g591(.A1(new_n682), .A2(new_n685), .B1(new_n702), .B2(new_n704), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n669), .B(new_n683), .C1(new_n596), .C2(new_n612), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n735), .A2(new_n778), .A3(KEYINPUT53), .A4(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n761), .ZN(new_n781));
  INV_X1    g595(.A(new_n397), .ZN(new_n782));
  NOR4_X1   g596(.A1(new_n781), .A2(new_n782), .A3(new_n620), .A4(new_n631), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n663), .A2(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n737), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n782), .A2(new_n464), .A3(KEYINPUT112), .A4(new_n468), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT112), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n464), .A2(new_n468), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n787), .B1(new_n788), .B2(new_n397), .ZN(new_n789));
  INV_X1    g603(.A(new_n591), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n786), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n525), .A2(new_n476), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n599), .A2(new_n601), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n571), .A2(new_n793), .A3(new_n624), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n728), .A2(new_n635), .ZN(new_n796));
  INV_X1    g610(.A(new_n713), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n700), .A2(new_n665), .A3(new_n627), .A4(new_n690), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n707), .A2(KEYINPUT113), .A3(new_n729), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n785), .A2(new_n794), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(new_n780), .B1(KEYINPUT117), .B2(new_n803), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n803), .A2(KEYINPUT117), .ZN(new_n805));
  AOI22_X1  g619(.A1(new_n663), .A2(new_n666), .B1(new_n707), .B2(new_n680), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n703), .A2(new_n480), .A3(new_n664), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n807), .A2(new_n654), .A3(new_n620), .A4(new_n796), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n645), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n645), .A2(new_n806), .A3(new_n808), .A4(KEYINPUT52), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n811), .A2(KEYINPUT114), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT114), .B1(new_n811), .B2(new_n812), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n804), .B(new_n805), .C1(new_n813), .C2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT116), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n735), .A2(new_n779), .A3(new_n778), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n803), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n811), .A2(new_n812), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n816), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n821), .ZN(new_n823));
  AOI211_X1 g637(.A(KEYINPUT116), .B(new_n823), .C1(new_n818), .C2(new_n819), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n777), .B(new_n815), .C1(new_n822), .C2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n813), .A2(new_n814), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n779), .A2(new_n686), .A3(new_n705), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n737), .A2(new_n784), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n571), .A2(new_n793), .A3(new_n624), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n828), .A2(new_n735), .A3(new_n802), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n827), .A2(new_n832), .ZN(new_n833));
  OAI22_X1  g647(.A1(new_n833), .A2(KEYINPUT53), .B1(new_n820), .B2(new_n821), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n826), .B1(KEYINPUT54), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n758), .A2(new_n472), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n702), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n837), .A2(new_n481), .A3(new_n658), .A4(new_n673), .ZN(new_n838));
  XNOR2_X1  g652(.A(new_n838), .B(KEYINPUT50), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n673), .A2(new_n781), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n570), .A3(new_n472), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n841), .A2(new_n654), .ZN(new_n842));
  OR3_X1    g656(.A1(new_n842), .A2(new_n788), .A3(new_n756), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n700), .A2(new_n627), .A3(new_n690), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n836), .A2(new_n840), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT120), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n839), .B(new_n843), .C1(new_n844), .C2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT51), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n836), .A2(new_n702), .A3(new_n761), .ZN(new_n849));
  INV_X1    g663(.A(new_n772), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n635), .A2(new_n672), .A3(new_n480), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n849), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OR3_X1    g666(.A1(new_n847), .A2(new_n848), .A3(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n851), .B(KEYINPUT119), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n849), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n848), .B1(new_n847), .B2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n680), .ZN(new_n857));
  OAI221_X1 g671(.A(new_n469), .B1(new_n790), .B2(new_n842), .C1(new_n837), .C2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n846), .A2(new_n670), .ZN(new_n859));
  INV_X1    g673(.A(new_n859), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n860), .A2(KEYINPUT48), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(KEYINPUT48), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n858), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n835), .A2(new_n853), .A3(new_n856), .A4(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(G952), .B2(G953), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n570), .A2(new_n712), .ZN(new_n866));
  OR3_X1    g680(.A1(new_n866), .A2(new_n757), .A3(new_n658), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n635), .A2(new_n672), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n868), .A2(KEYINPUT49), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(KEYINPUT49), .ZN(new_n870));
  NOR4_X1   g684(.A1(new_n867), .A2(new_n654), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT111), .Z(new_n872));
  NAND2_X1  g686(.A1(new_n865), .A2(new_n872), .ZN(G75));
  INV_X1    g687(.A(KEYINPUT56), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n815), .B1(new_n822), .B2(new_n824), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(G902), .ZN(new_n876));
  INV_X1    g690(.A(G210), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n517), .A2(new_n519), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(new_n520), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT55), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n878), .A2(new_n881), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n299), .A2(G952), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(G51));
  INV_X1    g699(.A(new_n671), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n811), .A2(new_n812), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n821), .B1(new_n887), .B2(new_n832), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT116), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n820), .A2(new_n816), .A3(new_n821), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n777), .B1(new_n891), .B2(new_n815), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n892), .A2(new_n826), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n742), .B(KEYINPUT57), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n886), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n876), .A2(new_n741), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n884), .B1(new_n895), .B2(new_n896), .ZN(G54));
  NAND4_X1  g711(.A1(new_n875), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n898));
  INV_X1    g712(.A(new_n453), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n898), .A2(new_n899), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n900), .A2(new_n901), .A3(new_n884), .ZN(G60));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT121), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n588), .A2(new_n589), .ZN(new_n905));
  NAND2_X1  g719(.A1(G478), .A2(G902), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT59), .Z(new_n907));
  NOR2_X1   g721(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  OAI211_X1 g722(.A(new_n904), .B(new_n908), .C1(new_n892), .C2(new_n826), .ZN(new_n909));
  INV_X1    g723(.A(new_n884), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n777), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n875), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n825), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n904), .B1(new_n914), .B2(new_n908), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n903), .B1(new_n911), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n908), .B1(new_n892), .B2(new_n826), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT121), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n918), .A2(KEYINPUT122), .A3(new_n910), .A4(new_n909), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n905), .B1(new_n835), .B2(new_n907), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(G63));
  NAND2_X1  g735(.A1(G217), .A2(G902), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT123), .Z(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n891), .B2(new_n815), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n910), .B1(new_n925), .B2(new_n556), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n619), .B2(new_n925), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT61), .ZN(G66));
  INV_X1    g742(.A(new_n475), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n299), .B1(new_n929), .B2(G224), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n828), .A2(new_n794), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n930), .B1(new_n931), .B2(new_n299), .ZN(new_n932));
  INV_X1    g746(.A(G898), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n879), .B1(new_n933), .B2(G953), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n932), .B(new_n934), .ZN(G69));
  OAI21_X1  g749(.A(new_n229), .B1(KEYINPUT30), .B2(new_n263), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT124), .Z(new_n937));
  NAND2_X1  g751(.A1(new_n445), .A2(new_n446), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n937), .B(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n645), .A2(new_n806), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n661), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(KEYINPUT62), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n791), .A2(new_n761), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n670), .A2(new_n649), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n945), .B1(new_n753), .B2(new_n764), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n661), .A2(new_n947), .A3(new_n941), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n943), .A2(new_n775), .A3(new_n946), .A4(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n939), .B1(new_n949), .B2(new_n299), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT125), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n670), .A2(new_n703), .ZN(new_n953));
  OAI211_X1 g767(.A(new_n750), .B(new_n752), .C1(new_n764), .C2(new_n953), .ZN(new_n954));
  AND4_X1   g768(.A1(new_n735), .A2(new_n954), .A3(new_n737), .A4(new_n941), .ZN(new_n955));
  AOI21_X1  g769(.A(G953), .B1(new_n955), .B2(new_n775), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n299), .A2(G900), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n957), .A2(KEYINPUT126), .A3(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n956), .B2(new_n958), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n960), .A2(new_n939), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n299), .B1(G227), .B2(G900), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n952), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n964), .B1(new_n952), .B2(new_n963), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n966), .A2(new_n967), .ZN(G72));
  XOR2_X1   g782(.A(KEYINPUT127), .B(KEYINPUT63), .Z(new_n969));
  NAND2_X1  g783(.A1(G472), .A2(G902), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n955), .A2(new_n775), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n971), .B1(new_n972), .B2(new_n931), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n281), .A2(new_n250), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n884), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n971), .B1(new_n949), .B2(new_n931), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n976), .A2(new_n250), .A3(new_n281), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n283), .A2(new_n255), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n834), .A2(new_n971), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n975), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(G57));
endmodule


