//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 0 0 1 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n602, new_n603, new_n604, new_n605, new_n607, new_n608, new_n609,
    new_n611, new_n612, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  INV_X1    g002(.A(G155gat), .ZN(new_n204));
  INV_X1    g003(.A(G162gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(new_n206), .B2(KEYINPUT2), .ZN(new_n207));
  XOR2_X1   g006(.A(G141gat), .B(G148gat), .Z(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT72), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(new_n203), .A3(new_n206), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n211), .A2(new_n212), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT29), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  XOR2_X1   g018(.A(G211gat), .B(G218gat), .Z(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT71), .ZN(new_n221));
  XNOR2_X1  g020(.A(G197gat), .B(G204gat), .ZN(new_n222));
  INV_X1    g021(.A(G211gat), .ZN(new_n223));
  INV_X1    g022(.A(G218gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n222), .B1(KEYINPUT22), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n221), .B(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n219), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n211), .A2(new_n215), .ZN(new_n230));
  INV_X1    g029(.A(new_n220), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n217), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n226), .A2(new_n231), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n212), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n202), .B1(new_n229), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n212), .B1(new_n227), .B2(KEYINPUT29), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(new_n230), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(G228gat), .A3(G233gat), .ZN(new_n239));
  OAI21_X1  g038(.A(KEYINPUT76), .B1(new_n219), .B2(new_n228), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT76), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n218), .A2(new_n241), .A3(new_n227), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n239), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT77), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  AOI211_X1 g044(.A(KEYINPUT77), .B(new_n239), .C1(new_n240), .C2(new_n242), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n236), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT78), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT78), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n249), .B(new_n236), .C1(new_n245), .C2(new_n246), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(G22gat), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT79), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n247), .A2(G22gat), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G78gat), .B(G106gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(KEYINPUT31), .B(G50gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n248), .A2(KEYINPUT79), .A3(G22gat), .A4(new_n250), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n253), .A2(new_n255), .A3(new_n258), .A4(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n258), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n247), .A2(G22gat), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n261), .B1(new_n262), .B2(new_n254), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(G120gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n265), .A2(G113gat), .ZN(new_n266));
  XOR2_X1   g065(.A(KEYINPUT67), .B(G120gat), .Z(new_n267));
  AOI21_X1  g066(.A(new_n266), .B1(new_n267), .B2(G113gat), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT1), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G127gat), .B(G134gat), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n270), .B(new_n271), .C1(new_n269), .C2(new_n268), .ZN(new_n272));
  INV_X1    g071(.A(new_n271), .ZN(new_n273));
  XNOR2_X1  g072(.A(G113gat), .B(G120gat), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n273), .B1(KEYINPUT1), .B2(new_n274), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n272), .A2(new_n211), .A3(new_n215), .A4(new_n275), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n276), .A2(KEYINPUT4), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n277), .A2(KEYINPUT75), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(KEYINPUT4), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(KEYINPUT75), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n230), .A2(KEYINPUT3), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n272), .A2(new_n275), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(new_n283), .A3(new_n216), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n282), .A2(new_n283), .A3(KEYINPUT73), .A4(new_n216), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n281), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(G225gat), .A2(G233gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n283), .A2(new_n230), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(new_n276), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n292), .B(KEYINPUT39), .C1(new_n291), .C2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G1gat), .B(G29gat), .ZN(new_n296));
  INV_X1    g095(.A(G85gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT0), .B(G57gat), .ZN(new_n299));
  XOR2_X1   g098(.A(new_n298), .B(new_n299), .Z(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n295), .B(new_n301), .C1(KEYINPUT39), .C2(new_n292), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT40), .ZN(new_n303));
  OR2_X1    g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT5), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n281), .A2(new_n305), .A3(new_n290), .A4(new_n288), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n276), .A2(KEYINPUT4), .A3(new_n290), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n277), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n288), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n291), .ZN(new_n311));
  AND4_X1   g110(.A1(new_n307), .A2(new_n310), .A3(KEYINPUT5), .A4(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n305), .B1(new_n288), .B2(new_n309), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n307), .B1(new_n313), .B2(new_n311), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n306), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(new_n300), .ZN(new_n316));
  NOR2_X1   g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(G169gat), .A2(G176gat), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n317), .B1(KEYINPUT23), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n317), .B(KEYINPUT64), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT23), .ZN(new_n322));
  NOR2_X1   g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323));
  XOR2_X1   g122(.A(new_n323), .B(KEYINPUT65), .Z(new_n324));
  NAND2_X1  g123(.A1(G183gat), .A2(G190gat), .ZN(new_n325));
  XOR2_X1   g124(.A(new_n325), .B(KEYINPUT24), .Z(new_n326));
  OAI221_X1 g125(.A(new_n320), .B1(new_n321), .B2(new_n322), .C1(new_n324), .C2(new_n326), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n323), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n328), .A2(new_n319), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT25), .B1(new_n317), .B2(KEYINPUT23), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n327), .A2(KEYINPUT25), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(KEYINPUT27), .B(G183gat), .ZN(new_n332));
  INV_X1    g131(.A(G190gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  XOR2_X1   g133(.A(new_n334), .B(KEYINPUT28), .Z(new_n335));
  NOR2_X1   g134(.A1(new_n321), .A2(KEYINPUT26), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT26), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n317), .B1(new_n337), .B2(new_n318), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n338), .B(KEYINPUT66), .Z(new_n339));
  OAI211_X1 g138(.A(new_n335), .B(new_n325), .C1(new_n336), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n331), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(G226gat), .A2(G233gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(new_n217), .A3(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n343), .B1(new_n342), .B2(new_n341), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(new_n228), .ZN(new_n345));
  XNOR2_X1  g144(.A(G8gat), .B(G36gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(G64gat), .B(G92gat), .ZN(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT30), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n350), .B1(new_n345), .B2(new_n348), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n349), .B(new_n351), .Z(new_n352));
  NAND2_X1  g151(.A1(new_n302), .A2(new_n303), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n304), .A2(new_n316), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT6), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n306), .B(new_n301), .C1(new_n312), .C2(new_n314), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n316), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n315), .A2(KEYINPUT6), .A3(new_n300), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT80), .ZN(new_n360));
  XOR2_X1   g159(.A(new_n345), .B(KEYINPUT37), .Z(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n348), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT38), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT80), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n358), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n360), .A2(new_n349), .A3(new_n363), .A4(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n362), .A2(KEYINPUT38), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n264), .B(new_n354), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n264), .ZN(new_n369));
  INV_X1    g168(.A(new_n352), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n359), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  XOR2_X1   g171(.A(new_n341), .B(new_n283), .Z(new_n373));
  NAND2_X1  g172(.A1(G227gat), .A2(G233gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(G15gat), .B(G43gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n376), .B(G71gat), .ZN(new_n377));
  INV_X1    g176(.A(G99gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(new_n377), .B(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n373), .A2(new_n374), .ZN(new_n380));
  XOR2_X1   g179(.A(KEYINPUT69), .B(KEYINPUT33), .Z(new_n381));
  OAI211_X1 g180(.A(new_n375), .B(new_n379), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(new_n381), .ZN(new_n383));
  INV_X1    g182(.A(new_n379), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n373), .B(new_n374), .C1(new_n383), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT32), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT34), .B1(new_n380), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT34), .ZN(new_n389));
  OAI211_X1 g188(.A(KEYINPUT32), .B(new_n389), .C1(new_n373), .C2(new_n374), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n386), .B(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT70), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(new_n394), .B(KEYINPUT36), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n368), .A2(new_n372), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT81), .ZN(new_n397));
  INV_X1    g196(.A(new_n392), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n264), .A2(new_n370), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT35), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n364), .B1(new_n357), .B2(new_n358), .ZN(new_n401));
  INV_X1    g200(.A(new_n365), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n397), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  AOI211_X1 g203(.A(new_n392), .B(new_n352), .C1(new_n260), .C2(new_n263), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT35), .B1(new_n360), .B2(new_n365), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT81), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n264), .A2(new_n398), .ZN(new_n408));
  OAI21_X1  g207(.A(KEYINPUT35), .B1(new_n408), .B2(new_n371), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n404), .A2(new_n407), .A3(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n396), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT85), .ZN(new_n412));
  INV_X1    g211(.A(G8gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(G15gat), .B(G22gat), .ZN(new_n414));
  INV_X1    g213(.A(G1gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT16), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n414), .A2(G1gat), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n412), .B(new_n413), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  OR2_X1    g218(.A1(new_n414), .A2(G1gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n414), .A2(new_n416), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n412), .A2(new_n413), .ZN(new_n422));
  NAND2_X1  g221(.A1(KEYINPUT85), .A2(G8gat), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n420), .A2(new_n421), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT87), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n425), .A2(new_n426), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT21), .ZN(new_n430));
  XOR2_X1   g229(.A(G71gat), .B(G78gat), .Z(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT9), .ZN(new_n433));
  INV_X1    g232(.A(G71gat), .ZN(new_n434));
  INV_X1    g233(.A(G78gat), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(G57gat), .B(G64gat), .Z(new_n437));
  NAND3_X1  g236(.A1(new_n432), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n436), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n431), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  OAI22_X1  g240(.A1(new_n428), .A2(new_n429), .B1(new_n430), .B2(new_n441), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n442), .B(G183gat), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n441), .A2(new_n430), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(new_n223), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n445), .B(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G127gat), .B(G155gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(G231gat), .A2(G233gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n448), .B(new_n451), .ZN(new_n452));
  AND2_X1   g251(.A1(G232gat), .A2(G233gat), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT41), .ZN(new_n454));
  INV_X1    g253(.A(G92gat), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT91), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n456), .A2(G85gat), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n297), .A2(KEYINPUT91), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n455), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  OR2_X1    g258(.A1(KEYINPUT90), .A2(KEYINPUT7), .ZN(new_n460));
  NAND2_X1  g259(.A1(G85gat), .A2(G92gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(KEYINPUT90), .A2(KEYINPUT7), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  OR2_X1    g263(.A1(G99gat), .A2(G106gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(G99gat), .A2(G106gat), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OR2_X1    g266(.A1(new_n467), .A2(KEYINPUT92), .ZN(new_n468));
  OR2_X1    g267(.A1(new_n461), .A2(new_n462), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT92), .B1(G99gat), .B2(G106gat), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT8), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(new_n466), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n464), .A2(new_n468), .A3(new_n469), .A4(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n473), .A2(new_n459), .A3(new_n469), .A4(new_n463), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n467), .A2(KEYINPUT92), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  OR3_X1    g277(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n479), .A2(new_n480), .B1(G29gat), .B2(G36gat), .ZN(new_n481));
  INV_X1    g280(.A(G50gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(G43gat), .ZN(new_n483));
  INV_X1    g282(.A(G43gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(G50gat), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT83), .ZN(new_n486));
  AND3_X1   g285(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n486), .B1(new_n483), .B2(new_n485), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT15), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G43gat), .B(G50gat), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(KEYINPUT15), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n481), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n483), .A2(new_n485), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT83), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n491), .A2(new_n486), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n495), .A2(new_n496), .A3(KEYINPUT15), .ZN(new_n497));
  INV_X1    g296(.A(new_n481), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n478), .A2(new_n493), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT84), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT17), .ZN(new_n502));
  INV_X1    g301(.A(new_n492), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n498), .B1(new_n497), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n490), .A2(new_n481), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n501), .B(new_n502), .C1(new_n504), .C2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(KEYINPUT84), .A2(KEYINPUT17), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n501), .A2(new_n502), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n493), .A2(new_n499), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n454), .B(new_n500), .C1(new_n511), .C2(new_n478), .ZN(new_n512));
  XNOR2_X1  g311(.A(G190gat), .B(G218gat), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n512), .B(new_n513), .Z(new_n514));
  OR2_X1    g313(.A1(new_n453), .A2(KEYINPUT41), .ZN(new_n515));
  XNOR2_X1  g314(.A(G134gat), .B(G162gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  OR2_X1    g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n514), .A2(new_n517), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n452), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n510), .A2(new_n425), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT86), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n419), .A2(new_n424), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT87), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n527), .A2(new_n493), .A3(new_n499), .A4(new_n427), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT88), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT18), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n510), .A2(KEYINPUT86), .A3(new_n425), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n525), .A2(new_n528), .A3(new_n531), .A4(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G229gat), .A2(G233gat), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  OAI22_X1  g334(.A1(new_n533), .A2(new_n535), .B1(new_n529), .B2(new_n530), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT86), .B1(new_n510), .B2(new_n425), .ZN(new_n537));
  AOI211_X1 g336(.A(new_n524), .B(new_n526), .C1(new_n506), .C2(new_n509), .ZN(new_n538));
  INV_X1    g337(.A(new_n528), .ZN(new_n539));
  NOR3_X1   g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n540), .A2(KEYINPUT88), .A3(KEYINPUT18), .A4(new_n534), .ZN(new_n541));
  OAI22_X1  g340(.A1(new_n428), .A2(new_n429), .B1(new_n504), .B2(new_n505), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n528), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n534), .B(KEYINPUT13), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT89), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n543), .A2(KEYINPUT89), .A3(new_n545), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n536), .A2(new_n541), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT82), .ZN(new_n552));
  XNOR2_X1  g351(.A(G113gat), .B(G141gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(G197gat), .ZN(new_n554));
  XOR2_X1   g353(.A(KEYINPUT11), .B(G169gat), .Z(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  XOR2_X1   g355(.A(new_n556), .B(KEYINPUT12), .Z(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n551), .A2(new_n552), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n558), .B1(new_n551), .B2(new_n552), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  AND2_X1   g361(.A1(new_n438), .A2(new_n440), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n475), .A2(new_n476), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n475), .A2(new_n476), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n563), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT10), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n474), .A2(new_n441), .A3(new_n477), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT93), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n478), .A2(KEYINPUT10), .A3(new_n563), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n566), .A2(KEYINPUT93), .A3(new_n568), .A4(new_n567), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G230gat), .A2(G233gat), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n566), .A2(new_n568), .ZN(new_n577));
  INV_X1    g376(.A(new_n575), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G120gat), .B(G148gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT94), .ZN(new_n582));
  XNOR2_X1  g381(.A(G176gat), .B(G204gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n582), .B(new_n583), .Z(new_n584));
  OAI21_X1  g383(.A(KEYINPUT95), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT95), .ZN(new_n586));
  INV_X1    g385(.A(new_n584), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n576), .A2(new_n586), .A3(new_n579), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n580), .A2(new_n584), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n562), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n522), .A2(new_n593), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n411), .A2(KEYINPUT96), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(KEYINPUT96), .B1(new_n411), .B2(new_n594), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n359), .B(KEYINPUT97), .Z(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(KEYINPUT98), .B(G1gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(G1324gat));
  NOR2_X1   g400(.A1(new_n597), .A2(new_n370), .ZN(new_n602));
  XOR2_X1   g401(.A(KEYINPUT16), .B(G8gat), .Z(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT42), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n605), .B1(new_n413), .B2(new_n602), .ZN(G1325gat));
  INV_X1    g405(.A(new_n597), .ZN(new_n607));
  AOI21_X1  g406(.A(G15gat), .B1(new_n607), .B2(new_n398), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n597), .A2(new_n395), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n608), .B1(G15gat), .B2(new_n609), .ZN(G1326gat));
  NOR2_X1   g409(.A1(new_n597), .A2(new_n264), .ZN(new_n611));
  XOR2_X1   g410(.A(KEYINPUT43), .B(G22gat), .Z(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(G1327gat));
  AOI21_X1  g412(.A(new_n521), .B1(new_n396), .B2(new_n410), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n593), .A2(new_n452), .ZN(new_n615));
  AND2_X1   g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(G29gat), .ZN(new_n617));
  INV_X1    g416(.A(new_n598), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT45), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n411), .A2(new_n520), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n621), .A2(KEYINPUT44), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT44), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n614), .A2(new_n623), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(new_n618), .A3(new_n615), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n620), .B1(new_n627), .B2(new_n617), .ZN(G1328gat));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n615), .ZN(new_n629));
  OAI21_X1  g428(.A(G36gat), .B1(new_n629), .B2(new_n370), .ZN(new_n630));
  INV_X1    g429(.A(G36gat), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n616), .A2(new_n631), .A3(new_n352), .ZN(new_n632));
  XOR2_X1   g431(.A(KEYINPUT99), .B(KEYINPUT46), .Z(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n630), .A2(new_n634), .ZN(G1329gat));
  INV_X1    g434(.A(new_n395), .ZN(new_n636));
  OAI211_X1 g435(.A(new_n636), .B(new_n615), .C1(new_n622), .C2(new_n624), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(G43gat), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n616), .A2(new_n484), .A3(new_n398), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT101), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT100), .B1(new_n637), .B2(G43gat), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n643), .A2(KEYINPUT47), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n642), .B(new_n644), .ZN(G1330gat));
  INV_X1    g444(.A(KEYINPUT102), .ZN(new_n646));
  OAI21_X1  g445(.A(G50gat), .B1(new_n629), .B2(new_n264), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n616), .A2(new_n482), .A3(new_n369), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n649), .B(KEYINPUT48), .Z(G1331gat));
  NOR2_X1   g449(.A1(new_n522), .A2(new_n562), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(new_n591), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT103), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n411), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n618), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g455(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n654), .A2(new_n352), .A3(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n658), .B(new_n659), .Z(G1333gat));
  AOI21_X1  g459(.A(new_n434), .B1(new_n654), .B2(new_n636), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n392), .B(KEYINPUT104), .Z(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(G71gat), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n661), .B1(new_n654), .B2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g464(.A1(new_n654), .A2(new_n369), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT105), .B(G78gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1335gat));
  OR2_X1    g467(.A1(new_n457), .A2(new_n458), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n622), .A2(new_n624), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(new_n592), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n452), .A2(new_n562), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n670), .B1(new_n674), .B2(new_n598), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n621), .A2(KEYINPUT106), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n614), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n676), .A2(new_n673), .A3(new_n678), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n679), .A2(KEYINPUT51), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(KEYINPUT51), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n680), .A2(new_n591), .A3(new_n618), .A4(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n675), .B1(new_n670), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT107), .ZN(G1336gat));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n676), .A2(new_n685), .A3(new_n673), .A4(new_n678), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT109), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT51), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n370), .A2(G92gat), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n685), .B1(new_n689), .B2(KEYINPUT109), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n679), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n690), .A2(new_n591), .A3(new_n691), .A4(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT110), .ZN(new_n695));
  OAI21_X1  g494(.A(G92gat), .B1(new_n674), .B2(new_n370), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n688), .A2(new_n689), .B1(new_n679), .B2(new_n692), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT110), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n697), .A2(new_n698), .A3(new_n591), .A4(new_n691), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n695), .A2(new_n696), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT52), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT52), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n680), .A2(new_n591), .A3(new_n681), .ZN(new_n703));
  INV_X1    g502(.A(new_n691), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n696), .B(new_n702), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n701), .A2(new_n705), .ZN(G1337gat));
  NOR2_X1   g505(.A1(new_n674), .A2(new_n395), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT111), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n398), .A2(new_n378), .ZN(new_n709));
  OAI22_X1  g508(.A1(new_n708), .A2(new_n378), .B1(new_n703), .B2(new_n709), .ZN(G1338gat));
  NAND3_X1  g509(.A1(new_n672), .A2(new_n369), .A3(new_n673), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT112), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT112), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n672), .A2(new_n713), .A3(new_n369), .A4(new_n673), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n712), .A2(new_n714), .A3(G106gat), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT53), .ZN(new_n716));
  NOR3_X1   g515(.A1(new_n264), .A2(G106gat), .A3(new_n592), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n680), .A2(new_n681), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n715), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  AOI22_X1  g518(.A1(new_n697), .A2(new_n717), .B1(new_n711), .B2(G106gat), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n719), .B1(new_n716), .B2(new_n720), .ZN(G1339gat));
  NAND2_X1  g520(.A1(new_n651), .A2(new_n592), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n571), .A2(new_n578), .A3(new_n572), .A4(new_n573), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n576), .A2(KEYINPUT54), .A3(new_n724), .ZN(new_n725));
  XOR2_X1   g524(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n726));
  NAND3_X1  g525(.A1(new_n574), .A2(new_n575), .A3(new_n726), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n725), .A2(KEYINPUT55), .A3(new_n584), .A4(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT114), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n727), .A2(new_n584), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n732), .A2(KEYINPUT114), .A3(KEYINPUT55), .A4(new_n725), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n730), .A2(new_n589), .A3(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT115), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT55), .ZN(new_n737));
  INV_X1    g536(.A(new_n725), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n738), .B2(new_n731), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n730), .A2(new_n733), .A3(new_n589), .A4(KEYINPUT115), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n736), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT116), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n736), .A2(KEYINPUT116), .A3(new_n739), .A4(new_n740), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n743), .A2(new_n562), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n540), .A2(new_n534), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n543), .A2(new_n545), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n556), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n591), .B(new_n748), .C1(new_n551), .C2(new_n557), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n520), .B1(new_n745), .B2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n748), .B1(new_n551), .B2(new_n557), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n521), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n743), .A2(new_n753), .A3(new_n744), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT117), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n743), .A2(KEYINPUT117), .A3(new_n753), .A4(new_n744), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n751), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n452), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n723), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OR3_X1    g560(.A1(new_n761), .A2(new_n408), .A3(new_n598), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(new_n352), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n562), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n591), .ZN(new_n766));
  MUX2_X1   g565(.A(new_n267), .B(G120gat), .S(new_n766), .Z(G1341gat));
  NAND2_X1  g566(.A1(new_n763), .A2(new_n452), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G127gat), .ZN(G1342gat));
  NOR2_X1   g568(.A1(new_n352), .A2(new_n521), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT118), .ZN(new_n771));
  OR3_X1    g570(.A1(new_n762), .A2(G134gat), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT56), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(KEYINPUT119), .ZN(new_n774));
  INV_X1    g573(.A(new_n763), .ZN(new_n775));
  OAI21_X1  g574(.A(G134gat), .B1(new_n775), .B2(new_n521), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n774), .B(new_n776), .C1(KEYINPUT56), .C2(new_n772), .ZN(G1343gat));
  INV_X1    g576(.A(KEYINPUT120), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n756), .A2(new_n757), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n760), .B1(new_n779), .B2(new_n750), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n264), .B1(new_n780), .B2(new_n722), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n778), .B1(new_n781), .B2(KEYINPUT57), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT57), .ZN(new_n783));
  OAI211_X1 g582(.A(KEYINPUT120), .B(new_n783), .C1(new_n761), .C2(new_n264), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n730), .A2(new_n739), .A3(new_n733), .A4(new_n589), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n785), .A2(new_n559), .A3(new_n560), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n592), .A2(new_n752), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT121), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT121), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n789), .B(new_n749), .C1(new_n561), .C2(new_n785), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n788), .A2(new_n790), .A3(new_n521), .ZN(new_n791));
  OAI211_X1 g590(.A(KEYINPUT122), .B(new_n760), .C1(new_n779), .C2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT122), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n791), .B1(new_n756), .B2(new_n757), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n794), .B2(new_n452), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n792), .A2(new_n722), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n796), .A2(KEYINPUT57), .A3(new_n369), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n782), .A2(new_n784), .A3(new_n797), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n636), .A2(new_n598), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n370), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(G141gat), .A3(new_n562), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n781), .A2(new_n801), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n804), .A2(new_n561), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(G141gat), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n806), .B(new_n807), .ZN(G1344gat));
  INV_X1    g607(.A(KEYINPUT59), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT57), .B1(new_n761), .B2(new_n264), .ZN(new_n810));
  INV_X1    g609(.A(new_n791), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n753), .A2(new_n739), .A3(new_n736), .A4(new_n740), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n452), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n783), .B(new_n369), .C1(new_n813), .C2(new_n723), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n810), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n815), .A2(new_n591), .A3(new_n801), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n809), .B1(new_n816), .B2(G148gat), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n798), .A2(new_n591), .A3(new_n801), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n809), .A2(G148gat), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT123), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT123), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n818), .A2(new_n822), .A3(new_n819), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n817), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n804), .A2(G148gat), .A3(new_n592), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT124), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT124), .ZN(new_n827));
  INV_X1    g626(.A(new_n825), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n818), .A2(new_n822), .A3(new_n819), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n822), .B1(new_n818), .B2(new_n819), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n827), .B(new_n828), .C1(new_n831), .C2(new_n817), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n826), .A2(new_n832), .ZN(G1345gat));
  INV_X1    g632(.A(new_n804), .ZN(new_n834));
  AOI21_X1  g633(.A(G155gat), .B1(new_n834), .B2(new_n452), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n760), .A2(new_n204), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n835), .B1(new_n802), .B2(new_n836), .ZN(G1346gat));
  NOR2_X1   g636(.A1(new_n771), .A2(G162gat), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n781), .A2(new_n799), .A3(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n802), .A2(new_n520), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(new_n205), .ZN(G1347gat));
  NOR2_X1   g640(.A1(new_n761), .A2(new_n618), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n662), .A2(new_n369), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n352), .A3(new_n843), .ZN(new_n844));
  OAI21_X1  g643(.A(G169gat), .B1(new_n844), .B2(new_n561), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n408), .A2(new_n370), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(KEYINPUT125), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n848), .A2(G169gat), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n845), .B1(new_n849), .B2(new_n561), .ZN(G1348gat));
  INV_X1    g649(.A(new_n848), .ZN(new_n851));
  AOI21_X1  g650(.A(G176gat), .B1(new_n851), .B2(new_n591), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n844), .A2(new_n592), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(G176gat), .B2(new_n853), .ZN(G1349gat));
  NAND3_X1  g653(.A1(new_n851), .A2(new_n332), .A3(new_n452), .ZN(new_n855));
  OAI21_X1  g654(.A(G183gat), .B1(new_n844), .B2(new_n760), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g657(.A(KEYINPUT61), .ZN(new_n859));
  OAI221_X1 g658(.A(G190gat), .B1(KEYINPUT126), .B2(new_n859), .C1(new_n844), .C2(new_n521), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(KEYINPUT126), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n860), .B(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n851), .A2(new_n333), .A3(new_n520), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(G1351gat));
  INV_X1    g663(.A(G197gat), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n618), .A2(new_n636), .A3(new_n370), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n815), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n865), .B1(new_n867), .B2(new_n562), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n781), .A2(new_n866), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n869), .A2(G197gat), .A3(new_n561), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n868), .A2(new_n870), .ZN(G1352gat));
  NOR3_X1   g670(.A1(new_n869), .A2(G204gat), .A3(new_n592), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT62), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n815), .A2(new_n591), .A3(new_n866), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(G204gat), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(G1353gat));
  NAND2_X1  g675(.A1(new_n867), .A2(new_n452), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n877), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n878));
  AOI21_X1  g677(.A(KEYINPUT63), .B1(new_n877), .B2(G211gat), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n452), .A2(new_n223), .ZN(new_n880));
  OAI22_X1  g679(.A1(new_n878), .A2(new_n879), .B1(new_n869), .B2(new_n880), .ZN(G1354gat));
  OAI21_X1  g680(.A(new_n224), .B1(new_n869), .B2(new_n521), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n882), .B(KEYINPUT127), .Z(new_n883));
  NOR2_X1   g682(.A1(new_n521), .A2(new_n224), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n883), .B1(new_n867), .B2(new_n884), .ZN(G1355gat));
endmodule


