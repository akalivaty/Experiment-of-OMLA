

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581;

  XNOR2_X1 U321 ( .A(n447), .B(n446), .ZN(n471) );
  AND2_X1 U322 ( .A1(G230GAT), .A2(G233GAT), .ZN(n289) );
  NAND2_X1 U323 ( .A1(n370), .A2(n369), .ZN(n456) );
  XNOR2_X1 U324 ( .A(n295), .B(KEYINPUT24), .ZN(n296) );
  XNOR2_X1 U325 ( .A(n430), .B(n289), .ZN(n432) );
  XNOR2_X1 U326 ( .A(n297), .B(n296), .ZN(n300) );
  XNOR2_X1 U327 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U328 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U329 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U330 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U331 ( .A(n440), .B(n439), .ZN(n444) );
  XNOR2_X1 U332 ( .A(n504), .B(KEYINPUT41), .ZN(n533) );
  AND2_X1 U333 ( .A1(n488), .A2(n459), .ZN(n446) );
  NOR2_X1 U334 ( .A1(n550), .A2(n549), .ZN(n561) );
  INV_X1 U335 ( .A(G50GAT), .ZN(n448) );
  XNOR2_X1 U336 ( .A(n448), .B(KEYINPUT108), .ZN(n449) );
  XNOR2_X1 U337 ( .A(n450), .B(n449), .ZN(G1331GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT86), .B(G197GAT), .Z(n291) );
  XNOR2_X1 U339 ( .A(G218GAT), .B(KEYINPUT21), .ZN(n290) );
  XNOR2_X1 U340 ( .A(n291), .B(n290), .ZN(n292) );
  XOR2_X1 U341 ( .A(G211GAT), .B(n292), .Z(n323) );
  XOR2_X1 U342 ( .A(G162GAT), .B(G50GAT), .Z(n396) );
  XOR2_X1 U343 ( .A(G141GAT), .B(KEYINPUT87), .Z(n294) );
  XNOR2_X1 U344 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n293) );
  XNOR2_X1 U345 ( .A(n294), .B(n293), .ZN(n346) );
  XOR2_X1 U346 ( .A(n396), .B(n346), .Z(n297) );
  NAND2_X1 U347 ( .A1(G228GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U348 ( .A(G148GAT), .B(G106GAT), .ZN(n298) );
  XNOR2_X1 U349 ( .A(n298), .B(G78GAT), .ZN(n442) );
  XOR2_X1 U350 ( .A(n442), .B(KEYINPUT22), .Z(n299) );
  XNOR2_X1 U351 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U352 ( .A(G155GAT), .B(G22GAT), .Z(n384) );
  XNOR2_X1 U353 ( .A(n384), .B(KEYINPUT23), .ZN(n302) );
  INV_X1 U354 ( .A(G204GAT), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n323), .B(n305), .ZN(n334) );
  XNOR2_X1 U356 ( .A(KEYINPUT28), .B(n334), .ZN(n494) );
  XNOR2_X1 U357 ( .A(KEYINPUT105), .B(KEYINPUT38), .ZN(n447) );
  XNOR2_X1 U358 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n306) );
  XNOR2_X1 U359 ( .A(n306), .B(G169GAT), .ZN(n307) );
  XOR2_X1 U360 ( .A(n307), .B(KEYINPUT85), .Z(n309) );
  XNOR2_X1 U361 ( .A(G183GAT), .B(KEYINPUT19), .ZN(n308) );
  XNOR2_X1 U362 ( .A(n309), .B(n308), .ZN(n322) );
  XOR2_X1 U363 ( .A(G120GAT), .B(G71GAT), .Z(n434) );
  XOR2_X1 U364 ( .A(n434), .B(G176GAT), .Z(n311) );
  NAND2_X1 U365 ( .A1(G227GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U366 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U367 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n313) );
  XNOR2_X1 U368 ( .A(G134GAT), .B(G43GAT), .ZN(n312) );
  XNOR2_X1 U369 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U370 ( .A(n315), .B(n314), .Z(n319) );
  XOR2_X1 U371 ( .A(KEYINPUT0), .B(G113GAT), .Z(n342) );
  XNOR2_X1 U372 ( .A(G190GAT), .B(G99GAT), .ZN(n316) );
  XOR2_X1 U373 ( .A(G127GAT), .B(G15GAT), .Z(n385) );
  XNOR2_X1 U374 ( .A(n316), .B(n385), .ZN(n317) );
  XNOR2_X1 U375 ( .A(n342), .B(n317), .ZN(n318) );
  XNOR2_X1 U376 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U377 ( .A(n322), .B(n320), .ZN(n550) );
  INV_X1 U378 ( .A(n334), .ZN(n547) );
  NAND2_X1 U379 ( .A1(n550), .A2(n547), .ZN(n321) );
  XNOR2_X1 U380 ( .A(n321), .B(KEYINPUT26), .ZN(n567) );
  XNOR2_X1 U381 ( .A(n323), .B(n322), .ZN(n332) );
  XOR2_X1 U382 ( .A(G176GAT), .B(G204GAT), .Z(n325) );
  XNOR2_X1 U383 ( .A(G92GAT), .B(G64GAT), .ZN(n324) );
  XNOR2_X1 U384 ( .A(n325), .B(n324), .ZN(n441) );
  XOR2_X1 U385 ( .A(KEYINPUT92), .B(n441), .Z(n327) );
  NAND2_X1 U386 ( .A1(G226GAT), .A2(G233GAT), .ZN(n326) );
  XNOR2_X1 U387 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U388 ( .A(n328), .B(KEYINPUT93), .Z(n330) );
  XOR2_X1 U389 ( .A(G190GAT), .B(G36GAT), .Z(n399) );
  XNOR2_X1 U390 ( .A(n399), .B(G8GAT), .ZN(n329) );
  XNOR2_X1 U391 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U392 ( .A(n332), .B(n331), .ZN(n490) );
  XNOR2_X1 U393 ( .A(n490), .B(KEYINPUT27), .ZN(n365) );
  NOR2_X1 U394 ( .A1(n567), .A2(n365), .ZN(n333) );
  XNOR2_X1 U395 ( .A(n333), .B(KEYINPUT97), .ZN(n340) );
  XNOR2_X1 U396 ( .A(KEYINPUT25), .B(KEYINPUT99), .ZN(n338) );
  INV_X1 U397 ( .A(n490), .ZN(n541) );
  INV_X1 U398 ( .A(n550), .ZN(n512) );
  NAND2_X1 U399 ( .A1(n541), .A2(n512), .ZN(n335) );
  NAND2_X1 U400 ( .A1(n335), .A2(n334), .ZN(n336) );
  XNOR2_X1 U401 ( .A(n336), .B(KEYINPUT98), .ZN(n337) );
  XNOR2_X1 U402 ( .A(n338), .B(n337), .ZN(n339) );
  NAND2_X1 U403 ( .A1(n340), .A2(n339), .ZN(n341) );
  XNOR2_X1 U404 ( .A(KEYINPUT100), .B(n341), .ZN(n364) );
  XOR2_X1 U405 ( .A(G162GAT), .B(G85GAT), .Z(n344) );
  XOR2_X1 U406 ( .A(KEYINPUT78), .B(G134GAT), .Z(n407) );
  XNOR2_X1 U407 ( .A(n407), .B(n342), .ZN(n343) );
  XNOR2_X1 U408 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U409 ( .A(n345), .B(G120GAT), .Z(n351) );
  XOR2_X1 U410 ( .A(n346), .B(KEYINPUT5), .Z(n348) );
  NAND2_X1 U411 ( .A1(G225GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U412 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U413 ( .A(G29GAT), .B(n349), .ZN(n350) );
  XNOR2_X1 U414 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U415 ( .A(G57GAT), .B(G155GAT), .Z(n353) );
  XNOR2_X1 U416 ( .A(G127GAT), .B(G148GAT), .ZN(n352) );
  XNOR2_X1 U417 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U418 ( .A(n355), .B(n354), .Z(n363) );
  XOR2_X1 U419 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n357) );
  XNOR2_X1 U420 ( .A(KEYINPUT91), .B(KEYINPUT1), .ZN(n356) );
  XNOR2_X1 U421 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U422 ( .A(KEYINPUT88), .B(KEYINPUT4), .Z(n359) );
  XNOR2_X1 U423 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n358) );
  XNOR2_X1 U424 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U425 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n363), .B(n362), .ZN(n545) );
  NAND2_X1 U427 ( .A1(n364), .A2(n545), .ZN(n370) );
  NOR2_X1 U428 ( .A1(n545), .A2(n365), .ZN(n366) );
  XNOR2_X1 U429 ( .A(KEYINPUT94), .B(n366), .ZN(n527) );
  NAND2_X1 U430 ( .A1(n494), .A2(n527), .ZN(n514) );
  XNOR2_X1 U431 ( .A(KEYINPUT95), .B(n514), .ZN(n367) );
  NAND2_X1 U432 ( .A1(n367), .A2(n550), .ZN(n368) );
  XNOR2_X1 U433 ( .A(n368), .B(KEYINPUT96), .ZN(n369) );
  XOR2_X1 U434 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n372) );
  XNOR2_X1 U435 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n371) );
  XNOR2_X1 U436 ( .A(n372), .B(n371), .ZN(n389) );
  XOR2_X1 U437 ( .A(KEYINPUT81), .B(KEYINPUT80), .Z(n374) );
  NAND2_X1 U438 ( .A1(G231GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U439 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U440 ( .A(n375), .B(KEYINPUT82), .Z(n379) );
  XNOR2_X1 U441 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n376) );
  XNOR2_X1 U442 ( .A(n376), .B(KEYINPUT72), .ZN(n431) );
  XNOR2_X1 U443 ( .A(G1GAT), .B(G8GAT), .ZN(n377) );
  XNOR2_X1 U444 ( .A(n377), .B(KEYINPUT71), .ZN(n422) );
  XNOR2_X1 U445 ( .A(n431), .B(n422), .ZN(n378) );
  XNOR2_X1 U446 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U447 ( .A(G211GAT), .B(G78GAT), .Z(n381) );
  XNOR2_X1 U448 ( .A(G71GAT), .B(G183GAT), .ZN(n380) );
  XNOR2_X1 U449 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U450 ( .A(n383), .B(n382), .Z(n387) );
  XNOR2_X1 U451 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U452 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U453 ( .A(n389), .B(n388), .Z(n501) );
  NAND2_X1 U454 ( .A1(n456), .A2(n501), .ZN(n390) );
  XOR2_X1 U455 ( .A(KEYINPUT104), .B(n390), .Z(n412) );
  XOR2_X1 U456 ( .A(KEYINPUT77), .B(KEYINPUT79), .Z(n392) );
  XNOR2_X1 U457 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n391) );
  XNOR2_X1 U458 ( .A(n392), .B(n391), .ZN(n411) );
  XOR2_X1 U459 ( .A(KEYINPUT67), .B(KEYINPUT9), .Z(n394) );
  XNOR2_X1 U460 ( .A(G106GAT), .B(G92GAT), .ZN(n393) );
  XNOR2_X1 U461 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U462 ( .A(n395), .B(KEYINPUT66), .Z(n398) );
  XNOR2_X1 U463 ( .A(n396), .B(G218GAT), .ZN(n397) );
  XNOR2_X1 U464 ( .A(n398), .B(n397), .ZN(n403) );
  XOR2_X1 U465 ( .A(G85GAT), .B(G99GAT), .Z(n430) );
  XOR2_X1 U466 ( .A(n399), .B(n430), .Z(n401) );
  NAND2_X1 U467 ( .A1(G232GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U468 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U469 ( .A(n403), .B(n402), .Z(n409) );
  XOR2_X1 U470 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n405) );
  XNOR2_X1 U471 ( .A(KEYINPUT70), .B(G43GAT), .ZN(n404) );
  XNOR2_X1 U472 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U473 ( .A(G29GAT), .B(n406), .Z(n423) );
  XNOR2_X1 U474 ( .A(n407), .B(n423), .ZN(n408) );
  XNOR2_X1 U475 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U476 ( .A(n411), .B(n410), .ZN(n560) );
  XNOR2_X1 U477 ( .A(KEYINPUT36), .B(n560), .ZN(n578) );
  NAND2_X1 U478 ( .A1(n412), .A2(n578), .ZN(n413) );
  XNOR2_X1 U479 ( .A(n413), .B(KEYINPUT37), .ZN(n488) );
  NAND2_X1 U480 ( .A1(G229GAT), .A2(G233GAT), .ZN(n419) );
  XOR2_X1 U481 ( .A(G169GAT), .B(G15GAT), .Z(n415) );
  XNOR2_X1 U482 ( .A(G141GAT), .B(G113GAT), .ZN(n414) );
  XNOR2_X1 U483 ( .A(n415), .B(n414), .ZN(n417) );
  XOR2_X1 U484 ( .A(G36GAT), .B(G50GAT), .Z(n416) );
  XNOR2_X1 U485 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U486 ( .A(n419), .B(n418), .ZN(n429) );
  XOR2_X1 U487 ( .A(KEYINPUT68), .B(KEYINPUT69), .Z(n421) );
  XNOR2_X1 U488 ( .A(G22GAT), .B(G197GAT), .ZN(n420) );
  XNOR2_X1 U489 ( .A(n421), .B(n420), .ZN(n427) );
  XOR2_X1 U490 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n425) );
  XNOR2_X1 U491 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U492 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U493 ( .A(n427), .B(n426), .Z(n428) );
  XNOR2_X1 U494 ( .A(n429), .B(n428), .ZN(n568) );
  XOR2_X1 U495 ( .A(n433), .B(KEYINPUT75), .Z(n440) );
  XNOR2_X1 U496 ( .A(n434), .B(KEYINPUT33), .ZN(n438) );
  XOR2_X1 U497 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n436) );
  XNOR2_X1 U498 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n435) );
  XNOR2_X1 U499 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U500 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U501 ( .A(n444), .B(n443), .ZN(n572) );
  INV_X1 U502 ( .A(n572), .ZN(n504) );
  NAND2_X1 U503 ( .A1(n568), .A2(n504), .ZN(n445) );
  XOR2_X1 U504 ( .A(KEYINPUT76), .B(n445), .Z(n459) );
  NOR2_X1 U505 ( .A1(n494), .A2(n471), .ZN(n450) );
  INV_X1 U506 ( .A(G36GAT), .ZN(n453) );
  NOR2_X1 U507 ( .A1(n490), .A2(n471), .ZN(n451) );
  XNOR2_X1 U508 ( .A(KEYINPUT106), .B(n451), .ZN(n452) );
  XNOR2_X1 U509 ( .A(n453), .B(n452), .ZN(G1329GAT) );
  NOR2_X1 U510 ( .A1(n501), .A2(n560), .ZN(n454) );
  XOR2_X1 U511 ( .A(KEYINPUT16), .B(n454), .Z(n455) );
  XNOR2_X1 U512 ( .A(KEYINPUT83), .B(n455), .ZN(n457) );
  NAND2_X1 U513 ( .A1(n457), .A2(n456), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n458), .B(KEYINPUT101), .ZN(n476) );
  NAND2_X1 U515 ( .A1(n476), .A2(n459), .ZN(n466) );
  NOR2_X1 U516 ( .A1(n545), .A2(n466), .ZN(n460) );
  XOR2_X1 U517 ( .A(KEYINPUT34), .B(n460), .Z(n461) );
  XNOR2_X1 U518 ( .A(G1GAT), .B(n461), .ZN(G1324GAT) );
  NOR2_X1 U519 ( .A1(n490), .A2(n466), .ZN(n462) );
  XOR2_X1 U520 ( .A(G8GAT), .B(n462), .Z(G1325GAT) );
  NOR2_X1 U521 ( .A1(n550), .A2(n466), .ZN(n464) );
  XNOR2_X1 U522 ( .A(KEYINPUT102), .B(KEYINPUT35), .ZN(n463) );
  XNOR2_X1 U523 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U524 ( .A(G15GAT), .B(n465), .ZN(G1326GAT) );
  NOR2_X1 U525 ( .A1(n494), .A2(n466), .ZN(n468) );
  XNOR2_X1 U526 ( .A(G22GAT), .B(KEYINPUT103), .ZN(n467) );
  XNOR2_X1 U527 ( .A(n468), .B(n467), .ZN(G1327GAT) );
  XNOR2_X1 U528 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n470) );
  NOR2_X1 U529 ( .A1(n545), .A2(n471), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n470), .B(n469), .ZN(G1328GAT) );
  NOR2_X1 U531 ( .A1(n471), .A2(n550), .ZN(n473) );
  XNOR2_X1 U532 ( .A(KEYINPUT40), .B(KEYINPUT107), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U534 ( .A(G43GAT), .B(n474), .ZN(G1330GAT) );
  XOR2_X1 U535 ( .A(KEYINPUT109), .B(n533), .Z(n554) );
  INV_X1 U536 ( .A(n554), .ZN(n475) );
  NOR2_X1 U537 ( .A1(n568), .A2(n475), .ZN(n487) );
  NAND2_X1 U538 ( .A1(n487), .A2(n476), .ZN(n482) );
  NOR2_X1 U539 ( .A1(n545), .A2(n482), .ZN(n477) );
  XOR2_X1 U540 ( .A(G57GAT), .B(n477), .Z(n478) );
  XNOR2_X1 U541 ( .A(KEYINPUT42), .B(n478), .ZN(G1332GAT) );
  NOR2_X1 U542 ( .A1(n490), .A2(n482), .ZN(n479) );
  XOR2_X1 U543 ( .A(KEYINPUT110), .B(n479), .Z(n480) );
  XNOR2_X1 U544 ( .A(G64GAT), .B(n480), .ZN(G1333GAT) );
  NOR2_X1 U545 ( .A1(n550), .A2(n482), .ZN(n481) );
  XOR2_X1 U546 ( .A(G71GAT), .B(n481), .Z(G1334GAT) );
  NOR2_X1 U547 ( .A1(n482), .A2(n494), .ZN(n486) );
  XOR2_X1 U548 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n484) );
  XNOR2_X1 U549 ( .A(G78GAT), .B(KEYINPUT112), .ZN(n483) );
  XNOR2_X1 U550 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U551 ( .A(n486), .B(n485), .ZN(G1335GAT) );
  NAND2_X1 U552 ( .A1(n488), .A2(n487), .ZN(n493) );
  NOR2_X1 U553 ( .A1(n545), .A2(n493), .ZN(n489) );
  XOR2_X1 U554 ( .A(G85GAT), .B(n489), .Z(G1336GAT) );
  NOR2_X1 U555 ( .A1(n490), .A2(n493), .ZN(n491) );
  XOR2_X1 U556 ( .A(G92GAT), .B(n491), .Z(G1337GAT) );
  NOR2_X1 U557 ( .A1(n550), .A2(n493), .ZN(n492) );
  XOR2_X1 U558 ( .A(G99GAT), .B(n492), .Z(G1338GAT) );
  NOR2_X1 U559 ( .A1(n494), .A2(n493), .ZN(n495) );
  XOR2_X1 U560 ( .A(KEYINPUT44), .B(n495), .Z(n496) );
  XNOR2_X1 U561 ( .A(G106GAT), .B(n496), .ZN(G1339GAT) );
  XNOR2_X1 U562 ( .A(G113GAT), .B(KEYINPUT114), .ZN(n516) );
  NAND2_X1 U563 ( .A1(n568), .A2(n533), .ZN(n497) );
  XOR2_X1 U564 ( .A(KEYINPUT46), .B(n497), .Z(n498) );
  NOR2_X1 U565 ( .A1(n560), .A2(n498), .ZN(n499) );
  NAND2_X1 U566 ( .A1(n501), .A2(n499), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n500), .B(KEYINPUT47), .ZN(n508) );
  INV_X1 U568 ( .A(n501), .ZN(n575) );
  NAND2_X1 U569 ( .A1(n575), .A2(n578), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n502), .B(KEYINPUT45), .ZN(n503) );
  XNOR2_X1 U571 ( .A(KEYINPUT65), .B(n503), .ZN(n505) );
  NAND2_X1 U572 ( .A1(n505), .A2(n504), .ZN(n506) );
  NOR2_X1 U573 ( .A1(n506), .A2(n568), .ZN(n507) );
  NOR2_X1 U574 ( .A1(n508), .A2(n507), .ZN(n511) );
  XOR2_X1 U575 ( .A(KEYINPUT64), .B(KEYINPUT113), .Z(n509) );
  XNOR2_X1 U576 ( .A(KEYINPUT48), .B(n509), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(n543) );
  INV_X1 U578 ( .A(n543), .ZN(n528) );
  NAND2_X1 U579 ( .A1(n512), .A2(n528), .ZN(n513) );
  NOR2_X1 U580 ( .A1(n514), .A2(n513), .ZN(n523) );
  NAND2_X1 U581 ( .A1(n568), .A2(n523), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(G1340GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT115), .B(KEYINPUT49), .Z(n518) );
  NAND2_X1 U584 ( .A1(n523), .A2(n554), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U586 ( .A(G120GAT), .B(n519), .Z(G1341GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n521) );
  NAND2_X1 U588 ( .A1(n523), .A2(n575), .ZN(n520) );
  XNOR2_X1 U589 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U590 ( .A(G127GAT), .B(n522), .Z(G1342GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n525) );
  NAND2_X1 U592 ( .A1(n523), .A2(n560), .ZN(n524) );
  XNOR2_X1 U593 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U594 ( .A(G134GAT), .B(n526), .Z(G1343GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n531) );
  NAND2_X1 U596 ( .A1(n527), .A2(n528), .ZN(n529) );
  NOR2_X1 U597 ( .A1(n567), .A2(n529), .ZN(n539) );
  NAND2_X1 U598 ( .A1(n539), .A2(n568), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(n532) );
  XNOR2_X1 U600 ( .A(G141GAT), .B(n532), .ZN(G1344GAT) );
  XNOR2_X1 U601 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n537) );
  XOR2_X1 U602 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n535) );
  NAND2_X1 U603 ( .A1(n539), .A2(n533), .ZN(n534) );
  XNOR2_X1 U604 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(G1345GAT) );
  NAND2_X1 U606 ( .A1(n575), .A2(n539), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n538), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U608 ( .A1(n560), .A2(n539), .ZN(n540) );
  XNOR2_X1 U609 ( .A(n540), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n552) );
  XNOR2_X1 U611 ( .A(KEYINPUT121), .B(n541), .ZN(n542) );
  NOR2_X1 U612 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n544), .B(KEYINPUT54), .ZN(n546) );
  NAND2_X1 U614 ( .A1(n546), .A2(n545), .ZN(n566) );
  NOR2_X1 U615 ( .A1(n547), .A2(n566), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n548), .B(KEYINPUT55), .ZN(n549) );
  NAND2_X1 U617 ( .A1(n561), .A2(n568), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G169GAT), .B(n553), .ZN(G1348GAT) );
  XNOR2_X1 U620 ( .A(KEYINPUT124), .B(KEYINPUT57), .ZN(n558) );
  XOR2_X1 U621 ( .A(G176GAT), .B(KEYINPUT56), .Z(n556) );
  NAND2_X1 U622 ( .A1(n561), .A2(n554), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1349GAT) );
  NAND2_X1 U625 ( .A1(n575), .A2(n561), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U627 ( .A(G190GAT), .B(KEYINPUT125), .ZN(n565) );
  XOR2_X1 U628 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n563) );
  NAND2_X1 U629 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(G1351GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n570) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n579) );
  NAND2_X1 U634 ( .A1(n579), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n574) );
  NAND2_X1 U638 ( .A1(n579), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  XOR2_X1 U640 ( .A(G211GAT), .B(KEYINPUT127), .Z(n577) );
  NAND2_X1 U641 ( .A1(n579), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1354GAT) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U644 ( .A(n580), .B(KEYINPUT62), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

