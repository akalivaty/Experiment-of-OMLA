//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:08 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1204, new_n1205, new_n1206,
    new_n1208, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1273, new_n1274;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G116), .A2(G270), .ZN(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  INV_X1    g0007(.A(G244), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G68), .ZN(new_n214));
  INV_X1    g0014(.A(G238), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n202), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI211_X1 g0016(.A(new_n211), .B(new_n216), .C1(G97), .C2(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G1), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT1), .Z(new_n222));
  OAI21_X1  g0022(.A(G50), .B1(G58), .B2(G68), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR3_X1   g0024(.A1(new_n223), .A2(new_n219), .A3(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(G13), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n220), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n222), .A2(new_n225), .A3(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT65), .B(G107), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND2_X1  g0048(.A1(new_n203), .A2(G20), .ZN(new_n249));
  INV_X1    g0049(.A(G150), .ZN(new_n250));
  NOR2_X1   g0050(.A1(G20), .A2(G33), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  INV_X1    g0053(.A(G33), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(G20), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n249), .B1(new_n250), .B2(new_n252), .C1(new_n253), .C2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  AND3_X1   g0058(.A1(new_n258), .A2(KEYINPUT66), .A3(new_n224), .ZN(new_n259));
  AOI21_X1  g0059(.A(KEYINPUT66), .B1(new_n258), .B2(new_n224), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n218), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  AOI22_X1  g0063(.A1(new_n257), .A2(new_n261), .B1(new_n202), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n261), .A2(new_n263), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n218), .A2(G20), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(G50), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT9), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G222), .ZN(new_n273));
  INV_X1    g0073(.A(G223), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n271), .B(new_n273), .C1(new_n274), .C2(new_n272), .ZN(new_n275));
  AND2_X1   g0075(.A1(G33), .A2(G41), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(new_n224), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n275), .B(new_n277), .C1(G77), .C2(new_n271), .ZN(new_n278));
  INV_X1    g0078(.A(G41), .ZN(new_n279));
  OAI211_X1 g0079(.A(G1), .B(G13), .C1(new_n254), .C2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n218), .B1(G41), .B2(G45), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G226), .ZN(new_n284));
  INV_X1    g0084(.A(G274), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n278), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G190), .ZN(new_n289));
  OR2_X1    g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(G200), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n264), .A2(KEYINPUT9), .A3(new_n267), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n270), .A2(new_n290), .A3(new_n291), .A4(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT10), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n293), .B(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n288), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n297), .B(new_n268), .C1(G179), .C2(new_n288), .ZN(new_n298));
  XNOR2_X1  g0098(.A(new_n298), .B(KEYINPUT67), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT69), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n262), .A2(G77), .ZN(new_n301));
  INV_X1    g0101(.A(new_n253), .ZN(new_n302));
  XOR2_X1   g0102(.A(KEYINPUT15), .B(G87), .Z(new_n303));
  AOI22_X1  g0103(.A1(new_n302), .A2(new_n251), .B1(new_n303), .B2(new_n255), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(new_n219), .B2(new_n207), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n258), .A2(new_n224), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n301), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n306), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n266), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n307), .B1(new_n207), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n272), .A2(G232), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n271), .B(new_n312), .C1(new_n215), .C2(new_n272), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n313), .B(new_n277), .C1(G107), .C2(new_n271), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n283), .A2(G244), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(new_n287), .A3(new_n315), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n316), .A2(KEYINPUT68), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(KEYINPUT68), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G200), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n311), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n289), .B1(new_n317), .B2(new_n318), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n317), .A2(new_n318), .A3(new_n296), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n310), .ZN(new_n325));
  AOI21_X1  g0125(.A(G179), .B1(new_n317), .B2(new_n318), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n300), .B1(new_n323), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n319), .A2(G190), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n329), .B(new_n311), .C1(new_n320), .C2(new_n319), .ZN(new_n330));
  INV_X1    g0130(.A(new_n326), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(new_n310), .A3(new_n324), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n330), .A2(new_n332), .A3(KEYINPUT69), .ZN(new_n333));
  AOI211_X1 g0133(.A(new_n295), .B(new_n299), .C1(new_n328), .C2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(G58), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n335), .A2(new_n214), .ZN(new_n336));
  OAI21_X1  g0136(.A(G20), .B1(new_n336), .B2(new_n201), .ZN(new_n337));
  INV_X1    g0137(.A(G159), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n337), .B1(new_n338), .B2(new_n252), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT7), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n340), .B1(new_n271), .B2(G20), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT3), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G33), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n340), .A2(G20), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n339), .B1(new_n348), .B2(G68), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n308), .B1(new_n349), .B2(KEYINPUT16), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT75), .ZN(new_n351));
  OAI21_X1  g0151(.A(new_n351), .B1(new_n254), .B2(KEYINPUT3), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n342), .A2(KEYINPUT75), .A3(G33), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n352), .A2(new_n344), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n346), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT76), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n354), .A2(KEYINPUT76), .A3(new_n346), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n357), .A2(new_n341), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n339), .B1(new_n359), .B2(G68), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n350), .B1(new_n360), .B2(KEYINPUT16), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n213), .A2(G1698), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n274), .A2(new_n272), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n271), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(G33), .A2(G87), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n280), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n280), .A2(G232), .A3(new_n281), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n366), .A2(new_n286), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n289), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n368), .B2(G200), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n253), .B1(new_n218), .B2(G20), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n265), .A2(new_n371), .B1(new_n263), .B2(new_n253), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n361), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  XNOR2_X1  g0173(.A(KEYINPUT77), .B(KEYINPUT17), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n373), .A2(new_n375), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n361), .A2(new_n372), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n364), .A2(new_n365), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n286), .B1(new_n379), .B2(new_n277), .ZN(new_n380));
  INV_X1    g0180(.A(new_n367), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n296), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G179), .ZN(new_n383));
  NOR4_X1   g0183(.A1(new_n366), .A2(new_n383), .A3(new_n367), .A4(new_n286), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT18), .B1(new_n378), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT18), .ZN(new_n388));
  AOI211_X1 g0188(.A(new_n388), .B(new_n385), .C1(new_n361), .C2(new_n372), .ZN(new_n389));
  OAI22_X1  g0189(.A1(new_n376), .A2(new_n377), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT78), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI221_X1 g0192(.A(KEYINPUT78), .B1(new_n387), .B2(new_n389), .C1(new_n377), .C2(new_n376), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT13), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n343), .A2(new_n344), .A3(G226), .A4(new_n272), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT70), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n271), .A2(KEYINPUT70), .A3(G226), .A4(new_n272), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G33), .A2(G97), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT71), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(KEYINPUT71), .A2(G33), .A3(G97), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  AND4_X1   g0206(.A1(G232), .A2(new_n343), .A3(new_n344), .A4(G1698), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n400), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n286), .B1(new_n409), .B2(new_n277), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n282), .A2(new_n215), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n395), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n407), .B1(new_n398), .B2(new_n399), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n280), .B1(new_n414), .B2(new_n406), .ZN(new_n415));
  NOR4_X1   g0215(.A1(new_n415), .A2(KEYINPUT13), .A3(new_n286), .A4(new_n411), .ZN(new_n416));
  OAI21_X1  g0216(.A(G169), .B1(new_n413), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT14), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n413), .A2(new_n416), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G179), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT14), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n421), .B(G169), .C1(new_n413), .C2(new_n416), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n418), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT74), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n256), .A2(new_n207), .B1(new_n219), .B2(G68), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n252), .A2(new_n202), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n261), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  XNOR2_X1  g0228(.A(KEYINPUT72), .B(KEYINPUT11), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n263), .A2(KEYINPUT73), .A3(new_n214), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT12), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT73), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n262), .B2(G68), .ZN(new_n434));
  XOR2_X1   g0234(.A(new_n432), .B(new_n434), .Z(new_n435));
  NOR2_X1   g0235(.A1(new_n309), .A2(new_n214), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n430), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n418), .A2(KEYINPUT74), .A3(new_n420), .A4(new_n422), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n425), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n438), .B1(new_n419), .B2(G190), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n320), .B2(new_n419), .ZN(new_n442));
  AND4_X1   g0242(.A1(new_n334), .A2(new_n394), .A3(new_n440), .A4(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT4), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n444), .B1(new_n345), .B2(new_n208), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(G1698), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n271), .A2(G244), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G33), .A2(G283), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n445), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n271), .A2(G250), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n272), .B1(new_n450), .B2(KEYINPUT4), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n277), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(G45), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n453), .A2(G1), .ZN(new_n454));
  NOR2_X1   g0254(.A1(KEYINPUT5), .A2(G41), .ZN(new_n455));
  AND2_X1   g0255(.A1(KEYINPUT5), .A2(G41), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n454), .B(G274), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n454), .B1(new_n456), .B2(new_n455), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n280), .ZN(new_n459));
  INV_X1    g0259(.A(G257), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT81), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT81), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n463), .B(new_n457), .C1(new_n459), .C2(new_n460), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n452), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n296), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n452), .A2(new_n462), .A3(new_n383), .A4(new_n464), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n359), .A2(G107), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT6), .ZN(new_n469));
  AND2_X1   g0269(.A1(G97), .A2(G107), .ZN(new_n470));
  NOR2_X1   g0270(.A1(G97), .A2(G107), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G107), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n473), .A2(KEYINPUT6), .A3(G97), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n219), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n252), .A2(new_n207), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT79), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT79), .ZN(new_n478));
  INV_X1    g0278(.A(new_n476), .ZN(new_n479));
  AND3_X1   g0279(.A1(new_n473), .A2(KEYINPUT6), .A3(G97), .ZN(new_n480));
  XNOR2_X1  g0280(.A(G97), .B(G107), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n480), .B1(new_n481), .B2(new_n469), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n478), .B(new_n479), .C1(new_n482), .C2(new_n219), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n308), .B1(new_n468), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n263), .A2(G97), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n218), .A2(G33), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n262), .B(new_n487), .C1(new_n259), .C2(new_n260), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n486), .B1(new_n488), .B2(G97), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT80), .ZN(new_n490));
  XNOR2_X1  g0290(.A(new_n489), .B(new_n490), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n466), .B(new_n467), .C1(new_n485), .C2(new_n491), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n354), .A2(KEYINPUT76), .A3(new_n346), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT76), .B1(new_n354), .B2(new_n346), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n473), .B1(new_n495), .B2(new_n341), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n477), .A2(new_n483), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n306), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n465), .A2(G200), .ZN(new_n499));
  XNOR2_X1  g0299(.A(new_n489), .B(KEYINPUT80), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n452), .A2(new_n462), .A3(G190), .A4(new_n464), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n498), .A2(new_n499), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n492), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT82), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT82), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n492), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(new_n488), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n303), .ZN(new_n509));
  INV_X1    g0309(.A(new_n303), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n263), .ZN(new_n511));
  NOR3_X1   g0311(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n512));
  AND3_X1   g0312(.A1(KEYINPUT71), .A2(G33), .A3(G97), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT71), .B1(G33), .B2(G97), .ZN(new_n514));
  OAI21_X1  g0314(.A(KEYINPUT19), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n512), .B1(new_n515), .B2(new_n219), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n345), .A2(G20), .A3(new_n214), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT19), .B1(new_n255), .B2(G97), .ZN(new_n518));
  NOR3_X1   g0318(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n509), .B(new_n511), .C1(new_n519), .C2(new_n308), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n454), .A2(G274), .ZN(new_n521));
  NOR2_X1   g0321(.A1(G238), .A2(G1698), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n208), .B2(G1698), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n523), .A2(new_n271), .B1(G33), .B2(G116), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n521), .B1(new_n524), .B2(new_n280), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n218), .A2(G45), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n526), .B(G250), .C1(new_n276), .C2(new_n224), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT83), .ZN(new_n528));
  XNOR2_X1  g0328(.A(new_n527), .B(new_n528), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n296), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g0330(.A(new_n527), .B(KEYINPUT83), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n208), .A2(G1698), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(G238), .B2(G1698), .ZN(new_n533));
  INV_X1    g0333(.A(G116), .ZN(new_n534));
  OAI22_X1  g0334(.A1(new_n533), .A2(new_n345), .B1(new_n254), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n277), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n531), .A2(new_n536), .A3(new_n383), .A4(new_n521), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n520), .A2(new_n530), .A3(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n271), .A2(new_n219), .A3(G68), .ZN(new_n539));
  INV_X1    g0339(.A(new_n518), .ZN(new_n540));
  AOI21_X1  g0340(.A(G20), .B1(new_n405), .B2(KEYINPUT19), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n539), .B(new_n540), .C1(new_n541), .C2(new_n512), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n542), .A2(new_n306), .B1(new_n263), .B2(new_n510), .ZN(new_n543));
  OAI21_X1  g0343(.A(G200), .B1(new_n525), .B2(new_n529), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n508), .A2(G87), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n531), .A2(new_n536), .A3(G190), .A4(new_n521), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n543), .A2(new_n544), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n538), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n343), .A2(new_n344), .A3(new_n219), .A4(G87), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT22), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT22), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n271), .A2(new_n551), .A3(new_n219), .A4(G87), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(KEYINPUT87), .A2(KEYINPUT23), .A3(G107), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT87), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(G20), .B2(new_n473), .ZN(new_n556));
  AOI22_X1  g0356(.A1(KEYINPUT87), .A2(KEYINPUT23), .B1(G33), .B2(G116), .ZN(new_n557));
  OAI22_X1  g0357(.A1(new_n556), .A2(KEYINPUT23), .B1(new_n557), .B2(G20), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n553), .A2(new_n554), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(KEYINPUT24), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n558), .B1(new_n550), .B2(new_n552), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT24), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n562), .A2(new_n563), .A3(new_n554), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n308), .B1(new_n561), .B2(new_n564), .ZN(new_n565));
  NOR4_X1   g0365(.A1(new_n226), .A2(new_n219), .A3(G1), .A4(G107), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT25), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n508), .A2(G107), .B1(new_n567), .B2(new_n566), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n565), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n210), .A2(new_n272), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n460), .A2(G1698), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n343), .A2(new_n572), .A3(new_n344), .A4(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(G294), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT88), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT88), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G294), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n578), .A3(G33), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n277), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n458), .A2(G264), .A3(new_n280), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n457), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT89), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n583), .A2(new_n584), .A3(G169), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n584), .B1(new_n583), .B2(G169), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n583), .A2(new_n383), .ZN(new_n587));
  NOR3_X1   g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AND3_X1   g0388(.A1(new_n562), .A2(new_n563), .A3(new_n554), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n563), .B1(new_n562), .B2(new_n554), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n306), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n568), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n583), .A2(G200), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n569), .A4(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n583), .A2(new_n289), .ZN(new_n595));
  OAI22_X1  g0395(.A1(new_n571), .A2(new_n588), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(G303), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n342), .A2(G33), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n272), .A2(G257), .ZN(new_n601));
  NAND2_X1  g0401(.A1(G264), .A2(G1698), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n343), .A2(new_n344), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n603), .A3(new_n277), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n458), .A2(G270), .A3(new_n280), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n604), .A2(new_n457), .A3(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT84), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n604), .A2(KEYINPUT84), .A3(new_n457), .A4(new_n605), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n608), .A2(G169), .A3(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT86), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n263), .A2(KEYINPUT85), .A3(new_n534), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT85), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n262), .B2(G116), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n308), .A2(G116), .A3(new_n262), .A4(new_n487), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n258), .A2(new_n224), .B1(G20), .B2(new_n534), .ZN(new_n617));
  INV_X1    g0417(.A(G97), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n448), .B(new_n219), .C1(G33), .C2(new_n618), .ZN(new_n619));
  AND3_X1   g0419(.A1(new_n617), .A2(KEYINPUT20), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT20), .B1(new_n617), .B2(new_n619), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n615), .B(new_n616), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n610), .A2(new_n611), .A3(KEYINPUT21), .A4(new_n622), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n608), .A2(G169), .A3(new_n622), .A4(new_n609), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT21), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(KEYINPUT86), .B1(new_n624), .B2(new_n625), .ZN(new_n627));
  OR2_X1    g0427(.A1(new_n606), .A2(new_n383), .ZN(new_n628));
  INV_X1    g0428(.A(new_n622), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n623), .A2(new_n626), .A3(new_n627), .A4(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n289), .B1(new_n608), .B2(new_n609), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n608), .A2(new_n609), .ZN(new_n633));
  AOI211_X1 g0433(.A(new_n622), .B(new_n632), .C1(new_n633), .C2(G200), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n596), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  AND4_X1   g0435(.A1(new_n443), .A2(new_n507), .A3(new_n548), .A4(new_n635), .ZN(G372));
  AND3_X1   g0436(.A1(new_n623), .A2(new_n627), .A3(new_n630), .ZN(new_n637));
  INV_X1    g0437(.A(new_n588), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n591), .A2(new_n592), .A3(new_n569), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT90), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n637), .A2(new_n640), .A3(new_n641), .A4(new_n626), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n548), .A2(new_n492), .A3(new_n502), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n594), .A2(new_n595), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n571), .A2(new_n588), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT90), .B1(new_n646), .B2(new_n631), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n642), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n538), .ZN(new_n649));
  AOI22_X1  g0449(.A1(new_n498), .A2(new_n500), .B1(new_n296), .B2(new_n465), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n548), .A2(new_n650), .A3(KEYINPUT26), .A4(new_n467), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT26), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n538), .A2(new_n547), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n652), .B1(new_n492), .B2(new_n653), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n649), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n648), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n443), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n299), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT91), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n295), .B(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n376), .A2(new_n377), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n442), .A2(new_n327), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n661), .B1(new_n440), .B2(new_n662), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n387), .A2(new_n389), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n660), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n657), .A2(new_n658), .A3(new_n666), .ZN(G369));
  NOR2_X1   g0467(.A1(new_n565), .A2(new_n570), .ZN(new_n668));
  INV_X1    g0468(.A(new_n595), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n668), .A2(new_n592), .A3(new_n669), .A4(new_n593), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n218), .A2(new_n219), .A3(G13), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT92), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n671), .B(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT93), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n676), .A2(G213), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(G343), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  OAI211_X1 g0481(.A(new_n640), .B(new_n670), .C1(new_n571), .C2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT94), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n682), .B(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n631), .A2(new_n681), .ZN(new_n685));
  OR2_X1    g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n640), .B2(new_n680), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n646), .A2(new_n680), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n631), .A2(new_n634), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n680), .A2(new_n622), .ZN(new_n692));
  MUX2_X1   g0492(.A(new_n631), .B(new_n691), .S(new_n692), .Z(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(G330), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n687), .A2(new_n695), .ZN(G399));
  NOR2_X1   g0496(.A1(new_n227), .A2(G41), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G1), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n512), .A2(new_n534), .ZN(new_n700));
  OAI22_X1  g0500(.A1(new_n699), .A2(new_n700), .B1(new_n223), .B2(new_n698), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT28), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n680), .B1(new_n648), .B2(new_n655), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT29), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n651), .A2(KEYINPUT97), .A3(new_n654), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT97), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n707), .B(new_n652), .C1(new_n492), .C2(new_n653), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n538), .A2(KEYINPUT96), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n646), .A2(new_n631), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n670), .A2(new_n492), .A3(new_n502), .A4(new_n548), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n538), .A2(KEYINPUT96), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n680), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n705), .B1(new_n716), .B2(new_n704), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n628), .A2(new_n525), .A3(new_n529), .ZN(new_n718));
  INV_X1    g0518(.A(new_n465), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n718), .A2(new_n719), .A3(new_n581), .A4(new_n582), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n525), .ZN(new_n723));
  AOI21_X1  g0523(.A(G179), .B1(new_n723), .B2(new_n531), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n633), .A2(new_n724), .A3(new_n465), .A4(new_n583), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  OR2_X1    g0527(.A1(new_n720), .A2(new_n721), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n681), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n635), .A2(new_n507), .A3(new_n548), .A4(new_n681), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(new_n730), .B2(KEYINPUT31), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT95), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n726), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n722), .A2(KEYINPUT95), .A3(new_n725), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(new_n728), .A3(new_n734), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n735), .A2(KEYINPUT31), .A3(new_n680), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n717), .B1(G330), .B2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n702), .B1(new_n738), .B2(G1), .ZN(G364));
  NOR2_X1   g0539(.A1(new_n219), .A2(new_n383), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G190), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(new_n320), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G326), .ZN(new_n743));
  INV_X1    g0543(.A(G283), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n219), .A2(G190), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n320), .A2(G179), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n743), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n740), .A2(new_n289), .A3(G200), .ZN(new_n749));
  INV_X1    g0549(.A(G317), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n749), .B1(KEYINPUT33), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(KEYINPUT33), .B2(new_n750), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n740), .A2(new_n289), .A3(new_n320), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n271), .B1(new_n754), .B2(G311), .ZN(new_n755));
  INV_X1    g0555(.A(G322), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n741), .A2(G200), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n752), .B(new_n755), .C1(new_n756), .C2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT100), .ZN(new_n760));
  INV_X1    g0560(.A(new_n745), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n383), .A2(new_n320), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n760), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n745), .A2(KEYINPUT100), .A3(new_n383), .A4(new_n320), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n748), .B(new_n759), .C1(G329), .C2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n746), .A2(G20), .A3(G190), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n576), .A2(new_n578), .ZN(new_n769));
  OAI21_X1  g0569(.A(G20), .B1(new_n762), .B2(new_n289), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT101), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n767), .B1(new_n597), .B2(new_n768), .C1(new_n769), .C2(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(G58), .A2(new_n757), .B1(new_n754), .B2(G77), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(KEYINPUT99), .ZN(new_n777));
  INV_X1    g0577(.A(new_n742), .ZN(new_n778));
  OAI221_X1 g0578(.A(new_n271), .B1(new_n747), .B2(new_n473), .C1(new_n778), .C2(new_n202), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(KEYINPUT99), .B2(new_n776), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n765), .A2(new_n338), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT32), .ZN(new_n782));
  INV_X1    g0582(.A(new_n774), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G97), .ZN(new_n784));
  INV_X1    g0584(.A(new_n749), .ZN(new_n785));
  INV_X1    g0585(.A(new_n768), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G68), .A2(new_n785), .B1(new_n786), .B2(G87), .ZN(new_n787));
  NAND4_X1  g0587(.A1(new_n780), .A2(new_n782), .A3(new_n784), .A4(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n775), .B1(new_n777), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n224), .B1(G20), .B2(new_n296), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  XOR2_X1   g0591(.A(new_n791), .B(KEYINPUT98), .Z(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(G20), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n790), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n227), .A2(new_n271), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n223), .A2(G45), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n796), .B(new_n797), .C1(new_n247), .C2(new_n453), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n228), .A2(G355), .A3(new_n271), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n798), .B(new_n799), .C1(G116), .C2(new_n228), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n789), .A2(new_n790), .B1(new_n795), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n226), .A2(G20), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n699), .B1(G45), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n794), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n801), .B(new_n803), .C1(new_n693), .C2(new_n804), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT102), .Z(new_n806));
  NOR2_X1   g0606(.A1(new_n693), .A2(G330), .ZN(new_n807));
  INV_X1    g0607(.A(new_n803), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n694), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n806), .B1(new_n807), .B2(new_n809), .ZN(G396));
  NAND2_X1  g0610(.A1(new_n737), .A2(G330), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n332), .A2(new_n680), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n330), .B1(new_n311), .B2(new_n681), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n812), .B1(new_n813), .B2(new_n332), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n703), .B(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n808), .B1(new_n811), .B2(new_n815), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT103), .Z(new_n817));
  NAND2_X1  g0617(.A1(new_n811), .A2(new_n815), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G143), .A2(new_n757), .B1(new_n785), .B2(G150), .ZN(new_n820));
  INV_X1    g0620(.A(G137), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n820), .B1(new_n821), .B2(new_n778), .C1(new_n338), .C2(new_n753), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT34), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(G132), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n824), .B1(new_n214), .B2(new_n747), .C1(new_n825), .C2(new_n765), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n345), .B1(new_n786), .B2(G50), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n827), .B1(new_n335), .B2(new_n774), .C1(new_n822), .C2(new_n823), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n345), .B1(new_n753), .B2(new_n534), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(G283), .B2(new_n785), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n830), .B1(new_n209), .B2(new_n747), .C1(new_n473), .C2(new_n768), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n766), .A2(G311), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G294), .A2(new_n757), .B1(new_n742), .B2(G303), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n784), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n826), .A2(new_n828), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n790), .A2(new_n791), .ZN(new_n836));
  AOI22_X1  g0636(.A1(new_n835), .A2(new_n790), .B1(new_n207), .B2(new_n836), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n803), .B(new_n837), .C1(new_n814), .C2(new_n793), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n819), .A2(new_n838), .ZN(G384));
  INV_X1    g0639(.A(KEYINPUT40), .ZN(new_n840));
  INV_X1    g0640(.A(new_n814), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n730), .A2(KEYINPUT31), .ZN(new_n842));
  INV_X1    g0642(.A(new_n729), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n729), .A2(KEYINPUT31), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n841), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n440), .A2(new_n442), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n681), .A2(new_n437), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n848), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n440), .A2(new_n442), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n846), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n678), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n349), .A2(KEYINPUT16), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n261), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n349), .A2(KEYINPUT16), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n372), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n390), .A2(new_n854), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n858), .B1(new_n854), .B2(new_n386), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n373), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n378), .A2(new_n386), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n378), .A2(new_n854), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n864), .A3(new_n373), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n862), .B1(KEYINPUT37), .B2(new_n865), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n859), .A2(KEYINPUT38), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT38), .B1(new_n859), .B2(new_n866), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n840), .B1(new_n853), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n859), .A2(KEYINPUT38), .A3(new_n866), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT107), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n865), .B(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n864), .B1(new_n664), .B2(KEYINPUT17), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT107), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n859), .A2(new_n878), .A3(KEYINPUT38), .A4(new_n866), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n872), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  NAND4_X1  g0680(.A1(new_n846), .A2(new_n880), .A3(KEYINPUT40), .A4(new_n852), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n870), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n844), .A2(new_n845), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n443), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n882), .B(new_n884), .Z(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(G330), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n440), .A2(new_n680), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT39), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n872), .A2(new_n888), .A3(new_n877), .A4(new_n879), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT106), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n890), .B(KEYINPUT39), .C1(new_n867), .C2(new_n868), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n859), .A2(new_n866), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n873), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n871), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n890), .B1(new_n895), .B2(KEYINPUT39), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n887), .B1(new_n892), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n703), .A2(new_n814), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT105), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n812), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n812), .A2(new_n899), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n898), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(new_n852), .A3(new_n895), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n665), .A2(new_n678), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n897), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n666), .A2(new_n658), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n717), .B2(new_n443), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n906), .B(new_n908), .Z(new_n909));
  XNOR2_X1  g0709(.A(new_n886), .B(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n218), .B2(new_n802), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT35), .ZN(new_n912));
  AOI211_X1 g0712(.A(new_n219), .B(new_n224), .C1(new_n482), .C2(new_n912), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n913), .B(G116), .C1(new_n912), .C2(new_n482), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT36), .ZN(new_n915));
  OAI21_X1  g0715(.A(G77), .B1(new_n335), .B2(new_n214), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n916), .A2(new_n223), .B1(G50), .B2(new_n214), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(G1), .A3(new_n226), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT104), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n911), .A2(new_n915), .A3(new_n919), .ZN(G367));
  OAI21_X1  g0720(.A(new_n680), .B1(new_n485), .B2(new_n491), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(new_n492), .A3(new_n502), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n686), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT42), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n492), .B1(new_n922), .B2(new_n640), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n681), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT108), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT43), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n543), .A2(new_n545), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n680), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n548), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n538), .B2(new_n931), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n929), .A2(new_n933), .A3(new_n927), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n933), .B2(new_n929), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n650), .A2(new_n467), .A3(new_n680), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n922), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n690), .A2(new_n694), .A3(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n935), .B(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n218), .B1(new_n802), .B2(G45), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n697), .B(KEYINPUT41), .Z(new_n943));
  NAND2_X1  g0743(.A1(new_n687), .A2(new_n938), .ZN(new_n944));
  XOR2_X1   g0744(.A(new_n944), .B(KEYINPUT44), .Z(new_n945));
  NAND2_X1  g0745(.A1(new_n695), .A2(KEYINPUT110), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n687), .A2(new_n938), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT45), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n695), .A2(KEYINPUT110), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n949), .B(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n685), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n686), .B1(new_n689), .B2(new_n952), .ZN(new_n953));
  XOR2_X1   g0753(.A(new_n953), .B(new_n694), .Z(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n738), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT109), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n951), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n943), .B1(new_n957), .B2(new_n738), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n940), .B1(new_n942), .B2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT111), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n768), .B2(new_n534), .ZN(new_n961));
  OR2_X1    g0761(.A1(new_n961), .A2(KEYINPUT46), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(KEYINPUT46), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n962), .B(new_n963), .C1(new_n750), .C2(new_n765), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n747), .A2(new_n618), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n271), .B(new_n965), .C1(G311), .C2(new_n742), .ZN(new_n966));
  INV_X1    g0766(.A(new_n769), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n967), .A2(new_n785), .B1(new_n754), .B2(G283), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n966), .B(new_n968), .C1(new_n473), .C2(new_n774), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n964), .B(new_n969), .C1(G303), .C2(new_n757), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n786), .A2(G58), .ZN(new_n971));
  AOI22_X1  g0771(.A1(G143), .A2(new_n742), .B1(new_n757), .B2(G150), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n821), .B2(new_n765), .ZN(new_n973));
  INV_X1    g0773(.A(new_n747), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n345), .B1(new_n974), .B2(G77), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n975), .B1(new_n202), .B2(new_n753), .C1(new_n338), .C2(new_n749), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n774), .A2(new_n214), .ZN(new_n977));
  NOR3_X1   g0777(.A1(new_n973), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n970), .B1(new_n971), .B2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT47), .Z(new_n980));
  AOI21_X1  g0780(.A(new_n808), .B1(new_n980), .B2(new_n790), .ZN(new_n981));
  INV_X1    g0781(.A(new_n796), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n795), .B1(new_n228), .B2(new_n510), .C1(new_n239), .C2(new_n982), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n981), .B(new_n983), .C1(new_n804), .C2(new_n933), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n959), .A2(new_n984), .ZN(G387));
  XOR2_X1   g0785(.A(new_n697), .B(KEYINPUT115), .Z(new_n986));
  NOR2_X1   g0786(.A1(new_n954), .A2(new_n738), .ZN(new_n987));
  OR3_X1    g0787(.A1(new_n956), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n954), .A2(new_n942), .ZN(new_n989));
  AND2_X1   g0789(.A1(new_n766), .A2(G326), .ZN(new_n990));
  AOI22_X1  g0790(.A1(G317), .A2(new_n757), .B1(new_n785), .B2(G311), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n597), .B2(new_n753), .C1(new_n756), .C2(new_n778), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n994));
  AOI22_X1  g0794(.A1(new_n993), .A2(new_n994), .B1(G283), .B2(new_n783), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n769), .B2(new_n768), .C1(new_n994), .C2(new_n993), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT49), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n271), .B(new_n990), .C1(new_n996), .C2(new_n997), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n997), .B2(new_n996), .C1(new_n534), .C2(new_n747), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n783), .A2(new_n303), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n202), .B2(new_n758), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT113), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n253), .A2(new_n749), .B1(new_n753), .B2(new_n214), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n768), .A2(new_n207), .ZN(new_n1004));
  OR3_X1    g0804(.A1(new_n1004), .A2(new_n965), .A3(new_n345), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(KEYINPUT112), .B(G150), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1003), .B(new_n1005), .C1(new_n766), .C2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1002), .B(new_n1007), .C1(new_n338), .C2(new_n778), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n999), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n790), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n302), .A2(new_n202), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n700), .B1(new_n1011), .B2(KEYINPUT50), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1012), .B(new_n453), .C1(KEYINPUT50), .C2(new_n1011), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(G68), .B2(G77), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n796), .B1(new_n236), .B2(new_n453), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n228), .A2(new_n271), .A3(new_n700), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n228), .A2(G107), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n795), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1010), .B(new_n1019), .C1(new_n689), .C2(new_n804), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n988), .B(new_n989), .C1(new_n808), .C2(new_n1020), .ZN(G393));
  NAND2_X1  g0821(.A1(new_n951), .A2(new_n942), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(G150), .A2(new_n742), .B1(new_n757), .B2(G159), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1023), .B(KEYINPUT51), .Z(new_n1024));
  OAI21_X1  g0824(.A(new_n271), .B1(new_n768), .B2(new_n214), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n766), .B2(G143), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n783), .A2(G77), .B1(G87), .B2(new_n974), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n202), .A2(new_n749), .B1(new_n753), .B2(new_n253), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT116), .Z(new_n1029));
  NAND4_X1  g0829(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G311), .A2(new_n757), .B1(new_n742), .B2(G317), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n1031), .A2(KEYINPUT52), .B1(new_n756), .B2(new_n765), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(KEYINPUT52), .B2(new_n1031), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n473), .B2(new_n747), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n575), .A2(new_n753), .B1(new_n749), .B2(new_n597), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(G283), .B2(new_n786), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1036), .B(new_n345), .C1(new_n534), .C2(new_n774), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1030), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n808), .B1(new_n1038), .B2(new_n790), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n795), .B1(new_n618), .B2(new_n228), .C1(new_n244), .C2(new_n982), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(new_n937), .C2(new_n804), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1022), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n986), .B1(new_n951), .B2(new_n956), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n951), .A2(new_n956), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1042), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(G390));
  OAI21_X1  g0847(.A(new_n271), .B1(new_n758), .B2(new_n825), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n742), .A2(G128), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n747), .A2(new_n202), .ZN(new_n1050));
  XOR2_X1   g0850(.A(KEYINPUT54), .B(G143), .Z(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n1052), .A2(new_n753), .B1(new_n821), .B2(new_n749), .ZN(new_n1053));
  NOR4_X1   g0853(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .A4(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(G125), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1054), .B1(new_n1055), .B2(new_n765), .C1(new_n338), .C2(new_n774), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n786), .A2(new_n1006), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1057), .B(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n778), .A2(new_n744), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n753), .A2(new_n618), .B1(new_n768), .B2(new_n209), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n271), .B(new_n1061), .C1(G107), .C2(new_n785), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n783), .A2(G77), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n766), .A2(G294), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n757), .A2(G116), .B1(new_n974), .B2(G68), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n1056), .A2(new_n1059), .B1(new_n1060), .B2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1067), .A2(new_n790), .B1(new_n253), .B2(new_n836), .ZN(new_n1068));
  OAI21_X1  g0868(.A(KEYINPUT39), .B1(new_n867), .B2(new_n868), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(KEYINPUT106), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1070), .A2(new_n889), .A3(new_n891), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n803), .B(new_n1068), .C1(new_n1071), .C2(new_n793), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n887), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n813), .A2(new_n332), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n812), .B1(new_n716), .B2(new_n1074), .ZN(new_n1075));
  AND3_X1   g0875(.A1(new_n440), .A2(new_n442), .A3(new_n850), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n850), .B1(new_n440), .B2(new_n442), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1073), .B(new_n880), .C1(new_n1075), .C2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n887), .B1(new_n903), .B2(new_n852), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1079), .B1(new_n1071), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n846), .A2(G330), .A3(new_n852), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI211_X1 g0883(.A(G330), .B(new_n814), .C1(new_n731), .C2(new_n736), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1084), .A2(new_n1078), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1079), .B(new_n1085), .C1(new_n1071), .C2(new_n1080), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n1087), .A2(KEYINPUT118), .A3(new_n942), .ZN(new_n1088));
  AOI21_X1  g0888(.A(KEYINPUT118), .B1(new_n1087), .B2(new_n942), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1072), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n883), .A2(new_n443), .A3(G330), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT117), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n883), .A2(new_n443), .A3(KEYINPUT117), .A4(G330), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n737), .A2(new_n852), .A3(G330), .A4(new_n814), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n845), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n814), .B1(new_n731), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g0898(.A(G330), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1078), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AND3_X1   g0900(.A1(new_n1096), .A2(new_n1100), .A3(new_n1075), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n902), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n900), .B(new_n1102), .C1(new_n703), .C2(new_n814), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1084), .A2(new_n1078), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1103), .B1(new_n1082), .B2(new_n1104), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n908), .B(new_n1095), .C1(new_n1101), .C2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1107), .A2(new_n1087), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1106), .B1(new_n1083), .B2(new_n1086), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n1108), .A2(new_n1109), .A3(new_n986), .ZN(new_n1110));
  OR2_X1    g0910(.A1(new_n1090), .A2(new_n1110), .ZN(G378));
  NOR3_X1   g0911(.A1(new_n1098), .A2(new_n1078), .A3(new_n869), .ZN(new_n1112));
  OAI211_X1 g0912(.A(G330), .B(new_n881), .C1(new_n1112), .C2(KEYINPUT40), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n854), .A2(new_n268), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n660), .A2(new_n298), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1114), .B1(new_n660), .B2(new_n298), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT121), .B(KEYINPUT56), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT55), .Z(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  OR3_X1    g0919(.A1(new_n1115), .A2(new_n1116), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1119), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1113), .A2(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n870), .A2(G330), .A3(new_n881), .A4(new_n1122), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n906), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n906), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1130), .A2(new_n942), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1123), .A2(new_n792), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n825), .A2(new_n749), .B1(new_n753), .B2(new_n821), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n778), .A2(new_n1055), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1133), .B(new_n1134), .C1(G128), .C2(new_n757), .ZN(new_n1135));
  OAI221_X1 g0935(.A(new_n1135), .B1(new_n250), .B2(new_n774), .C1(new_n768), .C2(new_n1052), .ZN(new_n1136));
  XOR2_X1   g0936(.A(new_n1136), .B(KEYINPUT59), .Z(new_n1137));
  AOI21_X1  g0937(.A(G41), .B1(new_n766), .B2(G124), .ZN(new_n1138));
  AOI21_X1  g0938(.A(G33), .B1(new_n974), .B2(G159), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n279), .B1(new_n342), .B2(new_n254), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n202), .ZN(new_n1142));
  OR2_X1    g0942(.A1(new_n1142), .A2(KEYINPUT120), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n279), .B1(new_n749), .B2(new_n618), .C1(new_n510), .C2(new_n753), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1144), .A2(new_n271), .A3(new_n1004), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n757), .A2(G107), .B1(new_n974), .B2(G58), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n744), .B2(new_n765), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n778), .A2(new_n534), .ZN(new_n1149));
  NOR4_X1   g0949(.A1(new_n1146), .A2(new_n1148), .A3(new_n977), .A4(new_n1149), .ZN(new_n1150));
  OR2_X1    g0950(.A1(new_n1150), .A2(KEYINPUT58), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1150), .A2(KEYINPUT58), .B1(KEYINPUT120), .B2(new_n1142), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1140), .A2(new_n1143), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1153), .A2(new_n790), .B1(new_n202), .B2(new_n836), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1132), .A2(new_n803), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1131), .A2(new_n1155), .ZN(new_n1156));
  AND2_X1   g0956(.A1(new_n1095), .A2(new_n908), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1105), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1096), .A2(new_n1100), .A3(new_n1075), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1086), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1082), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1073), .B1(new_n1103), .B2(new_n1078), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1163), .A2(new_n1070), .A3(new_n889), .A4(new_n891), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1162), .B1(new_n1164), .B2(new_n1079), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1157), .B(new_n1160), .C1(new_n1161), .C2(new_n1165), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1129), .A2(new_n1128), .B1(new_n1166), .B2(new_n1157), .ZN(new_n1167));
  AOI21_X1  g0967(.A(KEYINPUT122), .B1(new_n1167), .B2(KEYINPUT57), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1161), .A2(new_n1165), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1157), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  AND4_X1   g0971(.A1(KEYINPUT122), .A2(new_n1130), .A3(new_n1171), .A4(KEYINPUT57), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1095), .A2(new_n908), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n906), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n906), .B1(new_n1125), .B2(new_n1124), .ZN(new_n1176));
  OAI22_X1  g0976(.A1(new_n1109), .A2(new_n1174), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT57), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n986), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1156), .B1(new_n1173), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(G375));
  NAND2_X1  g0981(.A1(new_n1078), .A2(new_n791), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n766), .A2(G128), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n758), .A2(new_n821), .B1(new_n338), .B2(new_n768), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n271), .B1(new_n1052), .B2(new_n749), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n753), .A2(new_n250), .B1(new_n747), .B2(new_n335), .ZN(new_n1186));
  NOR4_X1   g0986(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .A4(new_n1186), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n202), .B2(new_n774), .C1(new_n825), .C2(new_n778), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n778), .A2(new_n575), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n758), .A2(new_n744), .B1(new_n618), .B2(new_n768), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(new_n766), .B2(G303), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n749), .A2(new_n534), .B1(new_n747), .B2(new_n207), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n271), .B(new_n1192), .C1(G107), .C2(new_n754), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1000), .A3(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1188), .B1(new_n1189), .B2(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1195), .A2(new_n790), .B1(new_n214), .B2(new_n836), .ZN(new_n1196));
  AND3_X1   g0996(.A1(new_n1182), .A2(new_n803), .A3(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(new_n1160), .B2(new_n942), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1170), .A2(new_n1174), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1200), .A2(new_n943), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1198), .B1(new_n1201), .B2(new_n1107), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT123), .Z(G381));
  NOR2_X1   g1003(.A1(G387), .A2(G390), .ZN(new_n1204));
  NOR4_X1   g1004(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(G375), .A2(G378), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .ZN(G407));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n679), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(G407), .A2(G213), .A3(new_n1208), .ZN(G409));
  INV_X1    g1009(.A(KEYINPUT126), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1155), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1130), .B2(new_n942), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n943), .B2(new_n1177), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1090), .A2(new_n1110), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1214), .A2(new_n1215), .B1(G213), .B2(new_n679), .ZN(new_n1216));
  OAI211_X1 g1016(.A(KEYINPUT125), .B(new_n1216), .C1(new_n1180), .C2(new_n1215), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT125), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1130), .A2(new_n1171), .A3(KEYINPUT57), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT122), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1167), .A2(KEYINPUT122), .A3(KEYINPUT57), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1179), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1215), .B1(new_n1223), .B2(new_n1212), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n679), .A2(G213), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(G378), .B2(new_n1213), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1218), .B1(new_n1224), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1217), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n986), .B1(new_n1200), .B2(KEYINPUT60), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1229), .B(new_n1106), .C1(KEYINPUT60), .C2(new_n1200), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(G384), .A3(new_n1198), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(G384), .B1(new_n1230), .B2(new_n1198), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(KEYINPUT62), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1210), .B1(new_n1228), .B2(new_n1236), .ZN(new_n1237));
  AOI211_X1 g1037(.A(KEYINPUT126), .B(new_n1235), .C1(new_n1217), .C2(new_n1227), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1239));
  AOI21_X1  g1039(.A(KEYINPUT62), .B1(new_n1239), .B2(new_n1234), .ZN(new_n1240));
  NOR3_X1   g1040(.A1(new_n1237), .A2(new_n1238), .A3(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n679), .A2(G213), .A3(G2897), .ZN(new_n1242));
  OR2_X1    g1042(.A1(new_n1225), .A2(KEYINPUT124), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1234), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1242), .B1(new_n1234), .B2(new_n1243), .ZN(new_n1245));
  NOR2_X1   g1045(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1246), .A2(new_n1227), .A3(new_n1217), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT61), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(KEYINPUT127), .B1(new_n1241), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1046), .B1(new_n959), .B2(new_n984), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1204), .A2(new_n1251), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(G393), .B(G396), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1252), .B(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1228), .A2(new_n1236), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(KEYINPUT126), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1240), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1228), .A2(new_n1210), .A3(new_n1236), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT127), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1250), .A2(new_n1254), .A3(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1253), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1252), .B(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1228), .A2(KEYINPUT63), .A3(new_n1234), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1246), .ZN(new_n1267));
  OAI21_X1  g1067(.A(KEYINPUT63), .B1(new_n1267), .B2(new_n1239), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1239), .A2(new_n1234), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT61), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1265), .A2(new_n1266), .A3(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1263), .A2(new_n1271), .ZN(G405));
  NOR2_X1   g1072(.A1(new_n1206), .A2(new_n1224), .ZN(new_n1273));
  XOR2_X1   g1073(.A(new_n1273), .B(new_n1234), .Z(new_n1274));
  XNOR2_X1  g1074(.A(new_n1265), .B(new_n1274), .ZN(G402));
endmodule


