//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 0 0 1 1 0 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n816, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027, new_n1028;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g002(.A1(G85gat), .A2(G92gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT7), .ZN(new_n205));
  INV_X1    g004(.A(G99gat), .ZN(new_n206));
  INV_X1    g005(.A(G106gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT8), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  OAI211_X1 g007(.A(new_n205), .B(new_n208), .C1(G85gat), .C2(G92gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(G99gat), .B(G106gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n209), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G57gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n212), .A2(G64gat), .ZN(new_n213));
  INV_X1    g012(.A(G64gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n214), .A2(G57gat), .ZN(new_n215));
  AND2_X1   g014(.A1(G71gat), .A2(G78gat), .ZN(new_n216));
  OAI22_X1  g015(.A1(new_n213), .A2(new_n215), .B1(new_n216), .B2(KEYINPUT9), .ZN(new_n217));
  XNOR2_X1  g016(.A(G71gat), .B(G78gat), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n210), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT104), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n211), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(new_n221), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n209), .A2(new_n220), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n209), .A2(new_n220), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT10), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n222), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n211), .A2(KEYINPUT10), .A3(new_n219), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n203), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n202), .B1(new_n222), .B2(new_n226), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G120gat), .B(G148gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(G176gat), .B(G204gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(KEYINPUT105), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT105), .ZN(new_n238));
  NOR4_X1   g037(.A1(new_n230), .A2(new_n238), .A3(new_n231), .A4(new_n235), .ZN(new_n239));
  OR2_X1    g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n235), .B1(new_n230), .B2(new_n231), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT18), .ZN(new_n244));
  XNOR2_X1  g043(.A(G15gat), .B(G22gat), .ZN(new_n245));
  INV_X1    g044(.A(G1gat), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(KEYINPUT16), .A3(new_n246), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(G8gat), .A3(new_n248), .ZN(new_n249));
  OR2_X1    g048(.A1(new_n249), .A2(KEYINPUT97), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(KEYINPUT97), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n247), .A2(new_n248), .ZN(new_n253));
  INV_X1    g052(.A(G8gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT98), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n253), .A2(KEYINPUT98), .A3(new_n254), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n252), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT14), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n261), .B1(G29gat), .B2(G36gat), .ZN(new_n262));
  OR3_X1    g061(.A1(new_n261), .A2(G29gat), .A3(G36gat), .ZN(new_n263));
  XOR2_X1   g062(.A(KEYINPUT95), .B(G36gat), .Z(new_n264));
  INV_X1    g063(.A(G29gat), .ZN(new_n265));
  OAI211_X1 g064(.A(new_n262), .B(new_n263), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT15), .ZN(new_n267));
  XOR2_X1   g066(.A(G43gat), .B(G50gat), .Z(new_n268));
  AOI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT96), .ZN(new_n270));
  OAI22_X1  g069(.A1(new_n266), .A2(new_n270), .B1(new_n267), .B2(new_n268), .ZN(new_n271));
  OR2_X1    g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT17), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n269), .A2(new_n271), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT99), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n260), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n272), .A2(new_n274), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n251), .A2(new_n250), .B1(new_n257), .B2(new_n258), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n273), .B1(new_n279), .B2(KEYINPUT99), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G229gat), .A2(G233gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n244), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n278), .A2(KEYINPUT100), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n279), .B1(KEYINPUT100), .B2(new_n278), .ZN(new_n287));
  OR2_X1    g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n282), .B(KEYINPUT13), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n286), .A2(new_n287), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n280), .A2(new_n278), .ZN(new_n293));
  OAI211_X1 g092(.A(KEYINPUT18), .B(new_n282), .C1(new_n293), .C2(new_n277), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n284), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G113gat), .B(G141gat), .ZN(new_n296));
  INV_X1    g095(.A(G197gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  XNOR2_X1  g097(.A(KEYINPUT11), .B(G169gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(KEYINPUT12), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n295), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n284), .A2(new_n292), .A3(new_n301), .A4(new_n294), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n243), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT77), .B(KEYINPUT6), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT71), .ZN(new_n308));
  AND2_X1   g107(.A1(KEYINPUT70), .A2(G120gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(KEYINPUT70), .A2(G120gat), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n308), .B(G113gat), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  OR2_X1    g110(.A1(G127gat), .A2(G134gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(G127gat), .A2(G134gat), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT1), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G113gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT70), .ZN(new_n316));
  INV_X1    g115(.A(G120gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(KEYINPUT70), .A2(G120gat), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n315), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n315), .A2(G120gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT71), .ZN(new_n322));
  OAI211_X1 g121(.A(new_n311), .B(new_n314), .C1(new_n320), .C2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n317), .A2(G113gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT1), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n313), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n323), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT4), .ZN(new_n332));
  AND2_X1   g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333));
  NOR2_X1   g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G141gat), .B(G148gat), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT2), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n337), .B1(G155gat), .B2(G162gat), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n335), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G148gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G141gat), .ZN(new_n341));
  INV_X1    g140(.A(G141gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G148gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G155gat), .B(G162gat), .ZN(new_n345));
  INV_X1    g144(.A(G155gat), .ZN(new_n346));
  INV_X1    g145(.A(G162gat), .ZN(new_n347));
  OAI21_X1  g146(.A(KEYINPUT2), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n344), .A2(new_n345), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n339), .A2(new_n349), .ZN(new_n350));
  NOR3_X1   g149(.A1(new_n331), .A2(new_n332), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  AOI22_X1  g151(.A1(KEYINPUT3), .A2(new_n350), .B1(new_n323), .B2(new_n330), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT3), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n349), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n332), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n350), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n339), .A2(new_n349), .A3(KEYINPUT74), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n331), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n352), .B1(new_n356), .B2(new_n360), .ZN(new_n361));
  XOR2_X1   g160(.A(KEYINPUT76), .B(KEYINPUT5), .Z(new_n362));
  NAND2_X1  g161(.A1(G225gat), .A2(G233gat), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  OR2_X1    g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT75), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n331), .A2(new_n350), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n344), .A2(new_n345), .A3(new_n348), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n345), .B1(new_n344), .B2(new_n348), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT3), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n371), .A2(new_n331), .A3(new_n355), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n368), .B1(new_n372), .B2(KEYINPUT4), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n328), .B1(new_n326), .B2(new_n325), .ZN(new_n374));
  AND2_X1   g173(.A1(G127gat), .A2(G134gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(G127gat), .A2(G134gat), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n326), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(G113gat), .B1(new_n309), .B2(new_n310), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n308), .B1(new_n315), .B2(G120gat), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n374), .B1(new_n380), .B2(new_n311), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n339), .A2(new_n349), .A3(KEYINPUT74), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT74), .B1(new_n339), .B2(new_n349), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n381), .B(KEYINPUT4), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(new_n363), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n367), .B1(new_n373), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n372), .A2(KEYINPUT4), .ZN(new_n387));
  INV_X1    g186(.A(new_n350), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n381), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n364), .B1(new_n360), .B2(KEYINPUT4), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT75), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n331), .B(new_n388), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n362), .B1(new_n394), .B2(new_n363), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n366), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G1gat), .B(G29gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n398), .B(G85gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT0), .B(G57gat), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n399), .B(new_n400), .Z(new_n401));
  AOI21_X1  g200(.A(new_n307), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT78), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n397), .ZN(new_n405));
  INV_X1    g204(.A(new_n401), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n405), .A2(KEYINPUT79), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n402), .A2(new_n403), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT79), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n409), .B1(new_n397), .B2(new_n401), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n404), .A2(new_n407), .A3(new_n408), .A4(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n395), .B1(new_n386), .B2(new_n392), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n406), .B(new_n307), .C1(new_n412), .C2(new_n366), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G211gat), .B(G218gat), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  AND2_X1   g215(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(KEYINPUT72), .A2(G211gat), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT22), .B1(new_n419), .B2(G218gat), .ZN(new_n420));
  INV_X1    g219(.A(G204gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n297), .A2(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(G197gat), .A2(G204gat), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n416), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT22), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT72), .B(G211gat), .ZN(new_n427));
  INV_X1    g226(.A(G218gat), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n424), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n430), .A3(new_n415), .ZN(new_n431));
  AND2_X1   g230(.A1(new_n425), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(G226gat), .A2(G233gat), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(G169gat), .ZN(new_n435));
  INV_X1    g234(.A(G176gat), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n436), .A3(KEYINPUT23), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT23), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n438), .B1(G169gat), .B2(G176gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(G169gat), .A2(G176gat), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n437), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT24), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(G183gat), .A3(G190gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(G183gat), .A2(G190gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT24), .ZN(new_n445));
  NOR2_X1   g244(.A1(G183gat), .A2(G190gat), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT65), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n441), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  OAI211_X1 g248(.A(KEYINPUT65), .B(new_n443), .C1(new_n445), .C2(new_n446), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(KEYINPUT25), .A3(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT25), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n452), .B1(new_n447), .B2(new_n441), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT64), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT64), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n455), .B(new_n452), .C1(new_n447), .C2(new_n441), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n451), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT68), .ZN(new_n458));
  AND4_X1   g257(.A1(KEYINPUT66), .A2(KEYINPUT67), .A3(KEYINPUT27), .A4(G183gat), .ZN(new_n459));
  AOI22_X1  g258(.A1(KEYINPUT66), .A2(KEYINPUT27), .B1(KEYINPUT67), .B2(G183gat), .ZN(new_n460));
  NOR2_X1   g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(G190gat), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT27), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n463), .A2(G183gat), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n462), .B1(new_n464), .B2(KEYINPUT66), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n458), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT28), .ZN(new_n467));
  INV_X1    g266(.A(G183gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT27), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT66), .ZN(new_n470));
  AOI21_X1  g269(.A(G190gat), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n471), .B(KEYINPUT68), .C1(new_n460), .C2(new_n459), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n466), .A2(new_n467), .A3(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT27), .B(G183gat), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n474), .A2(KEYINPUT28), .A3(new_n462), .ZN(new_n475));
  OR3_X1    g274(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(new_n477), .A3(new_n440), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n444), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT69), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n478), .A2(KEYINPUT69), .A3(new_n444), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n473), .A2(new_n475), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n434), .B1(new_n457), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(KEYINPUT73), .B(KEYINPUT29), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n473), .A2(new_n475), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n481), .A2(new_n482), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n451), .A2(new_n454), .A3(new_n456), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n432), .B(new_n484), .C1(new_n490), .C2(new_n434), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n433), .B1(new_n488), .B2(new_n489), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT29), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(new_n457), .B2(new_n483), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n492), .B1(new_n433), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n491), .B1(new_n495), .B2(new_n432), .ZN(new_n496));
  XNOR2_X1  g295(.A(G8gat), .B(G36gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(G64gat), .B(G92gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n497), .B(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n491), .B(new_n499), .C1(new_n495), .C2(new_n432), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(KEYINPUT30), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT30), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n496), .A2(new_n504), .A3(new_n500), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n414), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n382), .A2(new_n383), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n485), .B1(new_n425), .B2(new_n431), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n508), .B1(new_n509), .B2(KEYINPUT3), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT81), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OAI211_X1 g311(.A(KEYINPUT81), .B(new_n508), .C1(new_n509), .C2(KEYINPUT3), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT82), .ZN(new_n514));
  INV_X1    g313(.A(new_n485), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n355), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n425), .A2(new_n431), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n355), .A2(new_n515), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n432), .A2(KEYINPUT82), .A3(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n512), .A2(new_n513), .A3(new_n518), .A4(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(G228gat), .ZN(new_n522));
  INV_X1    g321(.A(G233gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n521), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT83), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT86), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT85), .B1(new_n432), .B2(new_n519), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT85), .ZN(new_n531));
  NOR3_X1   g330(.A1(new_n516), .A2(new_n517), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n524), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT84), .B1(new_n432), .B2(KEYINPUT29), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT29), .B1(new_n425), .B2(new_n431), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT84), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT3), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n388), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n529), .B1(new_n533), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n535), .A2(new_n536), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n354), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n535), .A2(new_n536), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n350), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n531), .B1(new_n516), .B2(new_n517), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n432), .A2(KEYINPUT85), .A3(new_n519), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n525), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n543), .A2(KEYINPUT86), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n539), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n521), .A2(KEYINPUT83), .A3(new_n525), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n528), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(G22gat), .ZN(new_n551));
  INV_X1    g350(.A(G22gat), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n528), .A2(new_n548), .A3(new_n552), .A4(new_n549), .ZN(new_n553));
  XNOR2_X1  g352(.A(G78gat), .B(G106gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(KEYINPUT31), .B(G50gat), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n551), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n557), .A2(KEYINPUT88), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT88), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n551), .A2(new_n559), .A3(new_n553), .A4(new_n556), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n551), .A2(new_n553), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n556), .B(KEYINPUT80), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT87), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT87), .ZN(new_n566));
  AOI211_X1 g365(.A(new_n566), .B(new_n563), .C1(new_n551), .C2(new_n553), .ZN(new_n567));
  OAI22_X1  g366(.A1(new_n558), .A2(new_n561), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G15gat), .B(G43gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(G71gat), .B(G99gat), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n569), .B(new_n570), .Z(new_n571));
  INV_X1    g370(.A(G227gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(new_n523), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n331), .B1(new_n457), .B2(new_n483), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n488), .A2(new_n381), .A3(new_n489), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n571), .B1(new_n577), .B2(KEYINPUT33), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n576), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(new_n573), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT34), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n580), .A2(KEYINPUT32), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT32), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT34), .B1(new_n577), .B2(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n579), .A2(new_n573), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n582), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n586), .B1(new_n582), .B2(new_n584), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n578), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n582), .A2(new_n584), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(new_n585), .ZN(new_n592));
  INV_X1    g391(.A(new_n578), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(new_n587), .A3(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n568), .A2(KEYINPUT35), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(KEYINPUT36), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n590), .A2(new_n594), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT36), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  AND3_X1   g400(.A1(new_n521), .A2(KEYINPUT83), .A3(new_n525), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT83), .B1(new_n521), .B2(new_n525), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n552), .B1(new_n604), .B2(new_n548), .ZN(new_n605));
  AND4_X1   g404(.A1(new_n552), .A2(new_n528), .A3(new_n548), .A4(new_n549), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n564), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(new_n566), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n562), .A2(KEYINPUT87), .A3(new_n564), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n557), .A2(KEYINPUT88), .ZN(new_n610));
  AOI22_X1  g409(.A1(new_n608), .A2(new_n609), .B1(new_n610), .B2(new_n560), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n601), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n507), .B1(new_n596), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n611), .B1(new_n597), .B2(new_n600), .ZN(new_n615));
  OAI21_X1  g414(.A(KEYINPUT91), .B1(new_n397), .B2(new_n401), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT91), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n617), .B(new_n406), .C1(new_n412), .C2(new_n366), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n619), .A2(new_n505), .A3(new_n503), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT89), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n351), .B1(new_n387), .B2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n621), .B1(new_n623), .B2(new_n363), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n361), .A2(KEYINPUT89), .A3(new_n364), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n406), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n627), .B1(new_n394), .B2(new_n363), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n624), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  AOI211_X1 g429(.A(KEYINPUT90), .B(KEYINPUT40), .C1(new_n628), .C2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT90), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n623), .A2(new_n621), .A3(new_n363), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT89), .B1(new_n361), .B2(new_n364), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n627), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n635), .A2(new_n401), .A3(new_n630), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT40), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n632), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n631), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n628), .A2(KEYINPUT40), .A3(new_n630), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n620), .A2(new_n639), .A3(KEYINPUT92), .A4(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT92), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n636), .A2(new_n637), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(KEYINPUT90), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n636), .A2(new_n632), .A3(new_n637), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n619), .A2(new_n505), .A3(new_n503), .A4(new_n640), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n642), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n413), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n649), .B1(new_n619), .B2(new_n402), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT37), .ZN(new_n651));
  INV_X1    g450(.A(new_n491), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n494), .A2(new_n433), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n432), .B1(new_n653), .B2(new_n484), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n651), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  OAI211_X1 g454(.A(KEYINPUT37), .B(new_n491), .C1(new_n495), .C2(new_n432), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n655), .A2(new_n499), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(KEYINPUT38), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT93), .ZN(new_n659));
  INV_X1    g458(.A(new_n501), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n653), .A2(new_n432), .A3(new_n484), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n515), .B1(new_n457), .B2(new_n483), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n492), .B1(new_n662), .B2(new_n433), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n661), .B(KEYINPUT37), .C1(new_n432), .C2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(KEYINPUT38), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n500), .B1(new_n496), .B2(new_n651), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n660), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT93), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n657), .A2(new_n669), .A3(KEYINPUT38), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n650), .A2(new_n659), .A3(new_n668), .A4(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n641), .A2(new_n648), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT94), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n598), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n590), .A2(KEYINPUT94), .A3(new_n594), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n506), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n650), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n676), .A2(new_n568), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT35), .ZN(new_n680));
  AOI22_X1  g479(.A1(new_n615), .A2(new_n672), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n306), .B1(new_n614), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n219), .A2(KEYINPUT21), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n279), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(G183gat), .ZN(new_n685));
  INV_X1    g484(.A(G231gat), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n685), .B1(new_n686), .B2(new_n523), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n684), .B(new_n468), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n688), .A2(G231gat), .A3(G233gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(G127gat), .B(G155gat), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT20), .Z(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n687), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n692), .B1(new_n687), .B2(new_n689), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n219), .A2(KEYINPUT21), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT101), .B(KEYINPUT19), .Z(new_n696));
  XOR2_X1   g495(.A(new_n696), .B(G211gat), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n695), .B(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  OR3_X1    g498(.A1(new_n693), .A2(new_n694), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n699), .B1(new_n693), .B2(new_n694), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n278), .A2(KEYINPUT17), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n704), .B(new_n275), .C1(new_n224), .C2(new_n225), .ZN(new_n705));
  XOR2_X1   g504(.A(G190gat), .B(G218gat), .Z(new_n706));
  INV_X1    g505(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT103), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n272), .A2(new_n211), .A3(new_n274), .ZN(new_n709));
  NAND3_X1  g508(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n710));
  AND3_X1   g509(.A1(new_n709), .A2(KEYINPUT102), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT102), .B1(new_n709), .B2(new_n710), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n705), .B(new_n708), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OR2_X1    g514(.A1(new_n711), .A2(new_n712), .ZN(new_n716));
  INV_X1    g515(.A(new_n714), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n716), .A2(new_n717), .A3(new_n708), .A4(new_n705), .ZN(new_n718));
  XNOR2_X1  g517(.A(G134gat), .B(G162gat), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  AND3_X1   g519(.A1(new_n715), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n720), .B1(new_n715), .B2(new_n718), .ZN(new_n722));
  OAI22_X1  g521(.A1(new_n721), .A2(new_n722), .B1(KEYINPUT103), .B2(new_n707), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n715), .A2(new_n718), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n719), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n707), .A2(KEYINPUT103), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n715), .A2(new_n718), .A3(new_n720), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n703), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n682), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(new_n414), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(new_n246), .ZN(G1324gat));
  NOR2_X1   g532(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n731), .A2(new_n506), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT42), .ZN(new_n736));
  NAND2_X1  g535(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n736), .B1(new_n735), .B2(new_n737), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n740));
  INV_X1    g539(.A(new_n731), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n677), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n740), .B1(new_n742), .B2(G8gat), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n740), .B(G8gat), .C1(new_n731), .C2(new_n506), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  OAI22_X1  g544(.A1(new_n738), .A2(new_n739), .B1(new_n743), .B2(new_n745), .ZN(G1325gat));
  INV_X1    g545(.A(G15gat), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n731), .A2(new_n747), .A3(new_n601), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n741), .A2(new_n676), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n748), .B1(new_n747), .B2(new_n749), .ZN(G1326gat));
  NOR2_X1   g549(.A1(new_n731), .A2(new_n568), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT43), .B(G22gat), .Z(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1327gat));
  NAND3_X1  g552(.A1(new_n672), .A2(new_n568), .A3(new_n601), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n674), .A2(new_n675), .ZN(new_n755));
  INV_X1    g554(.A(new_n678), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n611), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n754), .B1(new_n757), .B2(KEYINPUT35), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n729), .B1(new_n758), .B2(new_n613), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n702), .A2(new_n306), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n414), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n762), .A2(new_n265), .A3(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT45), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n759), .A2(new_n766), .ZN(new_n767));
  OAI211_X1 g566(.A(KEYINPUT44), .B(new_n729), .C1(new_n758), .C2(new_n613), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n769), .A2(new_n414), .A3(new_n761), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n765), .B1(new_n265), .B2(new_n770), .ZN(G1328gat));
  NAND3_X1  g570(.A1(new_n762), .A2(new_n264), .A3(new_n677), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n772), .B(KEYINPUT46), .Z(new_n773));
  NOR3_X1   g572(.A1(new_n769), .A2(new_n506), .A3(new_n761), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n264), .B2(new_n774), .ZN(G1329gat));
  NAND2_X1  g574(.A1(new_n614), .A2(new_n681), .ZN(new_n776));
  INV_X1    g575(.A(G43gat), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n776), .A2(new_n777), .A3(new_n729), .A4(new_n760), .ZN(new_n778));
  OAI21_X1  g577(.A(KEYINPUT107), .B1(new_n778), .B2(new_n755), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT107), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n762), .A2(new_n780), .A3(new_n777), .A4(new_n676), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(new_n601), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n767), .A2(new_n783), .A3(new_n768), .A4(new_n760), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G43gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT47), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n782), .A2(KEYINPUT47), .A3(new_n785), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(G1330gat));
  NAND4_X1  g589(.A1(new_n767), .A2(new_n611), .A3(new_n768), .A4(new_n760), .ZN(new_n791));
  AOI21_X1  g590(.A(KEYINPUT108), .B1(new_n791), .B2(G50gat), .ZN(new_n792));
  NOR4_X1   g591(.A1(new_n759), .A2(G50gat), .A3(new_n568), .A4(new_n761), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n793), .B1(new_n791), .B2(G50gat), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT48), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n792), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  AOI221_X4 g595(.A(new_n793), .B1(KEYINPUT108), .B2(KEYINPUT48), .C1(new_n791), .C2(G50gat), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n796), .A2(new_n797), .ZN(G1331gat));
  NOR3_X1   g597(.A1(new_n703), .A2(new_n729), .A3(new_n305), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n776), .A2(new_n242), .A3(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n800), .A2(new_n414), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(new_n212), .ZN(G1332gat));
  INV_X1    g601(.A(KEYINPUT49), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n776), .A2(new_n677), .A3(new_n242), .A4(new_n799), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n803), .A2(new_n214), .ZN(new_n805));
  OR3_X1    g604(.A1(new_n804), .A2(KEYINPUT109), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT109), .B1(new_n804), .B2(new_n805), .ZN(new_n807));
  AND4_X1   g606(.A1(new_n803), .A2(new_n806), .A3(new_n214), .A4(new_n807), .ZN(new_n808));
  AOI22_X1  g607(.A1(new_n806), .A2(new_n807), .B1(new_n803), .B2(new_n214), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n808), .A2(new_n809), .ZN(G1333gat));
  OAI21_X1  g609(.A(G71gat), .B1(new_n800), .B2(new_n601), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n755), .A2(G71gat), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n811), .B1(new_n800), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n813), .B(new_n814), .ZN(G1334gat));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n568), .ZN(new_n816));
  XOR2_X1   g615(.A(new_n816), .B(G78gat), .Z(G1335gat));
  INV_X1    g616(.A(KEYINPUT51), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n702), .A2(new_n305), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT110), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n776), .A2(new_n818), .A3(new_n729), .A4(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n821), .B(new_n729), .C1(new_n758), .C2(new_n613), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT51), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n822), .A2(new_n824), .A3(new_n242), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n825), .A2(new_n414), .ZN(new_n826));
  INV_X1    g625(.A(G85gat), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n821), .A2(new_n242), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n767), .A2(new_n768), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n414), .A2(new_n827), .ZN(new_n830));
  AOI22_X1  g629(.A1(new_n826), .A2(new_n827), .B1(new_n829), .B2(new_n830), .ZN(G1336gat));
  OAI21_X1  g630(.A(new_n823), .B1(KEYINPUT111), .B2(KEYINPUT51), .ZN(new_n832));
  NOR2_X1   g631(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n776), .A2(new_n729), .A3(new_n821), .A4(new_n833), .ZN(new_n834));
  AND3_X1   g633(.A1(new_n832), .A2(new_n834), .A3(new_n242), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n506), .A2(G92gat), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n767), .A2(new_n828), .A3(new_n677), .A4(new_n768), .ZN(new_n837));
  AOI22_X1  g636(.A1(new_n835), .A2(new_n836), .B1(G92gat), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n825), .A2(G92gat), .A3(new_n506), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(G92gat), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n839), .ZN(new_n842));
  OAI22_X1  g641(.A1(new_n838), .A2(new_n839), .B1(new_n840), .B2(new_n842), .ZN(G1337gat));
  NAND4_X1  g642(.A1(new_n767), .A2(new_n828), .A3(new_n783), .A4(new_n768), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n844), .A2(KEYINPUT112), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(KEYINPUT112), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n845), .A2(G99gat), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n676), .A2(new_n206), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n825), .B2(new_n848), .ZN(G1338gat));
  NOR2_X1   g648(.A1(new_n568), .A2(G106gat), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n767), .A2(new_n828), .A3(new_n611), .A4(new_n768), .ZN(new_n851));
  AOI22_X1  g650(.A1(new_n835), .A2(new_n850), .B1(G106gat), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n853));
  NAND4_X1  g652(.A1(new_n822), .A2(new_n824), .A3(new_n242), .A4(new_n850), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT113), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n853), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n851), .A2(G106gat), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n857), .B1(new_n854), .B2(KEYINPUT113), .ZN(new_n858));
  OAI22_X1  g657(.A1(new_n852), .A2(new_n853), .B1(new_n856), .B2(new_n858), .ZN(G1339gat));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n281), .A2(new_n283), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT115), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n281), .A2(new_n863), .A3(new_n283), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n290), .B1(new_n288), .B2(new_n291), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n300), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n242), .A3(new_n304), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n237), .A2(new_n239), .ZN(new_n869));
  INV_X1    g668(.A(new_n230), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n228), .A2(new_n203), .A3(new_n229), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(KEYINPUT54), .A3(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n236), .B1(new_n230), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n872), .A2(KEYINPUT55), .A3(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT114), .B1(new_n869), .B2(new_n875), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n872), .A2(new_n874), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n877), .A2(KEYINPUT55), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n872), .A2(KEYINPUT55), .A3(new_n874), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n879), .B(new_n880), .C1(new_n237), .C2(new_n239), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n876), .A2(new_n878), .A3(new_n881), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n303), .A2(new_n304), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n868), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n723), .A2(new_n728), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n867), .A2(new_n304), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n729), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n702), .B1(new_n886), .B2(new_n889), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n702), .A2(new_n885), .A3(new_n243), .A4(new_n883), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n860), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n885), .A2(new_n882), .A3(new_n887), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n305), .A2(new_n878), .A3(new_n881), .A4(new_n876), .ZN(new_n895));
  AOI22_X1  g694(.A1(new_n895), .A2(new_n868), .B1(new_n728), .B2(new_n723), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n703), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n897), .A2(KEYINPUT116), .A3(new_n891), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n611), .A2(new_n755), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n414), .A2(new_n677), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n893), .A2(new_n898), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(G113gat), .B1(new_n901), .B2(new_n883), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n611), .A2(new_n598), .ZN(new_n903));
  NAND4_X1  g702(.A1(new_n893), .A2(new_n898), .A3(new_n903), .A4(new_n900), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n305), .A2(new_n315), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n902), .B1(new_n904), .B2(new_n905), .ZN(G1340gat));
  OAI21_X1  g705(.A(G120gat), .B1(new_n901), .B2(new_n243), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n242), .B1(new_n310), .B2(new_n309), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT117), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n907), .B1(new_n904), .B2(new_n909), .ZN(G1341gat));
  INV_X1    g709(.A(G127gat), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n901), .A2(new_n911), .A3(new_n703), .ZN(new_n912));
  INV_X1    g711(.A(new_n904), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n702), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n911), .B2(new_n914), .ZN(G1342gat));
  OAI21_X1  g714(.A(G134gat), .B1(new_n901), .B2(new_n885), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT56), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n904), .A2(G134gat), .A3(new_n885), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n918), .A2(KEYINPUT118), .A3(new_n917), .ZN(new_n919));
  AOI21_X1  g718(.A(KEYINPUT118), .B1(new_n918), .B2(new_n917), .ZN(new_n920));
  OAI221_X1 g719(.A(new_n916), .B1(new_n917), .B2(new_n918), .C1(new_n919), .C2(new_n920), .ZN(G1343gat));
  INV_X1    g720(.A(KEYINPUT57), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n893), .A2(new_n898), .A3(new_n922), .A4(new_n611), .ZN(new_n923));
  INV_X1    g722(.A(new_n900), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n924), .A2(new_n783), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n867), .A2(new_n304), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n877), .A2(KEYINPUT119), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT55), .B1(new_n877), .B2(KEYINPUT119), .ZN(new_n928));
  AOI22_X1  g727(.A1(new_n927), .A2(new_n928), .B1(new_n303), .B2(new_n304), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n869), .A2(new_n875), .ZN(new_n930));
  AOI22_X1  g729(.A1(new_n242), .A2(new_n926), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n889), .B1(new_n931), .B2(new_n729), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n892), .B1(new_n932), .B2(new_n703), .ZN(new_n933));
  OAI21_X1  g732(.A(KEYINPUT57), .B1(new_n933), .B2(new_n568), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n923), .A2(new_n925), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(G141gat), .B1(new_n935), .B2(new_n883), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n893), .A2(new_n898), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n937), .A2(new_n612), .A3(new_n924), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n938), .A2(new_n342), .A3(new_n305), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(KEYINPUT58), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT58), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n936), .A2(new_n942), .A3(new_n939), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1344gat));
  NAND4_X1  g743(.A1(new_n923), .A2(new_n934), .A3(new_n242), .A4(new_n925), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n340), .A2(KEYINPUT59), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT121), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT121), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n945), .A2(new_n949), .A3(new_n946), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT59), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n893), .A2(new_n898), .A3(new_n611), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT57), .ZN(new_n954));
  OR3_X1    g753(.A1(new_n933), .A2(KEYINPUT57), .A3(new_n568), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n954), .A2(new_n955), .A3(new_n242), .A4(new_n925), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n952), .B1(new_n956), .B2(G148gat), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n938), .A2(new_n340), .A3(new_n242), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n958), .A2(KEYINPUT120), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n958), .A2(KEYINPUT120), .ZN(new_n960));
  OAI22_X1  g759(.A1(new_n951), .A2(new_n957), .B1(new_n959), .B2(new_n960), .ZN(G1345gat));
  NOR3_X1   g760(.A1(new_n935), .A2(new_n346), .A3(new_n703), .ZN(new_n962));
  AOI21_X1  g761(.A(G155gat), .B1(new_n938), .B2(new_n702), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n962), .A2(new_n963), .ZN(G1346gat));
  NOR3_X1   g763(.A1(new_n935), .A2(new_n347), .A3(new_n885), .ZN(new_n965));
  AOI21_X1  g764(.A(G162gat), .B1(new_n938), .B2(new_n729), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n965), .A2(new_n966), .ZN(G1347gat));
  NOR3_X1   g766(.A1(new_n763), .A2(KEYINPUT123), .A3(new_n506), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n969), .B1(new_n414), .B2(new_n677), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n893), .A2(new_n898), .A3(new_n899), .A4(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(G169gat), .B1(new_n972), .B2(new_n883), .ZN(new_n973));
  NOR2_X1   g772(.A1(new_n937), .A2(new_n763), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n611), .A2(new_n598), .A3(new_n506), .ZN(new_n975));
  OR2_X1    g774(.A1(new_n975), .A2(KEYINPUT122), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(KEYINPUT122), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n974), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n305), .A2(new_n435), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n973), .B1(new_n978), .B2(new_n979), .ZN(G1348gat));
  OAI21_X1  g779(.A(G176gat), .B1(new_n972), .B2(new_n243), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n242), .A2(new_n436), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n981), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n983), .B(KEYINPUT124), .ZN(G1349gat));
  AND2_X1   g783(.A1(new_n702), .A2(new_n474), .ZN(new_n985));
  NAND4_X1  g784(.A1(new_n974), .A2(new_n976), .A3(new_n977), .A4(new_n985), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT125), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n987), .A2(KEYINPUT60), .ZN(new_n988));
  OAI21_X1  g787(.A(G183gat), .B1(new_n972), .B2(new_n703), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n986), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  OR2_X1    g789(.A1(new_n987), .A2(KEYINPUT60), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n990), .B(new_n991), .ZN(G1350gat));
  OR3_X1    g791(.A1(new_n978), .A2(G190gat), .A3(new_n885), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT61), .ZN(new_n994));
  OR2_X1    g793(.A1(new_n972), .A2(new_n885), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n994), .B1(new_n995), .B2(G190gat), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n995), .A2(new_n994), .A3(G190gat), .ZN(new_n997));
  INV_X1    g796(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n993), .B1(new_n996), .B2(new_n998), .ZN(G1351gat));
  INV_X1    g798(.A(KEYINPUT127), .ZN(new_n1000));
  NOR3_X1   g799(.A1(new_n968), .A2(new_n783), .A3(new_n970), .ZN(new_n1001));
  XNOR2_X1  g800(.A(new_n1001), .B(KEYINPUT126), .ZN(new_n1002));
  NAND4_X1  g801(.A1(new_n954), .A2(new_n955), .A3(new_n305), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(G197gat), .ZN(new_n1004));
  INV_X1    g803(.A(new_n612), .ZN(new_n1005));
  NAND4_X1  g804(.A1(new_n893), .A2(new_n898), .A3(new_n414), .A4(new_n1005), .ZN(new_n1006));
  NOR2_X1   g805(.A1(new_n883), .A2(G197gat), .ZN(new_n1007));
  INV_X1    g806(.A(new_n1007), .ZN(new_n1008));
  NOR3_X1   g807(.A1(new_n1006), .A2(new_n506), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g808(.A(new_n1009), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n1000), .B1(new_n1004), .B2(new_n1010), .ZN(new_n1011));
  AOI211_X1 g810(.A(KEYINPUT127), .B(new_n1009), .C1(new_n1003), .C2(G197gat), .ZN(new_n1012));
  NOR2_X1   g811(.A1(new_n1011), .A2(new_n1012), .ZN(G1352gat));
  NOR2_X1   g812(.A1(new_n1006), .A2(new_n506), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n1014), .A2(new_n421), .A3(new_n242), .ZN(new_n1015));
  OR2_X1    g814(.A1(new_n1015), .A2(KEYINPUT62), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1015), .A2(KEYINPUT62), .ZN(new_n1017));
  AND2_X1   g816(.A1(new_n954), .A2(new_n955), .ZN(new_n1018));
  AND3_X1   g817(.A1(new_n1018), .A2(new_n242), .A3(new_n1002), .ZN(new_n1019));
  OAI211_X1 g818(.A(new_n1016), .B(new_n1017), .C1(new_n1019), .C2(new_n421), .ZN(G1353gat));
  NAND3_X1  g819(.A1(new_n1014), .A2(new_n702), .A3(new_n427), .ZN(new_n1021));
  NAND4_X1  g820(.A1(new_n954), .A2(new_n955), .A3(new_n702), .A4(new_n1001), .ZN(new_n1022));
  AND3_X1   g821(.A1(new_n1022), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1023));
  AOI21_X1  g822(.A(KEYINPUT63), .B1(new_n1022), .B2(G211gat), .ZN(new_n1024));
  OAI21_X1  g823(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(G1354gat));
  AOI21_X1  g824(.A(G218gat), .B1(new_n1014), .B2(new_n729), .ZN(new_n1026));
  AND2_X1   g825(.A1(new_n1018), .A2(new_n1002), .ZN(new_n1027));
  NOR2_X1   g826(.A1(new_n885), .A2(new_n428), .ZN(new_n1028));
  AOI21_X1  g827(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(G1355gat));
endmodule


