//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:21 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n560, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n583, new_n584, new_n585, new_n586, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n633, new_n634, new_n635, new_n636, new_n639,
    new_n640, new_n642, new_n643, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT66), .Z(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n460), .B1(new_n453), .B2(G2106), .ZN(new_n461));
  XNOR2_X1  g036(.A(new_n461), .B(KEYINPUT67), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT68), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n466), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n471), .A2(G137), .B1(G101), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n470), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n469), .A2(KEYINPUT68), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n475), .A2(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n471), .A2(G136), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n466), .A2(new_n472), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  OR2_X1    g060(.A1(new_n464), .A2(new_n465), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(new_n472), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n471), .A2(KEYINPUT4), .A3(G138), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G2105), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n479), .B2(G126), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n489), .A2(new_n490), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT69), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n489), .A2(new_n497), .A3(new_n494), .A4(new_n490), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n501), .B1(new_n502), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(KEYINPUT70), .A3(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n506), .B1(new_n504), .B2(KEYINPUT5), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n502), .A2(KEYINPUT71), .A3(G543), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n503), .A2(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AND2_X1   g087(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n504), .B1(new_n510), .B2(new_n511), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n513), .A2(G88), .B1(G50), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n503), .A2(new_n505), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n507), .A2(new_n508), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(G62), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G651), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n516), .A2(new_n524), .ZN(G166));
  NAND4_X1  g100(.A1(new_n518), .A2(new_n519), .A3(G89), .A4(new_n512), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT72), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n509), .A2(new_n531), .B1(G51), .B2(new_n514), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n526), .A2(new_n529), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT72), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(G286));
  INV_X1    g111(.A(G286), .ZN(G168));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n520), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n518), .A2(new_n519), .A3(G90), .A4(new_n512), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT73), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n514), .A2(G52), .ZN(new_n544));
  AND3_X1   g119(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n543), .B1(new_n542), .B2(new_n544), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n541), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(G171));
  AOI22_X1  g123(.A1(new_n513), .A2(G81), .B1(G43), .B2(new_n514), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n551));
  OAI21_X1  g126(.A(G651), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n520), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(KEYINPUT74), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n549), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT75), .Z(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  AND2_X1   g139(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n565));
  NOR2_X1   g140(.A1(KEYINPUT76), .A2(KEYINPUT9), .ZN(new_n566));
  OAI211_X1 g141(.A(new_n514), .B(G53), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n514), .A2(G53), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n567), .B1(new_n569), .B2(new_n566), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n513), .A2(G91), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n518), .A2(new_n519), .A3(G65), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT77), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n572), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(KEYINPUT78), .B1(new_n577), .B2(G651), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n579));
  INV_X1    g154(.A(G651), .ZN(new_n580));
  AOI211_X1 g155(.A(new_n579), .B(new_n580), .C1(new_n572), .C2(new_n576), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n570), .B(new_n571), .C1(new_n578), .C2(new_n581), .ZN(G299));
  NAND2_X1  g157(.A1(new_n547), .A2(KEYINPUT79), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n584));
  OAI211_X1 g159(.A(new_n541), .B(new_n584), .C1(new_n545), .C2(new_n546), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G301));
  INV_X1    g162(.A(G166), .ZN(G303));
  AOI22_X1  g163(.A1(new_n513), .A2(G87), .B1(G49), .B2(new_n514), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(G288));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n520), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G651), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n514), .A2(G48), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT80), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n514), .A2(KEYINPUT80), .A3(G48), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G86), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n509), .A2(new_n512), .ZN(new_n602));
  OAI211_X1 g177(.A(new_n595), .B(new_n600), .C1(new_n601), .C2(new_n602), .ZN(G305));
  NAND2_X1  g178(.A1(G72), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G60), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n520), .B2(new_n605), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n606), .A2(G651), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n514), .A2(G47), .ZN(new_n608));
  XNOR2_X1  g183(.A(KEYINPUT81), .B(G85), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n602), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(KEYINPUT82), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n610), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT82), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n606), .A2(G651), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n611), .A2(new_n615), .ZN(G290));
  NAND4_X1  g191(.A1(new_n518), .A2(new_n519), .A3(G92), .A4(new_n512), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(KEYINPUT83), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT83), .ZN(new_n619));
  NAND4_X1  g194(.A1(new_n509), .A2(new_n619), .A3(G92), .A4(new_n512), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT10), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g198(.A1(new_n618), .A2(new_n620), .A3(KEYINPUT10), .ZN(new_n624));
  NAND2_X1  g199(.A1(G79), .A2(G543), .ZN(new_n625));
  INV_X1    g200(.A(G66), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n520), .B2(new_n626), .ZN(new_n627));
  AOI22_X1  g202(.A1(new_n627), .A2(G651), .B1(G54), .B2(new_n514), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n623), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(G868), .B2(new_n586), .ZN(G321));
  XOR2_X1   g206(.A(G321), .B(KEYINPUT84), .Z(G284));
  INV_X1    g207(.A(G868), .ZN(new_n633));
  OR3_X1    g208(.A1(G168), .A2(KEYINPUT85), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(KEYINPUT85), .B1(G168), .B2(new_n633), .ZN(new_n635));
  INV_X1    g210(.A(G299), .ZN(new_n636));
  OAI211_X1 g211(.A(new_n634), .B(new_n635), .C1(G868), .C2(new_n636), .ZN(G297));
  OAI211_X1 g212(.A(new_n634), .B(new_n635), .C1(G868), .C2(new_n636), .ZN(G280));
  INV_X1    g213(.A(new_n629), .ZN(new_n639));
  INV_X1    g214(.A(G559), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n639), .B1(new_n640), .B2(G860), .ZN(G148));
  NAND2_X1  g216(.A1(new_n639), .A2(new_n640), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(G868), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g219(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g220(.A1(new_n486), .A2(new_n473), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT12), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT13), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2100), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n471), .A2(G135), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n479), .A2(G123), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n472), .A2(G111), .ZN(new_n652));
  OAI21_X1  g227(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n653));
  OAI211_X1 g228(.A(new_n650), .B(new_n651), .C1(new_n652), .C2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(KEYINPUT86), .B(G2096), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n649), .A2(new_n656), .ZN(G156));
  INV_X1    g232(.A(KEYINPUT14), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2427), .B(G2438), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2430), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT15), .B(G2435), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n662), .B1(new_n661), .B2(new_n660), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2451), .B(G2454), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT16), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1341), .B(G1348), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n663), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2443), .B(G2446), .ZN(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(G14), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n672), .B(KEYINPUT87), .Z(G401));
  INV_X1    g248(.A(KEYINPUT18), .ZN(new_n674));
  XOR2_X1   g249(.A(G2084), .B(G2090), .Z(new_n675));
  XNOR2_X1  g250(.A(G2067), .B(G2678), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(KEYINPUT17), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n675), .A2(new_n676), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n674), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n680), .B(G2100), .Z(new_n681));
  XOR2_X1   g256(.A(G2072), .B(G2078), .Z(new_n682));
  AOI21_X1  g257(.A(new_n682), .B1(new_n677), .B2(KEYINPUT18), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(G2096), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n681), .B(new_n684), .ZN(G227));
  XOR2_X1   g260(.A(G1971), .B(G1976), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT19), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1956), .B(G2474), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1961), .B(G1966), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NOR3_X1   g266(.A1(new_n687), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n687), .A2(new_n690), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT20), .Z(new_n694));
  AOI211_X1 g269(.A(new_n692), .B(new_n694), .C1(new_n687), .C2(new_n691), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1981), .B(G1986), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(G229));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G22), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G166), .B2(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(G1971), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT89), .Z(new_n707));
  NOR2_X1   g282(.A1(G16), .A2(G23), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT88), .Z(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G288), .B2(new_n702), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT33), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G1976), .ZN(new_n712));
  NOR2_X1   g287(.A1(G6), .A2(G16), .ZN(new_n713));
  INV_X1    g288(.A(G305), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n713), .B1(new_n714), .B2(G16), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT32), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G1981), .ZN(new_n717));
  NOR3_X1   g292(.A1(new_n707), .A2(new_n712), .A3(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT34), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n471), .A2(G131), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n479), .A2(G119), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n472), .A2(G107), .ZN(new_n724));
  OAI21_X1  g299(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n722), .B(new_n723), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  MUX2_X1   g301(.A(G25), .B(new_n726), .S(G29), .Z(new_n727));
  XOR2_X1   g302(.A(KEYINPUT35), .B(G1991), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n702), .A2(G24), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G290), .B2(G16), .ZN(new_n731));
  INV_X1    g306(.A(G1986), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n729), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n732), .B2(new_n731), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n720), .A2(new_n721), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g310(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT91), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n735), .A2(new_n737), .ZN(new_n739));
  INV_X1    g314(.A(G29), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G32), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n471), .A2(G141), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT96), .Z(new_n743));
  AND2_X1   g318(.A1(new_n473), .A2(G105), .ZN(new_n744));
  NAND3_X1  g319(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT26), .ZN(new_n746));
  AOI211_X1 g321(.A(new_n744), .B(new_n746), .C1(G129), .C2(new_n479), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n741), .B1(new_n749), .B2(new_n740), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT27), .B(G1996), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n740), .A2(G26), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT28), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n471), .A2(G140), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n479), .A2(G128), .ZN(new_n756));
  OR2_X1    g331(.A1(G104), .A2(G2105), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n757), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n754), .B1(new_n760), .B2(new_n740), .ZN(new_n761));
  INV_X1    g336(.A(G2067), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(G162), .A2(new_n740), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n740), .B2(G35), .ZN(new_n765));
  XOR2_X1   g340(.A(KEYINPUT29), .B(G2090), .Z(new_n766));
  AND2_X1   g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT30), .B(G28), .ZN(new_n769));
  OR2_X1    g344(.A1(KEYINPUT31), .A2(G11), .ZN(new_n770));
  NAND2_X1  g345(.A1(KEYINPUT31), .A2(G11), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n769), .A2(new_n740), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(new_n654), .B2(new_n740), .ZN(new_n773));
  NOR3_X1   g348(.A1(new_n767), .A2(new_n768), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n740), .B1(KEYINPUT24), .B2(G34), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(KEYINPUT24), .B2(G34), .ZN(new_n776));
  INV_X1    g351(.A(G160), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(G29), .ZN(new_n778));
  INV_X1    g353(.A(G2084), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n752), .A2(new_n763), .A3(new_n774), .A4(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G27), .A2(G29), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G164), .B2(G29), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G2078), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n781), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(G115), .A2(G2104), .ZN(new_n786));
  INV_X1    g361(.A(G127), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n466), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n472), .B1(new_n788), .B2(KEYINPUT93), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(KEYINPUT93), .B2(new_n788), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT92), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT25), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n471), .A2(G139), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n790), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  MUX2_X1   g370(.A(G33), .B(new_n795), .S(G29), .Z(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT94), .Z(new_n797));
  NAND2_X1  g372(.A1(new_n797), .A2(G2072), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n558), .A2(G16), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G16), .B2(G19), .ZN(new_n800));
  INV_X1    g375(.A(G1341), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(G168), .A2(new_n702), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(new_n702), .B2(G21), .ZN(new_n804));
  INV_X1    g379(.A(G1966), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n702), .A2(G5), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G171), .B2(new_n702), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(G1961), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n798), .A2(new_n802), .A3(new_n806), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n702), .A2(G20), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT23), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n636), .B2(new_n702), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(G1956), .ZN(new_n814));
  OAI22_X1  g389(.A1(new_n797), .A2(G2072), .B1(new_n800), .B2(new_n801), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n808), .A2(G1961), .ZN(new_n816));
  NOR4_X1   g391(.A1(new_n810), .A2(new_n814), .A3(new_n815), .A4(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n778), .A2(new_n779), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT95), .Z(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n805), .B2(new_n804), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n702), .A2(G4), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n639), .B2(new_n702), .ZN(new_n822));
  INV_X1    g397(.A(G1348), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  AND4_X1   g399(.A1(new_n785), .A2(new_n817), .A3(new_n820), .A4(new_n824), .ZN(new_n825));
  AND3_X1   g400(.A1(new_n738), .A2(new_n739), .A3(new_n825), .ZN(G311));
  NAND3_X1  g401(.A1(new_n738), .A2(new_n739), .A3(new_n825), .ZN(G150));
  INV_X1    g402(.A(G860), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n518), .A2(new_n519), .A3(G67), .ZN(new_n829));
  NAND2_X1  g404(.A1(G80), .A2(G543), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G651), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n518), .A2(new_n519), .A3(G93), .A4(new_n512), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n514), .A2(G55), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n828), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT37), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n639), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT98), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT38), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT97), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n832), .A2(new_n835), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n580), .B1(new_n829), .B2(new_n830), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n833), .A2(new_n834), .ZN(new_n844));
  OAI21_X1  g419(.A(KEYINPUT97), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(new_n557), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n550), .A2(new_n551), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n555), .A2(KEYINPUT74), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n848), .A2(new_n849), .A3(G651), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n850), .A2(new_n549), .A3(new_n845), .A4(new_n842), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n840), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n855), .A2(KEYINPUT39), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n828), .B1(new_n855), .B2(KEYINPUT39), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n837), .B1(new_n856), .B2(new_n857), .ZN(G145));
  INV_X1    g433(.A(G37), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n654), .B(KEYINPUT99), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(G162), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n777), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n726), .B(KEYINPUT101), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n647), .ZN(new_n864));
  AOI22_X1  g439(.A1(G130), .A2(new_n479), .B1(new_n471), .B2(G142), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n866), .A2(new_n472), .A3(G118), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n866), .B1(new_n472), .B2(G118), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n868), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n865), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n864), .B(new_n870), .Z(new_n871));
  XNOR2_X1  g446(.A(new_n495), .B(new_n759), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n795), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n748), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n871), .A2(new_n874), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(KEYINPUT102), .ZN(new_n878));
  INV_X1    g453(.A(new_n876), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n879), .A3(new_n862), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n875), .A2(KEYINPUT102), .ZN(new_n881));
  OAI221_X1 g456(.A(new_n859), .B1(new_n862), .B2(new_n877), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT40), .ZN(G395));
  OAI21_X1  g458(.A(new_n633), .B1(new_n843), .B2(new_n844), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n575), .B1(new_n509), .B2(G65), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n579), .B1(new_n885), .B2(new_n580), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n577), .A2(KEYINPUT78), .A3(G651), .ZN(new_n887));
  AOI22_X1  g462(.A1(new_n886), .A2(new_n887), .B1(G91), .B2(new_n513), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n629), .A2(new_n570), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(KEYINPUT10), .B1(new_n618), .B2(new_n620), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n514), .A2(G54), .ZN(new_n891));
  AOI22_X1  g466(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n891), .B1(new_n892), .B2(new_n580), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(G299), .A2(new_n894), .A3(new_n624), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n889), .A2(new_n895), .A3(KEYINPUT103), .ZN(new_n896));
  AOI21_X1  g471(.A(KEYINPUT103), .B1(new_n889), .B2(new_n895), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n889), .A2(new_n895), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT41), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n889), .A2(new_n895), .A3(KEYINPUT41), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n852), .B(new_n642), .ZN(new_n904));
  MUX2_X1   g479(.A(new_n898), .B(new_n903), .S(new_n904), .Z(new_n905));
  OAI211_X1 g480(.A(new_n590), .B(new_n589), .C1(new_n516), .C2(new_n524), .ZN(new_n906));
  NAND3_X1  g481(.A1(G288), .A2(new_n523), .A3(new_n515), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n611), .A2(new_n615), .A3(G305), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(G305), .B1(new_n611), .B2(new_n615), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(G290), .A2(new_n714), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n913), .A2(new_n907), .A3(new_n906), .A4(new_n909), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n915), .B(KEYINPUT42), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n905), .B(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n884), .B1(new_n917), .B2(new_n633), .ZN(G295));
  OAI21_X1  g493(.A(new_n884), .B1(new_n917), .B2(new_n633), .ZN(G331));
  AND3_X1   g494(.A1(new_n912), .A2(new_n914), .A3(KEYINPUT106), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT106), .B1(new_n912), .B2(new_n914), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(G286), .B1(new_n583), .B2(new_n585), .ZN(new_n923));
  INV_X1    g498(.A(new_n546), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AOI22_X1  g501(.A1(new_n926), .A2(new_n541), .B1(new_n533), .B2(new_n535), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n853), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n586), .A2(G168), .ZN(new_n929));
  INV_X1    g504(.A(new_n927), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(new_n852), .A3(new_n930), .ZN(new_n931));
  AOI22_X1  g506(.A1(new_n928), .A2(new_n931), .B1(new_n901), .B2(new_n902), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT105), .ZN(new_n933));
  AND4_X1   g508(.A1(new_n933), .A2(new_n929), .A3(new_n852), .A4(new_n930), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n927), .B1(new_n586), .B2(G168), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n933), .B1(new_n935), .B2(new_n852), .ZN(new_n936));
  OAI211_X1 g511(.A(new_n898), .B(new_n928), .C1(new_n934), .C2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n932), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n931), .A2(KEYINPUT105), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n935), .A2(new_n933), .A3(new_n852), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n942), .A2(KEYINPUT107), .A3(new_n898), .A4(new_n928), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n922), .B1(new_n939), .B2(new_n943), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n928), .A2(new_n899), .A3(new_n931), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n935), .A2(new_n852), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(new_n940), .B2(new_n941), .ZN(new_n947));
  INV_X1    g522(.A(new_n903), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n915), .B(new_n945), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n859), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT43), .B1(new_n944), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT108), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI211_X1 g528(.A(KEYINPUT108), .B(KEYINPUT43), .C1(new_n944), .C2(new_n950), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n928), .B1(new_n934), .B2(new_n936), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n903), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n922), .B1(new_n957), .B2(new_n945), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n950), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT43), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n955), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n953), .A2(new_n954), .A3(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n963));
  INV_X1    g538(.A(new_n950), .ZN(new_n964));
  INV_X1    g539(.A(new_n958), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n960), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n944), .A2(new_n950), .A3(KEYINPUT43), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n962), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n962), .A2(KEYINPUT109), .A3(new_n968), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(G397));
  INV_X1    g548(.A(G1384), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n495), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n476), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n977), .A2(G40), .A3(new_n474), .A4(new_n470), .ZN(new_n978));
  XNOR2_X1  g553(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n976), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n759), .B(G2067), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n983), .B1(new_n748), .B2(G1996), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G1996), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n981), .A2(new_n986), .A3(new_n749), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n988));
  OR2_X1    g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n987), .A2(new_n988), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n985), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n726), .B(new_n728), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n991), .B1(new_n982), .B2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n611), .A2(new_n615), .A3(new_n732), .ZN(new_n994));
  NAND2_X1  g569(.A1(G290), .A2(G1986), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n982), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(G8), .ZN(new_n998));
  NOR2_X1   g573(.A1(G166), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n999), .B(KEYINPUT55), .ZN(new_n1000));
  AOI21_X1  g575(.A(G1384), .B1(new_n496), .B2(new_n498), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1001), .A2(new_n980), .ZN(new_n1002));
  INV_X1    g577(.A(G40), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n475), .A2(new_n1003), .A3(new_n476), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT45), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1004), .B1(new_n1005), .B2(new_n975), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1007), .A2(G1971), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n978), .B1(new_n976), .B2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(new_n1009), .B2(new_n1001), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(G2090), .ZN(new_n1012));
  OAI211_X1 g587(.A(G8), .B(new_n1000), .C1(new_n1008), .C2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1981), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n714), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(G305), .A2(G1981), .ZN(new_n1016));
  OAI21_X1  g591(.A(KEYINPUT112), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1017), .A2(KEYINPUT49), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1004), .A2(new_n976), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(G8), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1021), .B1(new_n1017), .B2(KEYINPUT49), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n978), .A2(new_n975), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1024), .A2(new_n998), .ZN(new_n1025));
  INV_X1    g600(.A(G1976), .ZN(new_n1026));
  AOI21_X1  g601(.A(KEYINPUT52), .B1(G288), .B2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1025), .B(new_n1027), .C1(new_n1026), .C2(G288), .ZN(new_n1028));
  NOR2_X1   g603(.A1(G288), .A2(new_n1026), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT52), .B1(new_n1021), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1013), .A2(new_n1023), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT53), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n975), .A2(new_n1005), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(new_n978), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(new_n1001), .B2(new_n980), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1034), .B1(new_n1037), .B2(G2078), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1001), .A2(new_n980), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1004), .B1(new_n976), .B2(KEYINPUT45), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1034), .A2(G2078), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT123), .B(G1961), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1011), .A2(new_n1044), .ZN(new_n1045));
  AND3_X1   g620(.A1(new_n1038), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1046), .A2(G301), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1000), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1004), .B1(new_n976), .B2(new_n1009), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1049), .B1(new_n1009), .B2(new_n1001), .ZN(new_n1050));
  INV_X1    g625(.A(G2090), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1050), .A2(new_n1051), .B1(new_n1037), .B2(new_n705), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1048), .B1(new_n1052), .B2(new_n998), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1048), .B(KEYINPUT114), .C1(new_n1052), .C2(new_n998), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1033), .A2(new_n1047), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT62), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n805), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1010), .B(new_n779), .C1(new_n1009), .C2(new_n1001), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n998), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G286), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(G168), .A3(new_n1060), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n998), .A2(KEYINPUT122), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1063), .A2(KEYINPUT51), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT51), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1058), .B(new_n1062), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT125), .B1(new_n1057), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1031), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1070));
  AND4_X1   g645(.A1(new_n1055), .A2(new_n1056), .A3(new_n1013), .A4(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT125), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1071), .A2(new_n1072), .A3(new_n1047), .A4(new_n1067), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1062), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT62), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1069), .A2(new_n1073), .A3(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(G288), .A2(G1976), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1016), .B1(new_n1023), .B2(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1021), .B(KEYINPUT113), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1070), .ZN(new_n1080));
  OAI22_X1  g655(.A1(new_n1078), .A2(new_n1079), .B1(new_n1080), .B2(new_n1013), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT115), .B(KEYINPUT63), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1033), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1061), .A2(G168), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(G8), .B1(new_n1008), .B2(new_n1012), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n1048), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1084), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1033), .A2(new_n1087), .A3(KEYINPUT63), .A4(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1081), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1076), .A2(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n976), .A2(new_n980), .ZN(new_n1092));
  INV_X1    g667(.A(new_n474), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1093), .A2(KEYINPUT124), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(KEYINPUT124), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1095), .A2(G40), .A3(new_n469), .A4(new_n1042), .ZN(new_n1096));
  NOR4_X1   g671(.A1(new_n1092), .A2(new_n1035), .A3(new_n1094), .A4(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1097), .B1(new_n1011), .B2(new_n1044), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1098), .A2(G301), .A3(new_n1038), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1046), .B2(G301), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1098), .A2(new_n1038), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1101), .B1(new_n1102), .B2(G171), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1046), .A2(G301), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1100), .A2(new_n1101), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1105), .A2(new_n1071), .A3(new_n1074), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1011), .A2(new_n823), .B1(new_n762), .B2(new_n1024), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n639), .B1(new_n1107), .B2(KEYINPUT60), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT121), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1107), .A2(KEYINPUT60), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1111), .B(new_n639), .C1(new_n1107), .C2(KEYINPUT60), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1109), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1036), .B(new_n986), .C1(new_n1001), .C2(new_n980), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT58), .B(G1341), .Z(new_n1115));
  NAND2_X1  g690(.A1(new_n1020), .A2(new_n1115), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1114), .A2(KEYINPUT120), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT120), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n558), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(KEYINPUT59), .B(new_n558), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1113), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1110), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(KEYINPUT56), .B(G2072), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1007), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(G1956), .B2(new_n1050), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n636), .A2(KEYINPUT57), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n570), .A2(KEYINPUT117), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n570), .A2(KEYINPUT117), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n888), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT118), .ZN(new_n1134));
  XOR2_X1   g709(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n1135));
  AND3_X1   g710(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1134), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1130), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g715(.A(KEYINPUT119), .B(new_n1130), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1129), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1140), .A2(new_n1129), .A3(new_n1141), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1143), .A2(KEYINPUT61), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1144), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1146), .B1(new_n1147), .B2(new_n1142), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1123), .A2(new_n1126), .A3(new_n1145), .A4(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1144), .B1(new_n629), .B2(new_n1107), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n1143), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1106), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n997), .B1(new_n1091), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n981), .A2(new_n986), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT46), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n981), .B1(new_n748), .B2(new_n983), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT47), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n982), .A2(new_n994), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT127), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT48), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1158), .B1(new_n1161), .B2(new_n993), .ZN(new_n1162));
  INV_X1    g737(.A(new_n728), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n726), .A2(new_n1163), .ZN(new_n1164));
  AOI22_X1  g739(.A1(new_n991), .A2(new_n1164), .B1(new_n762), .B2(new_n760), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT126), .ZN(new_n1166));
  OR2_X1    g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n982), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1162), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1153), .A2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g745(.A(G227), .ZN(new_n1172));
  NAND3_X1  g746(.A1(G319), .A2(new_n672), .A3(new_n1172), .ZN(new_n1173));
  NOR2_X1   g747(.A1(G229), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g748(.A1(new_n1174), .A2(new_n882), .ZN(new_n1175));
  NOR2_X1   g749(.A1(new_n966), .A2(new_n967), .ZN(new_n1176));
  NOR2_X1   g750(.A1(new_n1175), .A2(new_n1176), .ZN(G308));
  INV_X1    g751(.A(G308), .ZN(G225));
endmodule


