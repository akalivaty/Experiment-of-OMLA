

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591;

  XOR2_X1 U323 ( .A(KEYINPUT71), .B(KEYINPUT13), .Z(n291) );
  XNOR2_X1 U324 ( .A(KEYINPUT47), .B(KEYINPUT113), .ZN(n382) );
  XNOR2_X1 U325 ( .A(n383), .B(n382), .ZN(n390) );
  XOR2_X1 U326 ( .A(n417), .B(n342), .Z(n586) );
  XOR2_X1 U327 ( .A(KEYINPUT41), .B(n586), .Z(n563) );
  XOR2_X1 U328 ( .A(n360), .B(n365), .Z(n582) );
  XNOR2_X1 U329 ( .A(n450), .B(KEYINPUT122), .ZN(n451) );
  XNOR2_X1 U330 ( .A(n452), .B(n451), .ZN(G1350GAT) );
  XOR2_X1 U331 ( .A(G183GAT), .B(KEYINPUT77), .Z(n309) );
  XOR2_X1 U332 ( .A(n309), .B(G155GAT), .Z(n293) );
  XOR2_X1 U333 ( .A(G1GAT), .B(KEYINPUT70), .Z(n345) );
  XNOR2_X1 U334 ( .A(n345), .B(G78GAT), .ZN(n292) );
  XNOR2_X1 U335 ( .A(n293), .B(n292), .ZN(n298) );
  XOR2_X1 U336 ( .A(G15GAT), .B(G127GAT), .Z(n432) );
  XNOR2_X1 U337 ( .A(G71GAT), .B(G57GAT), .ZN(n294) );
  XNOR2_X1 U338 ( .A(n291), .B(n294), .ZN(n332) );
  XOR2_X1 U339 ( .A(n432), .B(n332), .Z(n296) );
  NAND2_X1 U340 ( .A1(G231GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U341 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U342 ( .A(n298), .B(n297), .Z(n300) );
  XNOR2_X1 U343 ( .A(G22GAT), .B(G211GAT), .ZN(n299) );
  XNOR2_X1 U344 ( .A(n300), .B(n299), .ZN(n308) );
  XOR2_X1 U345 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n302) );
  XNOR2_X1 U346 ( .A(G8GAT), .B(G64GAT), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U348 ( .A(KEYINPUT78), .B(KEYINPUT15), .Z(n304) );
  XNOR2_X1 U349 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U351 ( .A(n306), .B(n305), .Z(n307) );
  XOR2_X1 U352 ( .A(n308), .B(n307), .Z(n590) );
  NAND2_X1 U353 ( .A1(G226GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U354 ( .A(n310), .B(n309), .ZN(n323) );
  XNOR2_X1 U355 ( .A(G176GAT), .B(G92GAT), .ZN(n311) );
  XNOR2_X1 U356 ( .A(n311), .B(G64GAT), .ZN(n331) );
  XOR2_X1 U357 ( .A(KEYINPUT76), .B(G218GAT), .Z(n313) );
  XNOR2_X1 U358 ( .A(G36GAT), .B(G190GAT), .ZN(n312) );
  XNOR2_X1 U359 ( .A(n313), .B(n312), .ZN(n376) );
  XOR2_X1 U360 ( .A(n331), .B(n376), .Z(n318) );
  XNOR2_X1 U361 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n314) );
  XNOR2_X1 U362 ( .A(n314), .B(KEYINPUT18), .ZN(n433) );
  XOR2_X1 U363 ( .A(G211GAT), .B(KEYINPUT21), .Z(n316) );
  XNOR2_X1 U364 ( .A(G197GAT), .B(KEYINPUT85), .ZN(n315) );
  XNOR2_X1 U365 ( .A(n316), .B(n315), .ZN(n412) );
  XNOR2_X1 U366 ( .A(n433), .B(n412), .ZN(n317) );
  XNOR2_X1 U367 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U368 ( .A(n319), .B(KEYINPUT91), .Z(n321) );
  XOR2_X1 U369 ( .A(G169GAT), .B(G8GAT), .Z(n346) );
  XNOR2_X1 U370 ( .A(n346), .B(G204GAT), .ZN(n320) );
  XNOR2_X1 U371 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U372 ( .A(n323), .B(n322), .Z(n506) );
  INV_X1 U373 ( .A(n506), .ZN(n529) );
  XNOR2_X1 U374 ( .A(G148GAT), .B(KEYINPUT73), .ZN(n324) );
  XNOR2_X1 U375 ( .A(n324), .B(KEYINPUT74), .ZN(n325) );
  XOR2_X1 U376 ( .A(n325), .B(G204GAT), .Z(n327) );
  XNOR2_X1 U377 ( .A(G78GAT), .B(G106GAT), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n327), .B(n326), .ZN(n417) );
  XOR2_X1 U379 ( .A(KEYINPUT31), .B(KEYINPUT72), .Z(n329) );
  NAND2_X1 U380 ( .A1(G230GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U382 ( .A(n330), .B(KEYINPUT33), .Z(n334) );
  XNOR2_X1 U383 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U384 ( .A(n334), .B(n333), .ZN(n337) );
  INV_X1 U385 ( .A(n337), .ZN(n335) );
  NAND2_X1 U386 ( .A1(n335), .A2(KEYINPUT32), .ZN(n339) );
  INV_X1 U387 ( .A(KEYINPUT32), .ZN(n336) );
  NAND2_X1 U388 ( .A1(n337), .A2(n336), .ZN(n338) );
  NAND2_X1 U389 ( .A1(n339), .A2(n338), .ZN(n341) );
  XOR2_X1 U390 ( .A(G99GAT), .B(G85GAT), .Z(n368) );
  XNOR2_X1 U391 ( .A(G120GAT), .B(n368), .ZN(n340) );
  XNOR2_X1 U392 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U393 ( .A(KEYINPUT67), .B(G15GAT), .Z(n344) );
  XNOR2_X1 U394 ( .A(G197GAT), .B(G113GAT), .ZN(n343) );
  XNOR2_X1 U395 ( .A(n344), .B(n343), .ZN(n356) );
  XOR2_X1 U396 ( .A(G50GAT), .B(G36GAT), .Z(n348) );
  XNOR2_X1 U397 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U398 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U399 ( .A(G141GAT), .B(G22GAT), .Z(n421) );
  XOR2_X1 U400 ( .A(n349), .B(n421), .Z(n354) );
  XOR2_X1 U401 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n351) );
  NAND2_X1 U402 ( .A1(G229GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U403 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U404 ( .A(KEYINPUT29), .B(n352), .ZN(n353) );
  XNOR2_X1 U405 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U406 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U407 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n358) );
  XNOR2_X1 U408 ( .A(G43GAT), .B(G29GAT), .ZN(n357) );
  XNOR2_X1 U409 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U410 ( .A(KEYINPUT69), .B(n359), .Z(n365) );
  NOR2_X1 U411 ( .A1(n563), .A2(n582), .ZN(n361) );
  XNOR2_X1 U412 ( .A(n361), .B(KEYINPUT46), .ZN(n362) );
  INV_X1 U413 ( .A(n590), .ZN(n496) );
  NOR2_X1 U414 ( .A1(n362), .A2(n496), .ZN(n364) );
  INV_X1 U415 ( .A(KEYINPUT112), .ZN(n363) );
  XNOR2_X1 U416 ( .A(n364), .B(n363), .ZN(n381) );
  INV_X1 U417 ( .A(n365), .ZN(n380) );
  XOR2_X1 U418 ( .A(KEYINPUT11), .B(KEYINPUT66), .Z(n367) );
  XNOR2_X1 U419 ( .A(G106GAT), .B(G92GAT), .ZN(n366) );
  XNOR2_X1 U420 ( .A(n367), .B(n366), .ZN(n372) );
  XOR2_X1 U421 ( .A(KEYINPUT10), .B(n368), .Z(n370) );
  XOR2_X1 U422 ( .A(G50GAT), .B(G162GAT), .Z(n413) );
  XNOR2_X1 U423 ( .A(G134GAT), .B(n413), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U425 ( .A(n372), .B(n371), .Z(n374) );
  NAND2_X1 U426 ( .A1(G232GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U427 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U428 ( .A(n375), .B(KEYINPUT9), .Z(n378) );
  XNOR2_X1 U429 ( .A(n376), .B(KEYINPUT64), .ZN(n377) );
  XNOR2_X1 U430 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U431 ( .A(n380), .B(n379), .Z(n480) );
  NOR2_X1 U432 ( .A1(n381), .A2(n480), .ZN(n383) );
  XOR2_X1 U433 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n386) );
  XOR2_X1 U434 ( .A(n480), .B(KEYINPUT101), .Z(n384) );
  XNOR2_X1 U435 ( .A(n384), .B(KEYINPUT36), .ZN(n494) );
  NAND2_X1 U436 ( .A1(n494), .A2(n496), .ZN(n385) );
  XNOR2_X1 U437 ( .A(n386), .B(n385), .ZN(n388) );
  NAND2_X1 U438 ( .A1(n582), .A2(n586), .ZN(n387) );
  NOR2_X1 U439 ( .A1(n388), .A2(n387), .ZN(n389) );
  NOR2_X1 U440 ( .A1(n390), .A2(n389), .ZN(n391) );
  XNOR2_X1 U441 ( .A(n391), .B(KEYINPUT48), .ZN(n555) );
  NOR2_X1 U442 ( .A1(n529), .A2(n555), .ZN(n392) );
  XNOR2_X1 U443 ( .A(n392), .B(KEYINPUT54), .ZN(n454) );
  XOR2_X1 U444 ( .A(G155GAT), .B(KEYINPUT2), .Z(n394) );
  XNOR2_X1 U445 ( .A(KEYINPUT86), .B(KEYINPUT3), .ZN(n393) );
  XNOR2_X1 U446 ( .A(n394), .B(n393), .ZN(n425) );
  XOR2_X1 U447 ( .A(n425), .B(G1GAT), .Z(n396) );
  NAND2_X1 U448 ( .A1(G225GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U449 ( .A(n396), .B(n395), .ZN(n411) );
  XOR2_X1 U450 ( .A(G85GAT), .B(G162GAT), .Z(n398) );
  XNOR2_X1 U451 ( .A(G29GAT), .B(G148GAT), .ZN(n397) );
  XNOR2_X1 U452 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U453 ( .A(KEYINPUT90), .B(KEYINPUT6), .Z(n400) );
  XNOR2_X1 U454 ( .A(KEYINPUT4), .B(G57GAT), .ZN(n399) );
  XNOR2_X1 U455 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U456 ( .A(n402), .B(n401), .Z(n409) );
  XOR2_X1 U457 ( .A(G120GAT), .B(KEYINPUT0), .Z(n404) );
  XNOR2_X1 U458 ( .A(G113GAT), .B(G134GAT), .ZN(n403) );
  XNOR2_X1 U459 ( .A(n404), .B(n403), .ZN(n436) );
  XOR2_X1 U460 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n406) );
  XNOR2_X1 U461 ( .A(G141GAT), .B(G127GAT), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U463 ( .A(n436), .B(n407), .ZN(n408) );
  XNOR2_X1 U464 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U465 ( .A(n411), .B(n410), .ZN(n527) );
  XOR2_X1 U466 ( .A(n413), .B(n412), .Z(n415) );
  NAND2_X1 U467 ( .A1(G228GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U468 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U469 ( .A(n417), .B(n416), .ZN(n429) );
  XOR2_X1 U470 ( .A(KEYINPUT23), .B(KEYINPUT88), .Z(n419) );
  XNOR2_X1 U471 ( .A(KEYINPUT84), .B(KEYINPUT87), .ZN(n418) );
  XNOR2_X1 U472 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U473 ( .A(n420), .B(KEYINPUT22), .Z(n423) );
  XNOR2_X1 U474 ( .A(n421), .B(G218GAT), .ZN(n422) );
  XNOR2_X1 U475 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U476 ( .A(n424), .B(KEYINPUT89), .Z(n427) );
  XNOR2_X1 U477 ( .A(KEYINPUT24), .B(n425), .ZN(n426) );
  XNOR2_X1 U478 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U479 ( .A(n429), .B(n428), .ZN(n470) );
  AND2_X1 U480 ( .A1(n527), .A2(n470), .ZN(n430) );
  NAND2_X1 U481 ( .A1(n454), .A2(n430), .ZN(n431) );
  XNOR2_X1 U482 ( .A(n431), .B(KEYINPUT55), .ZN(n449) );
  XOR2_X1 U483 ( .A(n433), .B(n432), .Z(n435) );
  XNOR2_X1 U484 ( .A(G190GAT), .B(G99GAT), .ZN(n434) );
  XNOR2_X1 U485 ( .A(n435), .B(n434), .ZN(n440) );
  XOR2_X1 U486 ( .A(n436), .B(G71GAT), .Z(n438) );
  NAND2_X1 U487 ( .A1(G227GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U488 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U489 ( .A(n440), .B(n439), .Z(n448) );
  XOR2_X1 U490 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n442) );
  XNOR2_X1 U491 ( .A(G43GAT), .B(KEYINPUT20), .ZN(n441) );
  XNOR2_X1 U492 ( .A(n442), .B(n441), .ZN(n446) );
  XOR2_X1 U493 ( .A(G176GAT), .B(G183GAT), .Z(n444) );
  XNOR2_X1 U494 ( .A(G169GAT), .B(KEYINPUT81), .ZN(n443) );
  XNOR2_X1 U495 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U496 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U497 ( .A(n448), .B(n447), .Z(n531) );
  INV_X1 U498 ( .A(n531), .ZN(n542) );
  NAND2_X1 U499 ( .A1(n449), .A2(n542), .ZN(n577) );
  NOR2_X1 U500 ( .A1(n590), .A2(n577), .ZN(n452) );
  INV_X1 U501 ( .A(G183GAT), .ZN(n450) );
  NOR2_X1 U502 ( .A1(n470), .A2(n542), .ZN(n453) );
  XOR2_X1 U503 ( .A(n453), .B(KEYINPUT26), .Z(n556) );
  INV_X1 U504 ( .A(n556), .ZN(n467) );
  AND2_X1 U505 ( .A1(n527), .A2(n467), .ZN(n455) );
  NAND2_X1 U506 ( .A1(n455), .A2(n454), .ZN(n456) );
  XNOR2_X1 U507 ( .A(n456), .B(KEYINPUT125), .ZN(n581) );
  NAND2_X1 U508 ( .A1(n581), .A2(n494), .ZN(n457) );
  XNOR2_X1 U509 ( .A(n457), .B(KEYINPUT62), .ZN(n458) );
  XNOR2_X1 U510 ( .A(n458), .B(KEYINPUT127), .ZN(n460) );
  XOR2_X1 U511 ( .A(G218GAT), .B(KEYINPUT126), .Z(n459) );
  XNOR2_X1 U512 ( .A(n460), .B(n459), .ZN(G1355GAT) );
  INV_X1 U513 ( .A(KEYINPUT120), .ZN(n463) );
  NOR2_X1 U514 ( .A1(n577), .A2(n582), .ZN(n461) );
  XNOR2_X1 U515 ( .A(G169GAT), .B(n461), .ZN(n462) );
  XNOR2_X1 U516 ( .A(n463), .B(n462), .ZN(G1348GAT) );
  INV_X1 U517 ( .A(n582), .ZN(n515) );
  AND2_X1 U518 ( .A1(n515), .A2(n586), .ZN(n464) );
  XOR2_X1 U519 ( .A(KEYINPUT75), .B(n464), .Z(n498) );
  XNOR2_X1 U520 ( .A(KEYINPUT27), .B(n506), .ZN(n468) );
  INV_X1 U521 ( .A(n527), .ZN(n501) );
  NAND2_X1 U522 ( .A1(n468), .A2(n501), .ZN(n465) );
  XOR2_X1 U523 ( .A(KEYINPUT92), .B(n465), .Z(n557) );
  XOR2_X1 U524 ( .A(n470), .B(KEYINPUT28), .Z(n512) );
  INV_X1 U525 ( .A(n512), .ZN(n535) );
  NAND2_X1 U526 ( .A1(n557), .A2(n535), .ZN(n541) );
  NOR2_X1 U527 ( .A1(n542), .A2(n541), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n466), .B(KEYINPUT93), .ZN(n479) );
  NAND2_X1 U529 ( .A1(n468), .A2(n467), .ZN(n476) );
  NOR2_X1 U530 ( .A1(n531), .A2(n529), .ZN(n469) );
  XOR2_X1 U531 ( .A(KEYINPUT94), .B(n469), .Z(n471) );
  NAND2_X1 U532 ( .A1(n471), .A2(n470), .ZN(n474) );
  XNOR2_X1 U533 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n472) );
  XNOR2_X1 U534 ( .A(n472), .B(KEYINPUT25), .ZN(n473) );
  XNOR2_X1 U535 ( .A(n474), .B(n473), .ZN(n475) );
  NAND2_X1 U536 ( .A1(n476), .A2(n475), .ZN(n477) );
  NAND2_X1 U537 ( .A1(n477), .A2(n527), .ZN(n478) );
  NAND2_X1 U538 ( .A1(n479), .A2(n478), .ZN(n493) );
  INV_X1 U539 ( .A(n480), .ZN(n578) );
  NAND2_X1 U540 ( .A1(n578), .A2(n496), .ZN(n481) );
  XOR2_X1 U541 ( .A(KEYINPUT16), .B(n481), .Z(n482) );
  AND2_X1 U542 ( .A1(n493), .A2(n482), .ZN(n516) );
  NAND2_X1 U543 ( .A1(n498), .A2(n516), .ZN(n491) );
  NOR2_X1 U544 ( .A1(n527), .A2(n491), .ZN(n484) );
  XNOR2_X1 U545 ( .A(KEYINPUT97), .B(KEYINPUT34), .ZN(n483) );
  XNOR2_X1 U546 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U547 ( .A(G1GAT), .B(n485), .ZN(G1324GAT) );
  NOR2_X1 U548 ( .A1(n529), .A2(n491), .ZN(n486) );
  XOR2_X1 U549 ( .A(KEYINPUT98), .B(n486), .Z(n487) );
  XNOR2_X1 U550 ( .A(G8GAT), .B(n487), .ZN(G1325GAT) );
  NOR2_X1 U551 ( .A1(n531), .A2(n491), .ZN(n489) );
  XNOR2_X1 U552 ( .A(KEYINPUT35), .B(KEYINPUT99), .ZN(n488) );
  XNOR2_X1 U553 ( .A(n489), .B(n488), .ZN(n490) );
  XOR2_X1 U554 ( .A(G15GAT), .B(n490), .Z(G1326GAT) );
  NOR2_X1 U555 ( .A1(n535), .A2(n491), .ZN(n492) );
  XOR2_X1 U556 ( .A(G22GAT), .B(n492), .Z(G1327GAT) );
  XOR2_X1 U557 ( .A(G29GAT), .B(KEYINPUT100), .Z(n503) );
  XOR2_X1 U558 ( .A(KEYINPUT38), .B(KEYINPUT102), .Z(n500) );
  NAND2_X1 U559 ( .A1(n494), .A2(n493), .ZN(n495) );
  NOR2_X1 U560 ( .A1(n496), .A2(n495), .ZN(n497) );
  XOR2_X1 U561 ( .A(KEYINPUT37), .B(n497), .Z(n526) );
  NAND2_X1 U562 ( .A1(n498), .A2(n526), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(n513) );
  NAND2_X1 U564 ( .A1(n513), .A2(n501), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(n505) );
  XOR2_X1 U566 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n504) );
  XNOR2_X1 U567 ( .A(n505), .B(n504), .ZN(G1328GAT) );
  NAND2_X1 U568 ( .A1(n506), .A2(n513), .ZN(n507) );
  XNOR2_X1 U569 ( .A(G36GAT), .B(n507), .ZN(G1329GAT) );
  XNOR2_X1 U570 ( .A(G43GAT), .B(KEYINPUT104), .ZN(n511) );
  XOR2_X1 U571 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n509) );
  NAND2_X1 U572 ( .A1(n513), .A2(n542), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n511), .B(n510), .ZN(G1330GAT) );
  NAND2_X1 U575 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U576 ( .A(n514), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U577 ( .A(n563), .B(KEYINPUT106), .ZN(n570) );
  NOR2_X1 U578 ( .A1(n515), .A2(n570), .ZN(n525) );
  NAND2_X1 U579 ( .A1(n525), .A2(n516), .ZN(n522) );
  NOR2_X1 U580 ( .A1(n527), .A2(n522), .ZN(n517) );
  XOR2_X1 U581 ( .A(G57GAT), .B(n517), .Z(n518) );
  XNOR2_X1 U582 ( .A(KEYINPUT42), .B(n518), .ZN(G1332GAT) );
  NOR2_X1 U583 ( .A1(n529), .A2(n522), .ZN(n520) );
  XNOR2_X1 U584 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(G1333GAT) );
  NOR2_X1 U586 ( .A1(n531), .A2(n522), .ZN(n521) );
  XOR2_X1 U587 ( .A(G71GAT), .B(n521), .Z(G1334GAT) );
  NOR2_X1 U588 ( .A1(n535), .A2(n522), .ZN(n524) );
  XNOR2_X1 U589 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n523) );
  XNOR2_X1 U590 ( .A(n524), .B(n523), .ZN(G1335GAT) );
  NAND2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n534) );
  NOR2_X1 U592 ( .A1(n527), .A2(n534), .ZN(n528) );
  XOR2_X1 U593 ( .A(G85GAT), .B(n528), .Z(G1336GAT) );
  NOR2_X1 U594 ( .A1(n529), .A2(n534), .ZN(n530) );
  XOR2_X1 U595 ( .A(G92GAT), .B(n530), .Z(G1337GAT) );
  NOR2_X1 U596 ( .A1(n531), .A2(n534), .ZN(n532) );
  XOR2_X1 U597 ( .A(KEYINPUT108), .B(n532), .Z(n533) );
  XNOR2_X1 U598 ( .A(G99GAT), .B(n533), .ZN(G1338GAT) );
  NOR2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n540) );
  XOR2_X1 U600 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n537) );
  XNOR2_X1 U601 ( .A(G106GAT), .B(KEYINPUT110), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U603 ( .A(KEYINPUT109), .B(n538), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(G1339GAT) );
  NOR2_X1 U605 ( .A1(n555), .A2(n541), .ZN(n543) );
  NAND2_X1 U606 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U607 ( .A(n544), .B(KEYINPUT114), .ZN(n551) );
  NOR2_X1 U608 ( .A1(n551), .A2(n582), .ZN(n545) );
  XOR2_X1 U609 ( .A(G113GAT), .B(n545), .Z(G1340GAT) );
  NOR2_X1 U610 ( .A1(n551), .A2(n570), .ZN(n547) );
  XNOR2_X1 U611 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U613 ( .A(G120GAT), .B(n548), .Z(G1341GAT) );
  NOR2_X1 U614 ( .A1(n590), .A2(n551), .ZN(n549) );
  XOR2_X1 U615 ( .A(KEYINPUT50), .B(n549), .Z(n550) );
  XNOR2_X1 U616 ( .A(G127GAT), .B(n550), .ZN(G1342GAT) );
  XNOR2_X1 U617 ( .A(KEYINPUT116), .B(KEYINPUT51), .ZN(n553) );
  NOR2_X1 U618 ( .A1(n578), .A2(n551), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G134GAT), .B(n554), .ZN(G1343GAT) );
  NOR2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n558) );
  NAND2_X1 U622 ( .A1(n558), .A2(n557), .ZN(n568) );
  NOR2_X1 U623 ( .A1(n582), .A2(n568), .ZN(n560) );
  XNOR2_X1 U624 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(G1344GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT52), .B(KEYINPUT118), .Z(n562) );
  XNOR2_X1 U627 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n565) );
  NOR2_X1 U629 ( .A1(n563), .A2(n568), .ZN(n564) );
  XOR2_X1 U630 ( .A(n565), .B(n564), .Z(G1345GAT) );
  NOR2_X1 U631 ( .A1(n590), .A2(n568), .ZN(n567) );
  XNOR2_X1 U632 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1346GAT) );
  NOR2_X1 U634 ( .A1(n578), .A2(n568), .ZN(n569) );
  XOR2_X1 U635 ( .A(G162GAT), .B(n569), .Z(G1347GAT) );
  NOR2_X1 U636 ( .A1(n577), .A2(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n574) );
  XOR2_X1 U639 ( .A(KEYINPUT56), .B(KEYINPUT121), .Z(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1349GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n576) );
  XNOR2_X1 U642 ( .A(G190GAT), .B(KEYINPUT124), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n576), .B(n575), .ZN(n580) );
  NOR2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U645 ( .A(n580), .B(n579), .Z(G1351GAT) );
  INV_X1 U646 ( .A(n581), .ZN(n589) );
  NOR2_X1 U647 ( .A1(n582), .A2(n589), .ZN(n584) );
  XNOR2_X1 U648 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(G197GAT), .B(n585), .ZN(G1352GAT) );
  NOR2_X1 U651 ( .A1(n586), .A2(n589), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1353GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U655 ( .A(G211GAT), .B(n591), .Z(G1354GAT) );
endmodule

