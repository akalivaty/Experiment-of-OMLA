//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n547, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n601, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1138, new_n1139;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT67), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT68), .Z(G325));
  XOR2_X1   g031(.A(G325), .B(KEYINPUT69), .Z(G261));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n452), .A2(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT70), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(KEYINPUT71), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT71), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(new_n465), .A3(G2104), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n463), .A2(new_n466), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G137), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n462), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT72), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n473), .B(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n465), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n468), .ZN(new_n478));
  INV_X1    g053(.A(G125), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n471), .A2(new_n475), .A3(new_n481), .ZN(G160));
  AND2_X1   g057(.A1(new_n466), .A2(new_n468), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n483), .A2(G2105), .A3(new_n463), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n467), .A2(G112), .ZN(new_n486));
  OAI21_X1  g061(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n487));
  OAI22_X1  g062(.A1(new_n484), .A2(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(G136), .B2(new_n470), .ZN(G162));
  XNOR2_X1  g064(.A(KEYINPUT73), .B(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n467), .A2(G138), .ZN(new_n491));
  NOR3_X1   g066(.A1(new_n478), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n483), .A2(G138), .A3(new_n467), .A4(new_n463), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(KEYINPUT4), .ZN(new_n494));
  OAI21_X1  g069(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G126), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n484), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT74), .B1(new_n494), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT4), .B1(new_n469), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n478), .A2(new_n491), .ZN(new_n504));
  INV_X1    g079(.A(new_n490), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT74), .ZN(new_n508));
  AND4_X1   g083(.A1(G2105), .A2(new_n463), .A3(new_n466), .A4(new_n468), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n497), .B1(new_n509), .B2(G126), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n507), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n501), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(G164));
  NAND2_X1  g088(.A1(KEYINPUT75), .A2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(KEYINPUT75), .A2(KEYINPUT5), .A3(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT6), .B(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G50), .ZN(new_n526));
  OAI22_X1  g101(.A1(new_n523), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n521), .A2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  INV_X1    g106(.A(G89), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n523), .B2(new_n532), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT76), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n522), .A2(G543), .ZN(new_n535));
  AND2_X1   g110(.A1(G63), .A2(G651), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n535), .A2(G51), .B1(new_n518), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(KEYINPUT77), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT77), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n534), .A2(new_n540), .A3(new_n537), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n541), .ZN(G168));
  AOI22_X1  g117(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n520), .ZN(new_n544));
  INV_X1    g119(.A(G90), .ZN(new_n545));
  INV_X1    g120(.A(G52), .ZN(new_n546));
  OAI22_X1  g121(.A1(new_n523), .A2(new_n545), .B1(new_n525), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n544), .A2(new_n547), .ZN(G171));
  AOI22_X1  g123(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n520), .ZN(new_n550));
  INV_X1    g125(.A(G81), .ZN(new_n551));
  XOR2_X1   g126(.A(KEYINPUT78), .B(G43), .Z(new_n552));
  OAI22_X1  g127(.A1(new_n523), .A2(new_n551), .B1(new_n525), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  AOI22_X1  g135(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n561), .A2(new_n520), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT79), .Z(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OR3_X1    g139(.A1(new_n525), .A2(KEYINPUT9), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT9), .B1(new_n525), .B2(new_n564), .ZN(new_n566));
  INV_X1    g141(.A(new_n523), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n565), .A2(new_n566), .B1(G91), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n563), .A2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  INV_X1    g145(.A(G168), .ZN(G286));
  NAND2_X1  g146(.A1(new_n567), .A2(G87), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n535), .A2(G49), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  AOI22_X1  g150(.A1(new_n518), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(new_n520), .ZN(new_n577));
  INV_X1    g152(.A(G86), .ZN(new_n578));
  INV_X1    g153(.A(G48), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n523), .A2(new_n578), .B1(new_n525), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n583), .A2(new_n520), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT80), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n567), .A2(G85), .B1(new_n535), .B2(G47), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n567), .A2(G92), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT10), .Z(new_n590));
  AOI22_X1  g165(.A1(new_n518), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G54), .ZN(new_n592));
  OAI22_X1  g167(.A1(new_n591), .A2(new_n520), .B1(new_n525), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT81), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n593), .B(new_n594), .ZN(new_n595));
  AND2_X1   g170(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n588), .B1(new_n596), .B2(G868), .ZN(G284));
  OAI21_X1  g172(.A(new_n588), .B1(new_n596), .B2(G868), .ZN(G321));
  MUX2_X1   g173(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g174(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n596), .B1(new_n601), .B2(G860), .ZN(G148));
  NAND2_X1  g177(.A1(new_n596), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g181(.A1(G99), .A2(G2105), .ZN(new_n607));
  OAI211_X1 g182(.A(new_n607), .B(G2104), .C1(G111), .C2(new_n467), .ZN(new_n608));
  INV_X1    g183(.A(G123), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n484), .B2(new_n609), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(G135), .B2(new_n470), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n612), .A2(G2096), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n612), .A2(G2096), .ZN(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT82), .B(KEYINPUT13), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2100), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n617));
  XOR2_X1   g192(.A(new_n617), .B(KEYINPUT12), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n616), .B(new_n618), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n613), .A2(new_n614), .A3(new_n619), .ZN(G156));
  XNOR2_X1  g195(.A(KEYINPUT15), .B(G2435), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2438), .Z(new_n622));
  XNOR2_X1  g197(.A(G2427), .B(G2430), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(KEYINPUT14), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT83), .ZN(new_n626));
  INV_X1    g201(.A(new_n622), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(new_n623), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2443), .B(G2446), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G1341), .B(G1348), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2451), .B(G2454), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n632), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(new_n636), .A3(G14), .ZN(new_n637));
  INV_X1    g212(.A(new_n637), .ZN(G401));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  XNOR2_X1  g214(.A(G2067), .B(G2678), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2072), .B(G2078), .Z(new_n642));
  NOR2_X1   g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT84), .B(KEYINPUT18), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT85), .B(KEYINPUT17), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n642), .B(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n639), .ZN(new_n648));
  INV_X1    g223(.A(new_n640), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n648), .A2(new_n642), .A3(new_n649), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(new_n641), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n645), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT86), .ZN(new_n654));
  XOR2_X1   g229(.A(G2096), .B(G2100), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(G227));
  XNOR2_X1  g231(.A(G1971), .B(G1976), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT87), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n660), .A2(new_n662), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n658), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(new_n663), .A3(new_n658), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n664), .B1(new_n663), .B2(new_n658), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1981), .B(G1986), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G229));
  INV_X1    g252(.A(G16), .ZN(new_n678));
  NOR2_X1   g253(.A1(G286), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT98), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g256(.A(KEYINPUT98), .B1(G16), .B2(G21), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n681), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(KEYINPUT99), .B(G1966), .Z(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT100), .ZN(new_n687));
  NAND2_X1  g262(.A1(G115), .A2(G2104), .ZN(new_n688));
  INV_X1    g263(.A(G127), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n688), .B1(new_n478), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G2105), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT95), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n467), .A2(G103), .A3(G2104), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT25), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(new_n470), .B2(G139), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n698), .B2(G33), .ZN(new_n700));
  INV_X1    g275(.A(G2072), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT96), .Z(new_n703));
  INV_X1    g278(.A(G34), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(KEYINPUT24), .ZN(new_n705));
  AOI21_X1  g280(.A(G29), .B1(new_n704), .B2(KEYINPUT24), .ZN(new_n706));
  AOI22_X1  g281(.A1(G160), .A2(G29), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n707), .A2(G2084), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n554), .A2(new_n678), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n678), .B2(G19), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  OAI22_X1  g286(.A1(new_n711), .A2(G1341), .B1(G2084), .B2(new_n707), .ZN(new_n712));
  AOI211_X1 g287(.A(new_n708), .B(new_n712), .C1(G1341), .C2(new_n711), .ZN(new_n713));
  NOR2_X1   g288(.A1(G171), .A2(new_n678), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G5), .B2(new_n678), .ZN(new_n715));
  INV_X1    g290(.A(G1961), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT101), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n698), .A2(G26), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  INV_X1    g295(.A(G104), .ZN(new_n721));
  AND3_X1   g296(.A1(new_n721), .A2(new_n467), .A3(KEYINPUT94), .ZN(new_n722));
  AOI21_X1  g297(.A(KEYINPUT94), .B1(new_n721), .B2(new_n467), .ZN(new_n723));
  OAI221_X1 g298(.A(G2104), .B1(G116), .B2(new_n467), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G128), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n484), .B2(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G140), .B2(new_n470), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n720), .B1(new_n727), .B2(new_n698), .ZN(new_n728));
  AOI22_X1  g303(.A1(new_n700), .A2(new_n701), .B1(G2067), .B2(new_n728), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n715), .A2(new_n716), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n728), .A2(G2067), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n612), .A2(new_n698), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT31), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n733), .A2(G11), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(G11), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT30), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n736), .A2(G28), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n698), .B1(new_n736), .B2(G28), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n734), .B(new_n735), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  NOR4_X1   g314(.A1(new_n730), .A2(new_n731), .A3(new_n732), .A4(new_n739), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n713), .A2(new_n718), .A3(new_n729), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n678), .A2(G20), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT23), .Z(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G299), .B2(G16), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(G1956), .Z(new_n745));
  NAND2_X1  g320(.A1(new_n698), .A2(G27), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G164), .B2(new_n698), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G2078), .ZN(new_n748));
  NOR4_X1   g323(.A1(new_n703), .A2(new_n741), .A3(new_n745), .A4(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(G4), .A2(G16), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n596), .B2(G16), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT93), .B(G1348), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n698), .A2(G35), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G162), .B2(new_n698), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT29), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2090), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n698), .A2(G32), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n470), .A2(G141), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n509), .A2(G129), .ZN(new_n760));
  NAND3_X1  g335(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT26), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  AOI22_X1  g339(.A1(new_n763), .A2(new_n764), .B1(G105), .B2(new_n472), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n759), .A2(new_n760), .A3(new_n765), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n766), .A2(KEYINPUT97), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(KEYINPUT97), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n758), .B1(new_n770), .B2(new_n698), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT27), .Z(new_n772));
  AOI211_X1 g347(.A(new_n753), .B(new_n757), .C1(G1996), .C2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n772), .ZN(new_n774));
  INV_X1    g349(.A(G1996), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n774), .A2(new_n775), .B1(new_n683), .B2(new_n685), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n687), .A2(new_n749), .A3(new_n773), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n678), .A2(G22), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G166), .B2(new_n678), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(G1971), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n678), .A2(G23), .ZN(new_n781));
  INV_X1    g356(.A(G288), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(new_n678), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT90), .Z(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT33), .B(G1976), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n780), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n678), .A2(G6), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n581), .B2(new_n678), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT89), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT32), .B(G1981), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n786), .B(new_n791), .C1(new_n784), .C2(new_n785), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT91), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n792), .A2(new_n793), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n794), .A2(KEYINPUT34), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT92), .ZN(new_n797));
  AOI21_X1  g372(.A(KEYINPUT34), .B1(new_n794), .B2(new_n795), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n698), .A2(G25), .ZN(new_n799));
  INV_X1    g374(.A(G119), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n467), .A2(G107), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n484), .A2(new_n800), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G131), .B2(new_n470), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n799), .B1(new_n804), .B2(new_n698), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT35), .B(G1991), .Z(new_n806));
  XOR2_X1   g381(.A(new_n805), .B(new_n806), .Z(new_n807));
  NOR2_X1   g382(.A1(G16), .A2(G24), .ZN(new_n808));
  INV_X1    g383(.A(G290), .ZN(new_n809));
  AOI21_X1  g384(.A(new_n808), .B1(new_n809), .B2(G16), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1986), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n798), .A2(new_n807), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n797), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(KEYINPUT36), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT36), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n797), .A2(new_n812), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n777), .B1(new_n814), .B2(new_n816), .ZN(G311));
  INV_X1    g392(.A(G311), .ZN(G150));
  AOI22_X1  g393(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(new_n520), .ZN(new_n820));
  INV_X1    g395(.A(G93), .ZN(new_n821));
  INV_X1    g396(.A(G55), .ZN(new_n822));
  OAI22_X1  g397(.A1(new_n523), .A2(new_n821), .B1(new_n525), .B2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT102), .ZN(new_n824));
  OR3_X1    g399(.A1(new_n820), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n554), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n824), .B1(new_n820), .B2(new_n823), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n825), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n554), .B1(new_n820), .B2(new_n823), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT103), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT103), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n828), .A2(new_n832), .A3(new_n829), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT38), .Z(new_n835));
  INV_X1    g410(.A(new_n596), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n836), .A2(new_n601), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n835), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT39), .ZN(new_n839));
  AOI21_X1  g414(.A(G860), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n825), .A2(new_n827), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G860), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT37), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n841), .A2(new_n844), .ZN(G145));
  NAND2_X1  g420(.A1(new_n507), .A2(new_n510), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT104), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT104), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n507), .A2(new_n848), .A3(new_n510), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n727), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n769), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT105), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n853), .B1(new_n696), .B2(KEYINPUT106), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(KEYINPUT105), .B2(new_n697), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n851), .B(new_n770), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n858), .A2(new_n855), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n509), .A2(G130), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n467), .A2(G118), .ZN(new_n861));
  OAI21_X1  g436(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n863), .B1(G142), .B2(new_n470), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(new_n618), .Z(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n804), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n857), .A2(new_n859), .A3(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n867), .B1(new_n859), .B2(new_n857), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(G162), .B(new_n611), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(G160), .Z(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(G37), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n870), .A2(new_n873), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n875), .A2(KEYINPUT107), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT107), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n870), .A2(new_n877), .A3(new_n873), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n874), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g455(.A(G290), .B(new_n782), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT109), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(G305), .B(G303), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n881), .A2(new_n882), .ZN(new_n886));
  MUX2_X1   g461(.A(new_n885), .B(new_n884), .S(new_n886), .Z(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT42), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n596), .A2(G299), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT108), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n596), .A2(G299), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n596), .A2(KEYINPUT108), .A3(G299), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(KEYINPUT41), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT41), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n889), .A2(new_n895), .A3(new_n891), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n892), .A2(new_n893), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n834), .B(new_n603), .ZN(new_n899));
  MUX2_X1   g474(.A(new_n897), .B(new_n898), .S(new_n899), .Z(new_n900));
  XNOR2_X1  g475(.A(new_n888), .B(new_n900), .ZN(new_n901));
  MUX2_X1   g476(.A(new_n842), .B(new_n901), .S(G868), .Z(G295));
  MUX2_X1   g477(.A(new_n842), .B(new_n901), .S(G868), .Z(G331));
  INV_X1    g478(.A(KEYINPUT110), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n539), .A2(new_n904), .A3(new_n541), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n905), .B1(new_n831), .B2(new_n833), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(G301), .B1(G168), .B2(KEYINPUT110), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n831), .A2(new_n905), .A3(new_n833), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n908), .ZN(new_n911));
  INV_X1    g486(.A(new_n909), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n911), .B1(new_n912), .B2(new_n906), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n895), .B1(new_n910), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n889), .A2(new_n891), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n887), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n898), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n916), .B1(new_n917), .B2(new_n914), .ZN(new_n918));
  NOR3_X1   g493(.A1(new_n912), .A2(new_n911), .A3(new_n906), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n908), .B1(new_n907), .B2(new_n909), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n897), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n910), .A2(new_n913), .A3(new_n898), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(G37), .B1(new_n923), .B2(new_n887), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n918), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n887), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n927), .A2(new_n921), .A3(new_n922), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n924), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n926), .B1(new_n929), .B2(new_n925), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n918), .A2(new_n924), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT111), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT112), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT111), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n918), .A2(new_n924), .A3(new_n936), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT43), .A4(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n931), .B1(new_n929), .B2(new_n925), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n925), .B1(new_n933), .B2(KEYINPUT111), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n935), .B1(new_n941), .B2(new_n937), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n932), .B1(new_n940), .B2(new_n942), .ZN(G397));
  INV_X1    g518(.A(G1384), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n850), .A2(new_n944), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n945), .A2(KEYINPUT45), .ZN(new_n946));
  AND4_X1   g521(.A1(G40), .A2(new_n471), .A3(new_n475), .A4(new_n481), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n770), .A2(new_n775), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n769), .A2(G1996), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n727), .B(G2067), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n804), .B(new_n806), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n949), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G1986), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n809), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(KEYINPUT113), .B1(G290), .B2(G1986), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n957), .B(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n949), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n955), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n961), .B(KEYINPUT114), .Z(new_n962));
  INV_X1    g537(.A(KEYINPUT51), .ZN(new_n963));
  AND3_X1   g538(.A1(new_n507), .A2(new_n508), .A3(new_n510), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n508), .B1(new_n507), .B2(new_n510), .ZN(new_n965));
  OAI211_X1 g540(.A(KEYINPUT45), .B(new_n944), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT116), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT116), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n512), .A2(new_n968), .A3(KEYINPUT45), .A4(new_n944), .ZN(new_n969));
  AOI21_X1  g544(.A(G1384), .B1(new_n507), .B2(new_n510), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n947), .B1(new_n970), .B2(KEYINPUT45), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n967), .A2(new_n969), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n684), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT117), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n971), .B1(new_n966), .B2(KEYINPUT116), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n685), .B1(new_n977), .B2(new_n969), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(KEYINPUT117), .ZN(new_n979));
  INV_X1    g554(.A(new_n970), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n947), .B1(new_n980), .B2(KEYINPUT50), .ZN(new_n981));
  AOI21_X1  g556(.A(G1384), .B1(new_n501), .B2(new_n511), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n981), .B1(new_n983), .B2(KEYINPUT50), .ZN(new_n984));
  XOR2_X1   g559(.A(KEYINPUT118), .B(G2084), .Z(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n976), .A2(new_n979), .A3(new_n986), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n963), .B(G8), .C1(new_n987), .C2(G286), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n986), .B1(new_n978), .B2(KEYINPUT117), .ZN(new_n989));
  AOI211_X1 g564(.A(new_n975), .B(new_n685), .C1(new_n977), .C2(new_n969), .ZN(new_n990));
  OAI21_X1  g565(.A(G8), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G8), .ZN(new_n992));
  NOR2_X1   g567(.A1(G168), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n991), .A2(KEYINPUT51), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT122), .B1(new_n987), .B2(new_n993), .ZN(new_n996));
  OAI211_X1 g571(.A(KEYINPUT122), .B(new_n993), .C1(new_n989), .C2(new_n990), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  OAI211_X1 g573(.A(new_n988), .B(new_n995), .C1(new_n996), .C2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT123), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT62), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT122), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n989), .A2(new_n990), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1002), .B1(new_n1003), .B2(new_n994), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n997), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT123), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1005), .A2(new_n1006), .A3(new_n988), .A4(new_n995), .ZN(new_n1007));
  AND3_X1   g582(.A1(new_n1000), .A2(new_n1001), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1001), .B1(new_n1000), .B2(new_n1007), .ZN(new_n1009));
  OR2_X1    g584(.A1(G305), .A2(G1981), .ZN(new_n1010));
  NAND2_X1  g585(.A1(G305), .A2(G1981), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT49), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n948), .A2(new_n980), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1015), .A2(new_n992), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1010), .A2(KEYINPUT49), .A3(new_n1011), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n782), .A2(G1976), .ZN(new_n1019));
  INV_X1    g594(.A(G1976), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(G288), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1016), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1018), .B1(new_n1022), .B2(KEYINPUT115), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1024), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1023), .B1(new_n1027), .B2(new_n1022), .ZN(new_n1028));
  NAND2_X1  g603(.A1(G303), .A2(G8), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(KEYINPUT55), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n847), .A2(KEYINPUT45), .A3(new_n944), .A4(new_n849), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1031), .B(new_n947), .C1(new_n982), .C2(KEYINPUT45), .ZN(new_n1032));
  INV_X1    g607(.A(G1971), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n947), .B1(new_n970), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1035), .B1(new_n982), .B2(new_n1034), .ZN(new_n1036));
  INV_X1    g611(.A(G2090), .ZN(new_n1037));
  AOI22_X1  g612(.A1(new_n1032), .A2(new_n1033), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1030), .B1(new_n1038), .B2(new_n992), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n984), .A2(new_n1037), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n992), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1030), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1028), .A2(new_n1039), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1047), .B1(new_n1032), .B2(G2078), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT124), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n948), .B1(new_n1034), .B2(new_n970), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n982), .B2(new_n1034), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1048), .A2(new_n1049), .B1(new_n716), .B2(new_n1051), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1053));
  OR3_X1    g628(.A1(new_n973), .A2(new_n1047), .A3(G2078), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1046), .A2(G171), .A3(new_n1055), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1008), .A2(new_n1009), .A3(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(G171), .B(KEYINPUT54), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1053), .A2(new_n1052), .A3(new_n1054), .A4(new_n1059), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n948), .A2(KEYINPUT125), .ZN(new_n1061));
  AOI211_X1 g636(.A(new_n1047), .B(G2078), .C1(new_n948), .C2(KEYINPUT125), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n946), .A2(new_n1031), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1053), .A2(new_n1063), .A3(new_n1052), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1060), .B1(new_n1064), .B2(new_n1059), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(new_n1046), .ZN(new_n1066));
  XOR2_X1   g641(.A(KEYINPUT58), .B(G1341), .Z(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n948), .B2(new_n980), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n1032), .B2(G1996), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT121), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1071), .B(new_n1068), .C1(new_n1032), .C2(G1996), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n826), .B1(new_n1070), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n1074));
  XNOR2_X1  g649(.A(new_n1073), .B(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(G1348), .ZN(new_n1076));
  INV_X1    g651(.A(G2067), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1051), .A2(new_n1076), .B1(new_n1077), .B2(new_n1015), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(new_n596), .ZN(new_n1079));
  OR2_X1    g654(.A1(new_n1079), .A2(KEYINPUT60), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT56), .B(G2072), .ZN(new_n1081));
  INV_X1    g656(.A(new_n1081), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n1032), .A2(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g658(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n1084));
  XNOR2_X1  g659(.A(G299), .B(new_n1084), .ZN(new_n1085));
  OR2_X1    g660(.A1(new_n1036), .A2(G1956), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1085), .ZN(new_n1088));
  OAI22_X1  g663(.A1(new_n1032), .A2(new_n1082), .B1(new_n1036), .B2(G1956), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1087), .A2(new_n1090), .A3(KEYINPUT61), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1015), .A2(new_n1077), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(new_n984), .B2(G1348), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n836), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1094), .A2(new_n1079), .A3(KEYINPUT60), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1080), .A2(new_n1091), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT61), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1087), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1090), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1075), .A2(new_n1096), .A3(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1078), .A2(new_n836), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1099), .B1(new_n1087), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1066), .B1(new_n1101), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1000), .A2(new_n1007), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1028), .A2(new_n1043), .A3(new_n1042), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1018), .A2(new_n1020), .A3(new_n782), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1010), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1016), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1028), .A2(new_n1044), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n987), .A2(G8), .A3(G168), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT63), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1114));
  OR3_X1    g689(.A1(new_n1112), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  XOR2_X1   g690(.A(KEYINPUT119), .B(KEYINPUT63), .Z(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(new_n1045), .B2(new_n1113), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1111), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1106), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n962), .B1(new_n1057), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n960), .B1(new_n770), .B2(new_n952), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT46), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n960), .A2(new_n1122), .A3(G1996), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT46), .B1(new_n949), .B2(new_n775), .ZN(new_n1124));
  NOR3_X1   g699(.A1(new_n1121), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n1126));
  XNOR2_X1  g701(.A(new_n1125), .B(new_n1126), .ZN(new_n1127));
  XOR2_X1   g702(.A(new_n955), .B(KEYINPUT127), .Z(new_n1128));
  NAND3_X1  g703(.A1(new_n949), .A2(new_n956), .A3(new_n809), .ZN(new_n1129));
  XOR2_X1   g704(.A(new_n1129), .B(KEYINPUT48), .Z(new_n1130));
  NAND2_X1  g705(.A1(new_n804), .A2(new_n806), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n953), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1132), .B1(new_n1077), .B2(new_n727), .ZN(new_n1133));
  OAI22_X1  g708(.A1(new_n1128), .A2(new_n1130), .B1(new_n960), .B2(new_n1133), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1127), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1120), .A2(new_n1135), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g711(.A(G319), .ZN(new_n1138));
  NOR4_X1   g712(.A1(G401), .A2(new_n1138), .A3(G227), .A4(G229), .ZN(new_n1139));
  NAND3_X1  g713(.A1(new_n879), .A2(new_n930), .A3(new_n1139), .ZN(G225));
  INV_X1    g714(.A(G225), .ZN(G308));
endmodule


