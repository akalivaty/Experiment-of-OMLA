//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:12 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n188), .A2(G143), .A3(G214), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  AOI21_X1  g004(.A(G143), .B1(new_n188), .B2(G214), .ZN(new_n191));
  OAI211_X1 g005(.A(KEYINPUT18), .B(G131), .C1(new_n190), .C2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G125), .B(G140), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT79), .A2(G125), .ZN(new_n196));
  INV_X1    g010(.A(G140), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(KEYINPUT79), .A2(G125), .A3(G140), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n198), .A2(G146), .A3(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n195), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(new_n191), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT18), .A2(G131), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n189), .A3(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n192), .A2(new_n201), .A3(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(G113), .B(G122), .ZN(new_n206));
  XNOR2_X1  g020(.A(new_n206), .B(G104), .ZN(new_n207));
  XNOR2_X1  g021(.A(new_n207), .B(KEYINPUT94), .ZN(new_n208));
  AND3_X1   g022(.A1(KEYINPUT79), .A2(G125), .A3(G140), .ZN(new_n209));
  AOI21_X1  g023(.A(G140), .B1(KEYINPUT79), .B2(G125), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT16), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT16), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n212), .A2(new_n197), .A3(G125), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT80), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT80), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n215), .A2(new_n212), .A3(new_n197), .A4(G125), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n211), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(new_n194), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT82), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n217), .A2(KEYINPUT82), .A3(new_n194), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n211), .A2(G146), .A3(new_n214), .A4(new_n216), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT81), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n222), .A2(new_n223), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n220), .B(new_n221), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(KEYINPUT64), .A2(G131), .ZN(new_n227));
  AND2_X1   g041(.A1(KEYINPUT64), .A2(G131), .ZN(new_n228));
  OAI22_X1  g042(.A1(new_n190), .A2(new_n191), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT17), .ZN(new_n230));
  OR2_X1    g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n228), .A2(new_n227), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n202), .A2(new_n232), .A3(new_n189), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n229), .A2(new_n233), .A3(new_n230), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n205), .B(new_n208), .C1(new_n226), .C2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n207), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n217), .A2(KEYINPUT82), .A3(new_n194), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT82), .B1(new_n217), .B2(new_n194), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(new_n222), .B(new_n223), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n241), .A2(new_n242), .A3(new_n231), .A4(new_n234), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n238), .B1(new_n243), .B2(new_n205), .ZN(new_n244));
  OAI211_X1 g058(.A(KEYINPUT95), .B(new_n187), .C1(new_n237), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G475), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n205), .B1(new_n226), .B2(new_n235), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n207), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n236), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT95), .B1(new_n249), .B2(new_n187), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT20), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT19), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n193), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n198), .A2(KEYINPUT19), .A3(new_n199), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(new_n194), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT93), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n255), .B(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n229), .A2(new_n233), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n222), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n205), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n207), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n236), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(G475), .A2(G902), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n251), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AND3_X1   g078(.A1(new_n262), .A2(new_n251), .A3(new_n263), .ZN(new_n265));
  OAI22_X1  g079(.A1(new_n246), .A2(new_n250), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G143), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G128), .ZN(new_n268));
  INV_X1    g082(.A(G128), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(G143), .ZN(new_n270));
  INV_X1    g084(.A(G134), .ZN(new_n271));
  AND3_X1   g085(.A1(new_n268), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G122), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G116), .ZN(new_n274));
  INV_X1    g088(.A(G116), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G122), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G107), .ZN(new_n278));
  INV_X1    g092(.A(G107), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n274), .A2(new_n276), .A3(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n272), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT13), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n268), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n270), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n268), .A2(new_n282), .ZN(new_n285));
  OAI21_X1  g099(.A(G134), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n275), .A2(KEYINPUT14), .A3(G122), .ZN(new_n288));
  OAI211_X1 g102(.A(G107), .B(new_n288), .C1(new_n277), .C2(KEYINPUT14), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n271), .B1(new_n268), .B2(new_n270), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n289), .B(new_n280), .C1(new_n272), .C2(new_n290), .ZN(new_n291));
  XOR2_X1   g105(.A(KEYINPUT75), .B(G217), .Z(new_n292));
  XOR2_X1   g106(.A(KEYINPUT9), .B(G234), .Z(new_n293));
  INV_X1    g107(.A(G953), .ZN(new_n294));
  AND3_X1   g108(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n287), .A2(new_n291), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n295), .B1(new_n287), .B2(new_n291), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n298), .A2(G902), .ZN(new_n299));
  INV_X1    g113(.A(G478), .ZN(new_n300));
  OR2_X1    g114(.A1(new_n300), .A2(KEYINPUT15), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n299), .A2(new_n301), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n266), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT87), .ZN(new_n307));
  INV_X1    g121(.A(G104), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G107), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT86), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT86), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(new_n308), .A3(G107), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n279), .A2(G104), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G101), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT3), .B1(new_n308), .B2(G107), .ZN(new_n316));
  AOI21_X1  g130(.A(G101), .B1(new_n308), .B2(G107), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT3), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(new_n279), .A3(G104), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n315), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT1), .B1(new_n267), .B2(G146), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n267), .A2(G146), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n194), .A2(G143), .ZN(new_n324));
  OAI211_X1 g138(.A(G128), .B(new_n322), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n194), .A2(G143), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n267), .A2(G146), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n326), .B(new_n327), .C1(KEYINPUT1), .C2(new_n269), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n325), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g143(.A(KEYINPUT10), .B1(new_n321), .B2(new_n329), .ZN(new_n330));
  AND2_X1   g144(.A1(new_n316), .A2(new_n319), .ZN(new_n331));
  AOI22_X1  g145(.A1(G101), .A2(new_n314), .B1(new_n331), .B2(new_n317), .ZN(new_n332));
  INV_X1    g146(.A(new_n329), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT10), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n316), .A2(new_n319), .A3(new_n309), .ZN(new_n337));
  INV_X1    g151(.A(G101), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n338), .A2(KEYINPUT4), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT84), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT84), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n337), .A2(new_n342), .A3(new_n339), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(KEYINPUT0), .A2(G128), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n326), .A2(new_n327), .A3(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(G143), .B(G146), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT0), .B(G128), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT67), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT67), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n346), .B(new_n351), .C1(new_n347), .C2(new_n348), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  AND2_X1   g167(.A1(new_n320), .A2(KEYINPUT4), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n337), .A2(G101), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n344), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n357), .A2(KEYINPUT85), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT85), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n350), .A2(new_n352), .B1(new_n354), .B2(new_n355), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n359), .B1(new_n360), .B2(new_n344), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n336), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT11), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n271), .B2(G137), .ZN(new_n364));
  INV_X1    g178(.A(G137), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(KEYINPUT11), .A3(G134), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n271), .A2(G137), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n364), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G131), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n232), .A2(new_n364), .A3(new_n366), .A4(new_n367), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n362), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n294), .A2(G227), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(KEYINPUT83), .ZN(new_n374));
  XNOR2_X1  g188(.A(G110), .B(G140), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n374), .B(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n357), .A2(KEYINPUT85), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n360), .A2(new_n359), .A3(new_n344), .ZN(new_n378));
  AOI22_X1  g192(.A1(new_n377), .A2(new_n378), .B1(new_n330), .B2(new_n335), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n364), .A2(new_n366), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n365), .A2(G134), .ZN(new_n381));
  NOR3_X1   g195(.A1(new_n381), .A2(new_n228), .A3(new_n227), .ZN(new_n382));
  AOI22_X1  g196(.A1(new_n380), .A2(new_n382), .B1(new_n368), .B2(G131), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n376), .B1(new_n379), .B2(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n383), .B(new_n336), .C1(new_n358), .C2(new_n361), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n321), .A2(new_n329), .ZN(new_n386));
  AOI22_X1  g200(.A1(new_n315), .A2(new_n320), .B1(new_n328), .B2(new_n325), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n371), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT12), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI211_X1 g204(.A(KEYINPUT12), .B(new_n371), .C1(new_n386), .C2(new_n387), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n385), .A2(new_n392), .ZN(new_n393));
  AOI22_X1  g207(.A1(new_n372), .A2(new_n384), .B1(new_n393), .B2(new_n376), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n307), .B(G469), .C1(new_n394), .C2(G902), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n384), .A2(new_n372), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n393), .A2(new_n376), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(G469), .ZN(new_n398));
  NAND2_X1  g212(.A1(G469), .A2(G902), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(KEYINPUT87), .A3(new_n399), .ZN(new_n400));
  XOR2_X1   g214(.A(KEYINPUT88), .B(G469), .Z(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n376), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n403), .B1(new_n372), .B2(new_n385), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n385), .A2(new_n403), .A3(new_n392), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n187), .B(new_n402), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n395), .A2(new_n400), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G221), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n408), .B1(new_n293), .B2(new_n187), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G952), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n411), .A2(G953), .ZN(new_n412));
  INV_X1    g226(.A(G234), .ZN(new_n413));
  INV_X1    g227(.A(G237), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  OAI211_X1 g229(.A(G902), .B(G953), .C1(new_n413), .C2(new_n414), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(KEYINPUT96), .ZN(new_n417));
  XOR2_X1   g231(.A(KEYINPUT21), .B(G898), .Z(new_n418));
  OAI21_X1  g232(.A(new_n415), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(G214), .B1(G237), .B2(G902), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G113), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT2), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT2), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G113), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G116), .B(G119), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G119), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G116), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n275), .A2(G119), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT2), .B(G113), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT66), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(KEYINPUT66), .B1(new_n426), .B2(new_n427), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n429), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n344), .A2(new_n438), .A3(new_n356), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT5), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(new_n430), .A3(G116), .ZN(new_n441));
  OAI211_X1 g255(.A(G113), .B(new_n441), .C1(new_n433), .C2(new_n440), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(new_n436), .B2(new_n437), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT89), .B1(new_n443), .B2(new_n321), .ZN(new_n444));
  XNOR2_X1  g258(.A(G110), .B(G122), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT89), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n435), .B1(new_n433), .B2(new_n434), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n426), .A2(new_n427), .A3(KEYINPUT66), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n332), .A2(new_n446), .A3(new_n449), .A4(new_n442), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n439), .A2(new_n444), .A3(new_n445), .A4(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G125), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n329), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n349), .A2(G125), .ZN(new_n454));
  INV_X1    g268(.A(G224), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT7), .B1(new_n455), .B2(G953), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n453), .A2(KEYINPUT91), .A3(new_n454), .A4(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n445), .B(KEYINPUT8), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n332), .B1(new_n449), .B2(new_n442), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n443), .A2(new_n321), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n451), .A2(new_n458), .A3(new_n462), .ZN(new_n463));
  OR2_X1    g277(.A1(new_n453), .A2(KEYINPUT90), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n453), .A2(KEYINPUT90), .B1(G125), .B2(new_n349), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n457), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT91), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n453), .A2(new_n454), .ZN(new_n468));
  OAI22_X1  g282(.A1(new_n466), .A2(new_n467), .B1(new_n468), .B2(new_n456), .ZN(new_n469));
  AOI21_X1  g283(.A(G902), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n439), .A2(new_n444), .A3(new_n450), .ZN(new_n471));
  INV_X1    g285(.A(new_n445), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n473), .A2(KEYINPUT6), .A3(new_n451), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n455), .A2(G953), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n468), .B(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n471), .A2(new_n477), .A3(new_n472), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n470), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(G210), .B1(G237), .B2(G902), .ZN(new_n481));
  XOR2_X1   g295(.A(new_n481), .B(KEYINPUT92), .Z(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n470), .A2(new_n479), .A3(new_n481), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n421), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND4_X1   g299(.A1(new_n306), .A2(new_n407), .A3(new_n410), .A4(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT32), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n271), .A2(G137), .ZN(new_n488));
  OAI21_X1  g302(.A(G131), .B1(new_n488), .B2(new_n381), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n364), .A2(new_n366), .ZN(new_n490));
  OR2_X1    g304(.A1(KEYINPUT64), .A2(G131), .ZN(new_n491));
  NAND2_X1  g305(.A1(KEYINPUT64), .A2(G131), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n491), .A2(new_n367), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n489), .B1(new_n490), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT68), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n370), .A2(KEYINPUT68), .A3(new_n489), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n333), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT69), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n438), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n352), .ZN(new_n501));
  NAND2_X1  g315(.A1(KEYINPUT0), .A2(G128), .ZN(new_n502));
  OR2_X1    g316(.A1(KEYINPUT0), .A2(G128), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n502), .B(new_n503), .C1(new_n323), .C2(new_n324), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n351), .B1(new_n504), .B2(new_n346), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n371), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n449), .A2(KEYINPUT69), .A3(new_n429), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n498), .A2(new_n500), .A3(new_n506), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT70), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n329), .B1(new_n495), .B2(new_n494), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n497), .A2(new_n510), .B1(new_n353), .B2(new_n371), .ZN(new_n511));
  AOI211_X1 g325(.A(new_n499), .B(new_n428), .C1(new_n447), .C2(new_n448), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT69), .B1(new_n449), .B2(new_n429), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT70), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n511), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n509), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT30), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n370), .A2(new_n489), .A3(new_n328), .A4(new_n325), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT65), .ZN(new_n520));
  OAI22_X1  g334(.A1(new_n519), .A2(new_n520), .B1(new_n383), .B2(new_n349), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n365), .A2(G134), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n367), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n380), .A2(new_n382), .B1(G131), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT65), .B1(new_n333), .B2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n518), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n498), .A2(new_n506), .A3(KEYINPUT30), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(new_n438), .A3(new_n527), .ZN(new_n528));
  XOR2_X1   g342(.A(KEYINPUT26), .B(G101), .Z(new_n529));
  NAND2_X1  g343(.A1(new_n188), .A2(G210), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n531), .B(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n517), .A2(KEYINPUT72), .A3(new_n528), .A4(new_n534), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n528), .A2(new_n509), .A3(new_n516), .A4(new_n534), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT72), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n535), .A2(KEYINPUT31), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n438), .B1(new_n521), .B2(new_n525), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n509), .A2(new_n516), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(KEYINPUT28), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT73), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT28), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n508), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n543), .B1(new_n508), .B2(new_n544), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n533), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n536), .A2(KEYINPUT31), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n539), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(G472), .A2(G902), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n487), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n553), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n550), .B1(new_n548), .B2(new_n533), .ZN(new_n556));
  AOI211_X1 g370(.A(KEYINPUT32), .B(new_n555), .C1(new_n556), .C2(new_n539), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n542), .A2(new_n534), .A3(new_n547), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n528), .A2(new_n509), .A3(new_n516), .ZN(new_n559));
  AOI21_X1  g373(.A(KEYINPUT29), .B1(new_n559), .B2(new_n533), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n558), .A2(KEYINPUT74), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT74), .B1(new_n558), .B2(new_n560), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n498), .A2(new_n506), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n563), .B1(new_n513), .B2(new_n512), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n509), .A2(new_n516), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT28), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n547), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n534), .A2(KEYINPUT29), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n187), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NOR3_X1   g383(.A1(new_n561), .A2(new_n562), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G472), .ZN(new_n571));
  OAI22_X1  g385(.A1(new_n554), .A2(new_n557), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT22), .B(G137), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n294), .A2(G221), .A3(G234), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n430), .A2(G128), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n269), .A2(G119), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT24), .B(G110), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT76), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT76), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(new_n579), .B2(new_n580), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT77), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n586), .B1(new_n430), .B2(G128), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(KEYINPUT23), .A3(new_n577), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT23), .B1(new_n269), .B2(G119), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n589), .A2(new_n586), .A3(new_n578), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(G110), .B1(new_n591), .B2(KEYINPUT78), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT78), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(new_n588), .B2(new_n590), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n585), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n595), .B1(new_n241), .B2(new_n242), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n579), .A2(new_n580), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n597), .B1(new_n591), .B2(G110), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(new_n222), .A3(new_n195), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n576), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n595), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n226), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n603), .A2(new_n575), .A3(new_n599), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n601), .A2(new_n604), .A3(new_n187), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT25), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n601), .A2(new_n604), .A3(KEYINPUT25), .A4(new_n187), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n292), .B1(new_n413), .B2(G902), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n601), .A2(new_n604), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n611), .A2(G902), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n486), .A2(new_n572), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  NAND2_X1  g433(.A1(new_n552), .A2(new_n553), .ZN(new_n620));
  AOI21_X1  g434(.A(G902), .B1(new_n556), .B2(new_n539), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n620), .B1(new_n571), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n407), .A2(new_n410), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n622), .A2(new_n623), .A3(new_n616), .ZN(new_n624));
  INV_X1    g438(.A(new_n420), .ZN(new_n625));
  INV_X1    g439(.A(new_n481), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n480), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n625), .B1(new_n627), .B2(new_n484), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n419), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n298), .B(KEYINPUT33), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(G478), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n299), .A2(new_n300), .ZN(new_n632));
  NAND2_X1  g446(.A1(G478), .A2(G902), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n266), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n629), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n624), .A2(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT34), .B(G104), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  INV_X1    g454(.A(new_n305), .ZN(new_n641));
  NOR3_X1   g455(.A1(new_n629), .A2(new_n641), .A3(new_n266), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n624), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G107), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT97), .B(KEYINPUT35), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  AOI21_X1  g460(.A(new_n610), .B1(new_n607), .B2(new_n608), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n603), .A2(new_n599), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT36), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n575), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(KEYINPUT98), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n648), .B(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n614), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n647), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n622), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n486), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT37), .B(G110), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  INV_X1    g473(.A(new_n266), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n417), .A2(G900), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n662), .A2(KEYINPUT99), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n415), .B1(new_n662), .B2(KEYINPUT99), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n660), .A2(new_n305), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n620), .A2(KEYINPUT32), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n552), .A2(new_n487), .A3(new_n553), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  OR2_X1    g484(.A1(new_n562), .A2(new_n569), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n671), .B2(new_n561), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n667), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n655), .ZN(new_n674));
  AND4_X1   g488(.A1(new_n410), .A2(new_n407), .A3(new_n628), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G128), .ZN(G30));
  NAND2_X1  g491(.A1(new_n483), .A2(new_n484), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n678), .B(KEYINPUT38), .Z(new_n679));
  NAND2_X1  g493(.A1(new_n266), .A2(new_n305), .ZN(new_n680));
  NOR4_X1   g494(.A1(new_n679), .A2(new_n625), .A3(new_n674), .A4(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n623), .ZN(new_n682));
  XOR2_X1   g496(.A(new_n665), .B(KEYINPUT39), .Z(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT40), .ZN(new_n685));
  INV_X1    g499(.A(new_n683), .ZN(new_n686));
  OR3_X1    g500(.A1(new_n623), .A2(KEYINPUT40), .A3(new_n686), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n535), .A2(new_n538), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n565), .A2(new_n533), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(G472), .B1(new_n690), .B2(G902), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n691), .B1(new_n554), .B2(new_n557), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n681), .A2(new_n685), .A3(new_n687), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT100), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G143), .ZN(G45));
  NAND3_X1  g509(.A1(new_n266), .A2(new_n635), .A3(new_n666), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n675), .A2(new_n572), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  INV_X1    g513(.A(new_n385), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n377), .A2(new_n378), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n383), .B1(new_n701), .B2(new_n336), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n376), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n385), .A2(new_n392), .A3(new_n403), .ZN(new_n704));
  AOI21_X1  g518(.A(G902), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(G469), .ZN(new_n706));
  OAI211_X1 g520(.A(new_n406), .B(new_n410), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT101), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n404), .A2(new_n405), .ZN(new_n710));
  OAI21_X1  g524(.A(G469), .B1(new_n710), .B2(G902), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n711), .A2(KEYINPUT101), .A3(new_n410), .A4(new_n406), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n713), .A2(new_n572), .A3(new_n617), .A4(new_n637), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  NAND4_X1  g530(.A1(new_n713), .A2(new_n642), .A3(new_n572), .A4(new_n617), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G116), .ZN(G18));
  INV_X1    g532(.A(new_n707), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(KEYINPUT102), .A3(new_n628), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT102), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n470), .A2(new_n479), .A3(new_n481), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n481), .B1(new_n470), .B2(new_n479), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n420), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n721), .B1(new_n707), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n674), .A2(new_n306), .A3(new_n419), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n572), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G119), .ZN(G21));
  AND3_X1   g543(.A1(new_n612), .A2(KEYINPUT103), .A3(new_n615), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT103), .B1(new_n612), .B2(new_n615), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n550), .B1(new_n567), .B2(new_n533), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n733), .A2(new_n539), .ZN(new_n734));
  OAI22_X1  g548(.A1(new_n734), .A2(new_n555), .B1(new_n621), .B2(new_n571), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n709), .A2(new_n419), .A3(new_n712), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT104), .B1(new_n680), .B2(new_n724), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT104), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n628), .A2(new_n739), .A3(new_n305), .A4(new_n266), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n736), .A2(new_n737), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G122), .ZN(G24));
  AOI21_X1  g557(.A(new_n696), .B1(new_n720), .B2(new_n725), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n555), .B1(new_n733), .B2(new_n539), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n552), .A2(new_n187), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n745), .B1(new_n746), .B2(G472), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT105), .B1(new_n747), .B2(new_n674), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n571), .B1(new_n552), .B2(new_n187), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT105), .ZN(new_n750));
  NOR4_X1   g564(.A1(new_n749), .A2(new_n750), .A3(new_n745), .A4(new_n655), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n744), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G125), .ZN(G27));
  OR2_X1    g567(.A1(new_n730), .A2(new_n731), .ZN(new_n754));
  AOI211_X1 g568(.A(G902), .B(new_n401), .C1(new_n703), .C2(new_n704), .ZN(new_n755));
  XOR2_X1   g569(.A(new_n399), .B(KEYINPUT106), .Z(new_n756));
  NAND2_X1  g570(.A1(new_n398), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n410), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n483), .A2(new_n484), .A3(new_n420), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n758), .A2(new_n696), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n572), .A2(new_n754), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(KEYINPUT42), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n572), .A2(new_n760), .A3(new_n763), .A4(new_n617), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g579(.A(KEYINPUT107), .B(G131), .Z(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(G33));
  NOR3_X1   g581(.A1(new_n667), .A2(new_n758), .A3(new_n759), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n572), .A2(new_n617), .A3(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  NAND2_X1  g584(.A1(new_n660), .A2(new_n635), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n771), .A2(KEYINPUT43), .ZN(new_n772));
  OR3_X1    g586(.A1(new_n266), .A2(KEYINPUT43), .A3(new_n634), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(KEYINPUT44), .A3(new_n622), .A4(new_n674), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n396), .A2(new_n397), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT45), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n394), .A2(KEYINPUT45), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n781), .A3(G469), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n756), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT46), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n782), .A2(KEYINPUT46), .A3(new_n756), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n786), .A2(KEYINPUT108), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(KEYINPUT108), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n406), .B(new_n785), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n410), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n790), .A2(new_n686), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n774), .A2(new_n622), .A3(new_n674), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT44), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n759), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n777), .A2(new_n791), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G137), .ZN(G39));
  NOR4_X1   g610(.A1(new_n572), .A2(new_n617), .A3(new_n696), .A4(new_n759), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n789), .A2(KEYINPUT47), .A3(new_n410), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT47), .B1(new_n789), .B2(new_n410), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n797), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(G140), .ZN(G42));
  NOR4_X1   g616(.A1(new_n732), .A2(new_n771), .A3(new_n409), .A4(new_n625), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT110), .ZN(new_n804));
  INV_X1    g618(.A(new_n692), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n711), .A2(new_n406), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n806), .B(KEYINPUT49), .Z(new_n807));
  NAND4_X1  g621(.A1(new_n804), .A2(new_n805), .A3(new_n679), .A4(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n398), .A2(new_n756), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n409), .B1(new_n810), .B2(new_n406), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n647), .A2(new_n654), .A3(new_n665), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT113), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n406), .A2(new_n398), .A3(new_n756), .ZN(new_n814));
  AND4_X1   g628(.A1(KEYINPUT113), .A2(new_n812), .A3(new_n814), .A4(new_n410), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n692), .B(new_n741), .C1(new_n813), .C2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n752), .A2(new_n676), .A3(new_n698), .A4(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n750), .B1(new_n735), .B2(new_n655), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n747), .A2(KEYINPUT105), .A3(new_n674), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n822), .A2(new_n744), .B1(new_n673), .B2(new_n675), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n816), .A2(new_n698), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT52), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n819), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n760), .B1(new_n748), .B2(new_n751), .ZN(new_n827));
  INV_X1    g641(.A(new_n759), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n305), .B(KEYINPUT112), .ZN(new_n829));
  NOR4_X1   g643(.A1(new_n829), .A2(new_n655), .A3(new_n266), .A4(new_n665), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n572), .A2(new_n682), .A3(new_n828), .A4(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n827), .A2(new_n769), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n765), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n622), .A2(new_n616), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n407), .A2(new_n410), .A3(new_n485), .ZN(new_n835));
  INV_X1    g649(.A(new_n636), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n618), .A3(KEYINPUT111), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT111), .B1(new_n837), .B2(new_n618), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n834), .A2(new_n835), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n829), .A2(new_n660), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n657), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n742), .A2(new_n728), .A3(new_n717), .A4(new_n714), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n833), .A2(new_n838), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n809), .B1(new_n826), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n843), .A2(new_n838), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n817), .A2(new_n818), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n823), .A2(new_n824), .A3(KEYINPUT52), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n844), .A2(new_n832), .A3(new_n765), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n849), .A2(new_n852), .A3(KEYINPUT53), .A4(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n847), .A2(new_n848), .A3(new_n854), .ZN(new_n855));
  OAI211_X1 g669(.A(KEYINPUT114), .B(new_n809), .C1(new_n826), .C2(new_n846), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n855), .A2(KEYINPUT54), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n847), .A2(new_n858), .A3(new_n854), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n857), .A2(KEYINPUT115), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT115), .B1(new_n857), .B2(new_n859), .ZN(new_n861));
  INV_X1    g675(.A(new_n415), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n772), .A2(new_n862), .A3(new_n773), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n736), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  AOI211_X1 g679(.A(new_n411), .B(G953), .C1(new_n865), .C2(new_n726), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n719), .A2(new_n617), .A3(new_n862), .A4(new_n828), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n692), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n868), .A2(new_n836), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n863), .A2(new_n719), .A3(new_n828), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT48), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n732), .B1(new_n670), .B2(new_n672), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n872), .B1(new_n871), .B2(new_n873), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n864), .A2(new_n759), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n799), .A2(new_n800), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n711), .A2(new_n409), .A3(new_n406), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n707), .A2(new_n420), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n863), .A2(new_n679), .A3(new_n736), .A4(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT50), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n882), .B(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n266), .A2(new_n635), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n871), .A2(new_n822), .B1(new_n868), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n884), .A2(KEYINPUT51), .A3(new_n886), .ZN(new_n887));
  OAI221_X1 g701(.A(new_n870), .B1(new_n874), .B2(new_n875), .C1(new_n880), .C2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT47), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n785), .A2(new_n406), .ZN(new_n890));
  INV_X1    g704(.A(new_n788), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n786), .A2(KEYINPUT108), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n889), .B1(new_n893), .B2(new_n409), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n894), .A2(KEYINPUT116), .A3(new_n798), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n879), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT116), .B1(new_n894), .B2(new_n798), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n876), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n884), .A2(new_n886), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT51), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT117), .B1(new_n888), .B2(new_n901), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n866), .B(new_n869), .C1(new_n874), .C2(new_n875), .ZN(new_n903));
  INV_X1    g717(.A(new_n880), .ZN(new_n904));
  INV_X1    g718(.A(new_n887), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT117), .ZN(new_n907));
  INV_X1    g721(.A(new_n897), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n895), .A3(new_n879), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n899), .B1(new_n909), .B2(new_n876), .ZN(new_n910));
  OAI211_X1 g724(.A(new_n906), .B(new_n907), .C1(new_n910), .C2(KEYINPUT51), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n902), .A2(new_n911), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n860), .A2(new_n861), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(G952), .A2(G953), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n808), .B1(new_n913), .B2(new_n914), .ZN(G75));
  NAND2_X1  g729(.A1(new_n474), .A2(new_n478), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(new_n476), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT55), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n187), .B1(new_n847), .B2(new_n854), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(G210), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT56), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n918), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n294), .A2(G952), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n918), .A2(new_n921), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n919), .B2(new_n482), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(G51));
  AOI211_X1 g740(.A(new_n187), .B(new_n782), .C1(new_n847), .C2(new_n854), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n847), .A2(new_n854), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT54), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n859), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n756), .B(KEYINPUT57), .Z(new_n931));
  AOI21_X1  g745(.A(new_n710), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT118), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n927), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n931), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n929), .B2(new_n859), .ZN(new_n936));
  OAI21_X1  g750(.A(KEYINPUT118), .B1(new_n936), .B2(new_n710), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n923), .B1(new_n934), .B2(new_n937), .ZN(G54));
  NAND3_X1  g752(.A1(new_n919), .A2(KEYINPUT58), .A3(G475), .ZN(new_n939));
  INV_X1    g753(.A(new_n262), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n941), .A2(new_n942), .A3(new_n923), .ZN(G60));
  INV_X1    g757(.A(new_n923), .ZN(new_n944));
  INV_X1    g758(.A(new_n930), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n630), .B(KEYINPUT119), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n633), .B(KEYINPUT59), .Z(new_n947));
  OR2_X1    g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n944), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n947), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n860), .B2(new_n861), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n949), .B1(new_n951), .B2(new_n946), .ZN(G63));
  NAND2_X1  g766(.A1(G217), .A2(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT60), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(new_n847), .B2(new_n854), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n652), .B(KEYINPUT121), .Z(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n957), .B(new_n944), .C1(new_n613), .C2(new_n955), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n958), .A2(KEYINPUT120), .A3(KEYINPUT61), .ZN(new_n959));
  AOI21_X1  g773(.A(KEYINPUT61), .B1(new_n958), .B2(KEYINPUT120), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(G66));
  AOI21_X1  g775(.A(new_n294), .B1(new_n418), .B2(G224), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n849), .A2(new_n845), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(new_n963), .B2(new_n294), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n916), .B1(G898), .B2(new_n294), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT122), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n964), .B(new_n966), .ZN(G69));
  NAND2_X1  g781(.A1(new_n526), .A2(new_n527), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n253), .A2(new_n254), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n795), .A2(new_n801), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT100), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n693), .B(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n823), .A2(new_n698), .ZN(new_n975));
  OAI21_X1  g789(.A(KEYINPUT62), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT62), .ZN(new_n977));
  INV_X1    g791(.A(new_n975), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n694), .A2(new_n977), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n841), .A2(new_n636), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT123), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n759), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n982), .B1(new_n981), .B2(new_n980), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n572), .A2(new_n617), .ZN(new_n984));
  NOR3_X1   g798(.A1(new_n983), .A2(new_n984), .A3(new_n684), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT124), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n972), .A2(new_n976), .A3(new_n979), .A4(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n970), .B1(new_n987), .B2(new_n294), .ZN(new_n988));
  NAND2_X1  g802(.A1(G900), .A2(G953), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n970), .A2(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n791), .A2(new_n741), .A3(new_n873), .ZN(new_n991));
  AND3_X1   g805(.A1(new_n762), .A2(new_n764), .A3(new_n769), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n991), .A2(new_n978), .A3(new_n992), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n971), .A2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n990), .B1(new_n994), .B2(new_n294), .ZN(new_n995));
  OAI21_X1  g809(.A(KEYINPUT125), .B1(new_n988), .B2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n995), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT125), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n977), .B1(new_n694), .B2(new_n978), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n986), .A2(new_n795), .A3(new_n801), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(G953), .B1(new_n1001), .B2(new_n979), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n997), .B(new_n998), .C1(new_n1002), .C2(new_n970), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n294), .B1(G227), .B2(G900), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n996), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1004), .ZN(new_n1006));
  OAI211_X1 g820(.A(KEYINPUT125), .B(new_n1006), .C1(new_n988), .C2(new_n995), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n1005), .A2(new_n1007), .ZN(G72));
  XNOR2_X1  g822(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n571), .A2(new_n187), .ZN(new_n1010));
  XOR2_X1   g824(.A(new_n1009), .B(new_n1010), .Z(new_n1011));
  NAND2_X1  g825(.A1(new_n559), .A2(new_n533), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1011), .B1(new_n688), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n855), .A2(new_n856), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1011), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1015), .B1(new_n987), .B2(new_n963), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n533), .B1(new_n517), .B2(new_n528), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT127), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(new_n994), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1015), .B1(new_n1021), .B2(new_n963), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n559), .A2(new_n534), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n923), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1016), .A2(KEYINPUT127), .A3(new_n1017), .ZN(new_n1025));
  AND4_X1   g839(.A1(new_n1014), .A2(new_n1020), .A3(new_n1024), .A4(new_n1025), .ZN(G57));
endmodule


