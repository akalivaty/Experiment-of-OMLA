

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589;

  INV_X1 U325 ( .A(KEYINPUT47), .ZN(n422) );
  XNOR2_X1 U326 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U327 ( .A(n418), .B(n417), .ZN(n581) );
  XNOR2_X1 U328 ( .A(n459), .B(KEYINPUT41), .ZN(n545) );
  INV_X1 U329 ( .A(G218GAT), .ZN(n456) );
  XNOR2_X1 U330 ( .A(n456), .B(KEYINPUT62), .ZN(n457) );
  XNOR2_X1 U331 ( .A(n458), .B(n457), .ZN(G1355GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT8), .B(KEYINPUT72), .Z(n294) );
  XNOR2_X1 U333 ( .A(G36GAT), .B(G29GAT), .ZN(n293) );
  XNOR2_X1 U334 ( .A(n294), .B(n293), .ZN(n295) );
  XNOR2_X1 U335 ( .A(KEYINPUT7), .B(n295), .ZN(n402) );
  INV_X1 U336 ( .A(n402), .ZN(n302) );
  XOR2_X1 U337 ( .A(G43GAT), .B(G134GAT), .Z(n335) );
  XOR2_X1 U338 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n297) );
  XNOR2_X1 U339 ( .A(G218GAT), .B(KEYINPUT64), .ZN(n296) );
  XNOR2_X1 U340 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U341 ( .A(n335), .B(n298), .Z(n300) );
  NAND2_X1 U342 ( .A1(G232GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U343 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U344 ( .A(n302), .B(n301), .ZN(n315) );
  XOR2_X1 U345 ( .A(KEYINPUT10), .B(KEYINPUT67), .Z(n304) );
  XNOR2_X1 U346 ( .A(G99GAT), .B(KEYINPUT82), .ZN(n303) );
  XNOR2_X1 U347 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U348 ( .A(KEYINPUT65), .B(KEYINPUT66), .Z(n306) );
  XNOR2_X1 U349 ( .A(G190GAT), .B(G106GAT), .ZN(n305) );
  XNOR2_X1 U350 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U351 ( .A(n308), .B(n307), .Z(n313) );
  XNOR2_X1 U352 ( .A(G50GAT), .B(KEYINPUT81), .ZN(n309) );
  XNOR2_X1 U353 ( .A(n309), .B(G162GAT), .ZN(n321) );
  XOR2_X1 U354 ( .A(G85GAT), .B(G92GAT), .Z(n310) );
  XNOR2_X1 U355 ( .A(KEYINPUT76), .B(n310), .ZN(n412) );
  INV_X1 U356 ( .A(n412), .ZN(n311) );
  XNOR2_X1 U357 ( .A(n321), .B(n311), .ZN(n312) );
  XNOR2_X1 U358 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U359 ( .A(n315), .B(n314), .ZN(n573) );
  XNOR2_X1 U360 ( .A(KEYINPUT36), .B(n573), .ZN(n486) );
  XOR2_X1 U361 ( .A(G211GAT), .B(KEYINPUT21), .Z(n317) );
  XNOR2_X1 U362 ( .A(G197GAT), .B(G218GAT), .ZN(n316) );
  XNOR2_X1 U363 ( .A(n317), .B(n316), .ZN(n357) );
  XOR2_X1 U364 ( .A(G22GAT), .B(G155GAT), .Z(n367) );
  XOR2_X1 U365 ( .A(n357), .B(n367), .Z(n319) );
  NAND2_X1 U366 ( .A1(G228GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U368 ( .A(n320), .B(G204GAT), .Z(n323) );
  XNOR2_X1 U369 ( .A(n321), .B(KEYINPUT22), .ZN(n322) );
  XNOR2_X1 U370 ( .A(n323), .B(n322), .ZN(n327) );
  XOR2_X1 U371 ( .A(KEYINPUT95), .B(KEYINPUT23), .Z(n325) );
  XNOR2_X1 U372 ( .A(KEYINPUT94), .B(KEYINPUT24), .ZN(n324) );
  XNOR2_X1 U373 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U374 ( .A(n327), .B(n326), .Z(n332) );
  XOR2_X1 U375 ( .A(G78GAT), .B(G148GAT), .Z(n329) );
  XNOR2_X1 U376 ( .A(G106GAT), .B(KEYINPUT75), .ZN(n328) );
  XNOR2_X1 U377 ( .A(n329), .B(n328), .ZN(n405) );
  XNOR2_X1 U378 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n330) );
  XNOR2_X1 U379 ( .A(n330), .B(KEYINPUT3), .ZN(n448) );
  XNOR2_X1 U380 ( .A(n405), .B(n448), .ZN(n331) );
  XNOR2_X1 U381 ( .A(n332), .B(n331), .ZN(n558) );
  XOR2_X1 U382 ( .A(KEYINPUT89), .B(KEYINPUT92), .Z(n334) );
  XNOR2_X1 U383 ( .A(G176GAT), .B(KEYINPUT91), .ZN(n333) );
  XNOR2_X1 U384 ( .A(n334), .B(n333), .ZN(n339) );
  XOR2_X1 U385 ( .A(KEYINPUT20), .B(KEYINPUT90), .Z(n337) );
  XOR2_X1 U386 ( .A(G15GAT), .B(G127GAT), .Z(n371) );
  XNOR2_X1 U387 ( .A(n335), .B(n371), .ZN(n336) );
  XNOR2_X1 U388 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U389 ( .A(n339), .B(n338), .Z(n341) );
  NAND2_X1 U390 ( .A1(G227GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U391 ( .A(n341), .B(n340), .ZN(n343) );
  XNOR2_X1 U392 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n342) );
  XNOR2_X1 U393 ( .A(n342), .B(KEYINPUT88), .ZN(n440) );
  XOR2_X1 U394 ( .A(n343), .B(n440), .Z(n350) );
  XNOR2_X1 U395 ( .A(G183GAT), .B(KEYINPUT17), .ZN(n344) );
  XNOR2_X1 U396 ( .A(n344), .B(KEYINPUT18), .ZN(n345) );
  XOR2_X1 U397 ( .A(n345), .B(KEYINPUT19), .Z(n347) );
  XNOR2_X1 U398 ( .A(G169GAT), .B(G190GAT), .ZN(n346) );
  XOR2_X1 U399 ( .A(n347), .B(n346), .Z(n363) );
  XNOR2_X1 U400 ( .A(G99GAT), .B(G71GAT), .ZN(n348) );
  XNOR2_X1 U401 ( .A(n348), .B(G120GAT), .ZN(n413) );
  XOR2_X1 U402 ( .A(n363), .B(n413), .Z(n349) );
  XNOR2_X1 U403 ( .A(n350), .B(n349), .ZN(n562) );
  INV_X1 U404 ( .A(n562), .ZN(n498) );
  NAND2_X1 U405 ( .A1(n558), .A2(n498), .ZN(n351) );
  XNOR2_X1 U406 ( .A(KEYINPUT26), .B(n351), .ZN(n540) );
  XOR2_X1 U407 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n353) );
  NAND2_X1 U408 ( .A1(G226GAT), .A2(G233GAT), .ZN(n352) );
  XNOR2_X1 U409 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U410 ( .A(n354), .B(KEYINPUT101), .Z(n359) );
  XOR2_X1 U411 ( .A(G64GAT), .B(KEYINPUT78), .Z(n356) );
  XNOR2_X1 U412 ( .A(G176GAT), .B(G204GAT), .ZN(n355) );
  XNOR2_X1 U413 ( .A(n356), .B(n355), .ZN(n404) );
  XNOR2_X1 U414 ( .A(n357), .B(n404), .ZN(n358) );
  XNOR2_X1 U415 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U416 ( .A(G8GAT), .B(KEYINPUT83), .Z(n372) );
  XOR2_X1 U417 ( .A(n360), .B(n372), .Z(n362) );
  XNOR2_X1 U418 ( .A(G36GAT), .B(G92GAT), .ZN(n361) );
  XNOR2_X1 U419 ( .A(n362), .B(n361), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n364), .B(n363), .ZN(n495) );
  XOR2_X1 U421 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n366) );
  XNOR2_X1 U422 ( .A(G1GAT), .B(G64GAT), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n384) );
  XOR2_X1 U424 ( .A(n367), .B(KEYINPUT12), .Z(n369) );
  NAND2_X1 U425 ( .A1(G231GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U426 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U427 ( .A(n371), .B(n370), .ZN(n382) );
  XOR2_X1 U428 ( .A(G57GAT), .B(KEYINPUT13), .Z(n414) );
  XOR2_X1 U429 ( .A(n414), .B(n372), .Z(n374) );
  XNOR2_X1 U430 ( .A(G78GAT), .B(G211GAT), .ZN(n373) );
  XNOR2_X1 U431 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U432 ( .A(KEYINPUT14), .B(KEYINPUT85), .Z(n376) );
  XNOR2_X1 U433 ( .A(KEYINPUT84), .B(KEYINPUT15), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U435 ( .A(n378), .B(n377), .Z(n380) );
  XNOR2_X1 U436 ( .A(G183GAT), .B(G71GAT), .ZN(n379) );
  XNOR2_X1 U437 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U438 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U439 ( .A(n384), .B(n383), .ZN(n569) );
  INV_X1 U440 ( .A(n569), .ZN(n586) );
  XOR2_X1 U441 ( .A(G22GAT), .B(G197GAT), .Z(n386) );
  XNOR2_X1 U442 ( .A(G169GAT), .B(G141GAT), .ZN(n385) );
  XNOR2_X1 U443 ( .A(n386), .B(n385), .ZN(n390) );
  XOR2_X1 U444 ( .A(G1GAT), .B(KEYINPUT74), .Z(n388) );
  XNOR2_X1 U445 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n387) );
  XNOR2_X1 U446 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U447 ( .A(n390), .B(n389), .Z(n401) );
  XOR2_X1 U448 ( .A(KEYINPUT73), .B(KEYINPUT30), .Z(n392) );
  XNOR2_X1 U449 ( .A(KEYINPUT71), .B(KEYINPUT70), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n392), .B(n391), .ZN(n399) );
  XOR2_X1 U451 ( .A(G15GAT), .B(G113GAT), .Z(n394) );
  XNOR2_X1 U452 ( .A(G50GAT), .B(G43GAT), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U454 ( .A(KEYINPUT69), .B(n395), .Z(n397) );
  NAND2_X1 U455 ( .A1(G229GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U457 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n401), .B(n400), .ZN(n403) );
  XOR2_X1 U459 ( .A(n403), .B(n402), .Z(n576) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n410) );
  XOR2_X1 U461 ( .A(KEYINPUT77), .B(KEYINPUT32), .Z(n407) );
  NAND2_X1 U462 ( .A1(G230GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U463 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U464 ( .A(n408), .B(KEYINPUT79), .Z(n409) );
  XNOR2_X1 U465 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U466 ( .A(n411), .B(KEYINPUT33), .Z(n418) );
  XNOR2_X1 U467 ( .A(n413), .B(n412), .ZN(n416) );
  XNOR2_X1 U468 ( .A(n414), .B(KEYINPUT31), .ZN(n415) );
  INV_X1 U469 ( .A(n581), .ZN(n459) );
  NAND2_X1 U470 ( .A1(n576), .A2(n545), .ZN(n419) );
  XNOR2_X1 U471 ( .A(KEYINPUT46), .B(n419), .ZN(n420) );
  NAND2_X1 U472 ( .A1(n420), .A2(n573), .ZN(n421) );
  NOR2_X1 U473 ( .A1(n586), .A2(n421), .ZN(n423) );
  XNOR2_X1 U474 ( .A(n423), .B(n422), .ZN(n429) );
  NOR2_X1 U475 ( .A1(n486), .A2(n569), .ZN(n424) );
  XOR2_X1 U476 ( .A(KEYINPUT45), .B(n424), .Z(n425) );
  NOR2_X1 U477 ( .A1(n581), .A2(n425), .ZN(n426) );
  XOR2_X1 U478 ( .A(KEYINPUT114), .B(n426), .Z(n427) );
  NOR2_X1 U479 ( .A1(n576), .A2(n427), .ZN(n428) );
  NOR2_X1 U480 ( .A1(n429), .A2(n428), .ZN(n430) );
  XNOR2_X1 U481 ( .A(KEYINPUT48), .B(n430), .ZN(n539) );
  NOR2_X1 U482 ( .A1(n495), .A2(n539), .ZN(n431) );
  XNOR2_X1 U483 ( .A(KEYINPUT54), .B(n431), .ZN(n453) );
  XOR2_X1 U484 ( .A(KEYINPUT98), .B(KEYINPUT97), .Z(n433) );
  XNOR2_X1 U485 ( .A(G1GAT), .B(G57GAT), .ZN(n432) );
  XNOR2_X1 U486 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U487 ( .A(G155GAT), .B(G148GAT), .Z(n435) );
  XNOR2_X1 U488 ( .A(G120GAT), .B(G127GAT), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U490 ( .A(n437), .B(n436), .ZN(n452) );
  XOR2_X1 U491 ( .A(G85GAT), .B(G162GAT), .Z(n439) );
  XNOR2_X1 U492 ( .A(G29GAT), .B(G134GAT), .ZN(n438) );
  XNOR2_X1 U493 ( .A(n439), .B(n438), .ZN(n444) );
  XOR2_X1 U494 ( .A(KEYINPUT4), .B(n440), .Z(n442) );
  NAND2_X1 U495 ( .A1(G225GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U496 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U497 ( .A(n444), .B(n443), .Z(n450) );
  XOR2_X1 U498 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n446) );
  XNOR2_X1 U499 ( .A(KEYINPUT6), .B(KEYINPUT96), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U502 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U503 ( .A(n452), .B(n451), .ZN(n491) );
  NAND2_X1 U504 ( .A1(n453), .A2(n491), .ZN(n557) );
  NOR2_X1 U505 ( .A1(n540), .A2(n557), .ZN(n454) );
  XOR2_X1 U506 ( .A(KEYINPUT123), .B(n454), .Z(n587) );
  INV_X1 U507 ( .A(n587), .ZN(n455) );
  NOR2_X1 U508 ( .A1(n486), .A2(n455), .ZN(n458) );
  INV_X1 U509 ( .A(n491), .ZN(n516) );
  NAND2_X1 U510 ( .A1(n576), .A2(n459), .ZN(n460) );
  XNOR2_X1 U511 ( .A(n460), .B(KEYINPUT80), .ZN(n488) );
  NAND2_X1 U512 ( .A1(n573), .A2(n586), .ZN(n461) );
  XOR2_X1 U513 ( .A(KEYINPUT16), .B(n461), .Z(n474) );
  XNOR2_X1 U514 ( .A(n495), .B(KEYINPUT27), .ZN(n467) );
  NOR2_X1 U515 ( .A1(n491), .A2(n467), .ZN(n542) );
  XOR2_X1 U516 ( .A(n558), .B(KEYINPUT68), .Z(n462) );
  XNOR2_X1 U517 ( .A(KEYINPUT28), .B(n462), .ZN(n502) );
  NAND2_X1 U518 ( .A1(n542), .A2(n502), .ZN(n528) );
  XNOR2_X1 U519 ( .A(KEYINPUT93), .B(n498), .ZN(n463) );
  NOR2_X1 U520 ( .A1(n528), .A2(n463), .ZN(n472) );
  NOR2_X1 U521 ( .A1(n495), .A2(n498), .ZN(n464) );
  NOR2_X1 U522 ( .A1(n558), .A2(n464), .ZN(n465) );
  XOR2_X1 U523 ( .A(n465), .B(KEYINPUT102), .Z(n466) );
  XNOR2_X1 U524 ( .A(KEYINPUT25), .B(n466), .ZN(n469) );
  NOR2_X1 U525 ( .A1(n540), .A2(n467), .ZN(n468) );
  NOR2_X1 U526 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U527 ( .A1(n516), .A2(n470), .ZN(n471) );
  NOR2_X1 U528 ( .A1(n472), .A2(n471), .ZN(n483) );
  INV_X1 U529 ( .A(n483), .ZN(n473) );
  NAND2_X1 U530 ( .A1(n474), .A2(n473), .ZN(n505) );
  NOR2_X1 U531 ( .A1(n488), .A2(n505), .ZN(n481) );
  NAND2_X1 U532 ( .A1(n516), .A2(n481), .ZN(n477) );
  XOR2_X1 U533 ( .A(G1GAT), .B(KEYINPUT34), .Z(n475) );
  XNOR2_X1 U534 ( .A(KEYINPUT103), .B(n475), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n477), .B(n476), .ZN(G1324GAT) );
  INV_X1 U536 ( .A(n495), .ZN(n519) );
  NAND2_X1 U537 ( .A1(n519), .A2(n481), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n478), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U539 ( .A(G15GAT), .B(KEYINPUT35), .Z(n480) );
  NAND2_X1 U540 ( .A1(n481), .A2(n562), .ZN(n479) );
  XNOR2_X1 U541 ( .A(n480), .B(n479), .ZN(G1326GAT) );
  INV_X1 U542 ( .A(n502), .ZN(n524) );
  NAND2_X1 U543 ( .A1(n481), .A2(n524), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n482), .B(G22GAT), .ZN(G1327GAT) );
  XNOR2_X1 U545 ( .A(KEYINPUT106), .B(KEYINPUT39), .ZN(n493) );
  NOR2_X1 U546 ( .A1(n586), .A2(n483), .ZN(n484) );
  XOR2_X1 U547 ( .A(KEYINPUT104), .B(n484), .Z(n485) );
  NOR2_X1 U548 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U549 ( .A(KEYINPUT37), .B(n487), .ZN(n513) );
  NOR2_X1 U550 ( .A1(n488), .A2(n513), .ZN(n490) );
  XNOR2_X1 U551 ( .A(KEYINPUT38), .B(KEYINPUT105), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n490), .B(n489), .ZN(n503) );
  NOR2_X1 U553 ( .A1(n491), .A2(n503), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G29GAT), .B(n494), .ZN(G1328GAT) );
  XNOR2_X1 U556 ( .A(G36GAT), .B(KEYINPUT107), .ZN(n497) );
  NOR2_X1 U557 ( .A1(n495), .A2(n503), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n497), .B(n496), .ZN(G1329GAT) );
  NOR2_X1 U559 ( .A1(n503), .A2(n498), .ZN(n500) );
  XNOR2_X1 U560 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U562 ( .A(G43GAT), .B(n501), .Z(G1330GAT) );
  NOR2_X1 U563 ( .A1(n503), .A2(n502), .ZN(n504) );
  XOR2_X1 U564 ( .A(G50GAT), .B(n504), .Z(G1331GAT) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n507) );
  XNOR2_X1 U566 ( .A(KEYINPUT109), .B(n545), .ZN(n565) );
  OR2_X1 U567 ( .A1(n576), .A2(n565), .ZN(n514) );
  NOR2_X1 U568 ( .A1(n514), .A2(n505), .ZN(n510) );
  NAND2_X1 U569 ( .A1(n510), .A2(n516), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n507), .B(n506), .ZN(G1332GAT) );
  NAND2_X1 U571 ( .A1(n519), .A2(n510), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n508), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U573 ( .A1(n510), .A2(n562), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n509), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U575 ( .A(G78GAT), .B(KEYINPUT43), .Z(n512) );
  NAND2_X1 U576 ( .A1(n510), .A2(n524), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  XOR2_X1 U578 ( .A(G85GAT), .B(KEYINPUT111), .Z(n518) );
  NOR2_X1 U579 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n515), .B(KEYINPUT110), .ZN(n525) );
  NAND2_X1 U581 ( .A1(n525), .A2(n516), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(G1336GAT) );
  NAND2_X1 U583 ( .A1(n525), .A2(n519), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n520), .B(KEYINPUT112), .ZN(n521) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(n521), .ZN(G1337GAT) );
  XOR2_X1 U586 ( .A(G99GAT), .B(KEYINPUT113), .Z(n523) );
  NAND2_X1 U587 ( .A1(n562), .A2(n525), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(G1338GAT) );
  NAND2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n526), .B(KEYINPUT44), .ZN(n527) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  INV_X1 U592 ( .A(n576), .ZN(n563) );
  NOR2_X1 U593 ( .A1(n539), .A2(n528), .ZN(n529) );
  NAND2_X1 U594 ( .A1(n562), .A2(n529), .ZN(n536) );
  NOR2_X1 U595 ( .A1(n563), .A2(n536), .ZN(n530) );
  XOR2_X1 U596 ( .A(G113GAT), .B(n530), .Z(G1340GAT) );
  NOR2_X1 U597 ( .A1(n565), .A2(n536), .ZN(n532) );
  XNOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  NOR2_X1 U600 ( .A1(n569), .A2(n536), .ZN(n534) );
  XNOR2_X1 U601 ( .A(KEYINPUT50), .B(KEYINPUT115), .ZN(n533) );
  XNOR2_X1 U602 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  NOR2_X1 U604 ( .A1(n573), .A2(n536), .ZN(n538) );
  XNOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n537) );
  XNOR2_X1 U606 ( .A(n538), .B(n537), .ZN(G1343GAT) );
  NOR2_X1 U607 ( .A1(n540), .A2(n539), .ZN(n541) );
  NAND2_X1 U608 ( .A1(n542), .A2(n541), .ZN(n553) );
  NOR2_X1 U609 ( .A1(n563), .A2(n553), .ZN(n543) );
  XOR2_X1 U610 ( .A(KEYINPUT116), .B(n543), .Z(n544) );
  XNOR2_X1 U611 ( .A(G141GAT), .B(n544), .ZN(G1344GAT) );
  XOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT117), .Z(n547) );
  INV_X1 U613 ( .A(n553), .ZN(n550) );
  NAND2_X1 U614 ( .A1(n550), .A2(n545), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(n549) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n548) );
  XNOR2_X1 U617 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  NAND2_X1 U618 ( .A1(n550), .A2(n586), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n551), .B(KEYINPUT118), .ZN(n552) );
  XNOR2_X1 U620 ( .A(G155GAT), .B(n552), .ZN(G1346GAT) );
  NOR2_X1 U621 ( .A1(n573), .A2(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n554) );
  XNOR2_X1 U623 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U624 ( .A(G162GAT), .B(n556), .ZN(G1347GAT) );
  NOR2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n560) );
  XNOR2_X1 U626 ( .A(KEYINPUT121), .B(KEYINPUT55), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n572) );
  NOR2_X1 U629 ( .A1(n563), .A2(n572), .ZN(n564) );
  XOR2_X1 U630 ( .A(G169GAT), .B(n564), .Z(G1348GAT) );
  NOR2_X1 U631 ( .A1(n565), .A2(n572), .ZN(n567) );
  XNOR2_X1 U632 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(G176GAT), .B(n568), .ZN(G1349GAT) );
  NOR2_X1 U635 ( .A1(n569), .A2(n572), .ZN(n570) );
  XOR2_X1 U636 ( .A(KEYINPUT122), .B(n570), .Z(n571) );
  XNOR2_X1 U637 ( .A(G183GAT), .B(n571), .ZN(G1350GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U639 ( .A(KEYINPUT58), .B(n574), .Z(n575) );
  XNOR2_X1 U640 ( .A(G190GAT), .B(n575), .ZN(G1351GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n587), .ZN(n580) );
  XOR2_X1 U642 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n583) );
  NAND2_X1 U647 ( .A1(n587), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n585) );
  XOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT125), .Z(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  XOR2_X1 U651 ( .A(G211GAT), .B(KEYINPUT127), .Z(n589) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n589), .B(n588), .ZN(G1354GAT) );
endmodule

