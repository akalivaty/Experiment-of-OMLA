

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U553 ( .A(n686), .B(KEYINPUT90), .ZN(n768) );
  NOR2_X1 U554 ( .A1(n751), .A2(n752), .ZN(n697) );
  BUF_X1 U555 ( .A(n695), .Z(n807) );
  NAND2_X1 U556 ( .A1(n882), .A2(G137), .ZN(n540) );
  XOR2_X1 U557 ( .A(n543), .B(KEYINPUT23), .Z(n520) );
  XOR2_X1 U558 ( .A(KEYINPUT30), .B(KEYINPUT100), .Z(n521) );
  XOR2_X1 U559 ( .A(n730), .B(KEYINPUT28), .Z(n522) );
  NOR2_X1 U560 ( .A1(n753), .A2(n752), .ZN(n523) );
  NOR2_X1 U561 ( .A1(n714), .A2(n713), .ZN(n719) );
  BUF_X1 U562 ( .A(n703), .Z(n704) );
  BUF_X1 U563 ( .A(n704), .Z(n737) );
  INV_X1 U564 ( .A(G168), .ZN(n700) );
  AND2_X1 U565 ( .A1(n701), .A2(n700), .ZN(n702) );
  INV_X1 U566 ( .A(n991), .ZN(n760) );
  NOR2_X1 U567 ( .A1(n761), .A2(n760), .ZN(n762) );
  AND2_X1 U568 ( .A1(n763), .A2(n762), .ZN(n764) );
  INV_X1 U569 ( .A(KEYINPUT17), .ZN(n537) );
  NOR2_X1 U570 ( .A1(G543), .A2(G651), .ZN(n641) );
  AND2_X2 U571 ( .A1(n542), .A2(G2104), .ZN(n883) );
  NOR2_X1 U572 ( .A1(n621), .A2(G651), .ZN(n640) );
  NAND2_X1 U573 ( .A1(n641), .A2(G89), .ZN(n524) );
  XNOR2_X1 U574 ( .A(n524), .B(KEYINPUT4), .ZN(n526) );
  XOR2_X1 U575 ( .A(KEYINPUT0), .B(G543), .Z(n621) );
  INV_X1 U576 ( .A(G651), .ZN(n528) );
  NOR2_X1 U577 ( .A1(n621), .A2(n528), .ZN(n634) );
  NAND2_X1 U578 ( .A1(G76), .A2(n634), .ZN(n525) );
  NAND2_X1 U579 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U580 ( .A(KEYINPUT5), .B(n527), .ZN(n535) );
  NOR2_X1 U581 ( .A1(G543), .A2(n528), .ZN(n529) );
  XOR2_X1 U582 ( .A(KEYINPUT1), .B(n529), .Z(n637) );
  NAND2_X1 U583 ( .A1(n637), .A2(G63), .ZN(n530) );
  XOR2_X1 U584 ( .A(KEYINPUT75), .B(n530), .Z(n532) );
  NAND2_X1 U585 ( .A1(n640), .A2(G51), .ZN(n531) );
  NAND2_X1 U586 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U587 ( .A(KEYINPUT6), .B(n533), .Z(n534) );
  NAND2_X1 U588 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U589 ( .A(KEYINPUT7), .B(n536), .ZN(G168) );
  NOR2_X1 U590 ( .A1(G2105), .A2(G2104), .ZN(n538) );
  XNOR2_X2 U591 ( .A(n538), .B(n537), .ZN(n882) );
  AND2_X1 U592 ( .A1(G2105), .A2(G2104), .ZN(n878) );
  NAND2_X1 U593 ( .A1(n878), .A2(G113), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U595 ( .A(n541), .B(KEYINPUT65), .ZN(n685) );
  INV_X1 U596 ( .A(G2105), .ZN(n542) );
  NOR2_X2 U597 ( .A1(G2104), .A2(n542), .ZN(n879) );
  NAND2_X1 U598 ( .A1(G125), .A2(n879), .ZN(n544) );
  NAND2_X1 U599 ( .A1(n883), .A2(G101), .ZN(n543) );
  AND2_X1 U600 ( .A1(n544), .A2(n520), .ZN(n683) );
  AND2_X1 U601 ( .A1(n685), .A2(n683), .ZN(G160) );
  NAND2_X1 U602 ( .A1(G60), .A2(n637), .ZN(n546) );
  NAND2_X1 U603 ( .A1(G47), .A2(n640), .ZN(n545) );
  NAND2_X1 U604 ( .A1(n546), .A2(n545), .ZN(n550) );
  NAND2_X1 U605 ( .A1(G85), .A2(n641), .ZN(n548) );
  NAND2_X1 U606 ( .A1(G72), .A2(n634), .ZN(n547) );
  NAND2_X1 U607 ( .A1(n548), .A2(n547), .ZN(n549) );
  OR2_X1 U608 ( .A1(n550), .A2(n549), .ZN(G290) );
  NAND2_X1 U609 ( .A1(G64), .A2(n637), .ZN(n552) );
  NAND2_X1 U610 ( .A1(G52), .A2(n640), .ZN(n551) );
  NAND2_X1 U611 ( .A1(n552), .A2(n551), .ZN(n558) );
  NAND2_X1 U612 ( .A1(n634), .A2(G77), .ZN(n553) );
  XNOR2_X1 U613 ( .A(n553), .B(KEYINPUT66), .ZN(n555) );
  NAND2_X1 U614 ( .A1(G90), .A2(n641), .ZN(n554) );
  NAND2_X1 U615 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U616 ( .A(KEYINPUT9), .B(n556), .Z(n557) );
  NOR2_X1 U617 ( .A1(n558), .A2(n557), .ZN(G171) );
  AND2_X1 U618 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U619 ( .A(G57), .ZN(G237) );
  INV_X1 U620 ( .A(G132), .ZN(G219) );
  XOR2_X1 U621 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U622 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n560) );
  NAND2_X1 U623 ( .A1(G7), .A2(G661), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n560), .B(n559), .ZN(G223) );
  INV_X1 U625 ( .A(G223), .ZN(n833) );
  NAND2_X1 U626 ( .A1(n833), .A2(G567), .ZN(n561) );
  XOR2_X1 U627 ( .A(KEYINPUT11), .B(n561), .Z(G234) );
  NAND2_X1 U628 ( .A1(n637), .A2(G56), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(KEYINPUT14), .ZN(n564) );
  NAND2_X1 U630 ( .A1(G43), .A2(n640), .ZN(n563) );
  NAND2_X1 U631 ( .A1(n564), .A2(n563), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n641), .A2(G81), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n565), .B(KEYINPUT12), .ZN(n567) );
  NAND2_X1 U634 ( .A1(G68), .A2(n634), .ZN(n566) );
  NAND2_X1 U635 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U636 ( .A(KEYINPUT72), .B(n568), .Z(n569) );
  XNOR2_X1 U637 ( .A(KEYINPUT13), .B(n569), .ZN(n570) );
  NOR2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U639 ( .A(KEYINPUT73), .B(n572), .ZN(n980) );
  INV_X1 U640 ( .A(G860), .ZN(n593) );
  OR2_X1 U641 ( .A1(n980), .A2(n593), .ZN(G153) );
  INV_X1 U642 ( .A(G171), .ZN(G301) );
  NAND2_X1 U643 ( .A1(G868), .A2(G301), .ZN(n582) );
  NAND2_X1 U644 ( .A1(G66), .A2(n637), .ZN(n574) );
  NAND2_X1 U645 ( .A1(G92), .A2(n641), .ZN(n573) );
  NAND2_X1 U646 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U647 ( .A(KEYINPUT74), .B(n575), .ZN(n579) );
  NAND2_X1 U648 ( .A1(G54), .A2(n640), .ZN(n577) );
  NAND2_X1 U649 ( .A1(G79), .A2(n634), .ZN(n576) );
  NAND2_X1 U650 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U651 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U652 ( .A(KEYINPUT15), .B(n580), .Z(n973) );
  OR2_X1 U653 ( .A1(n973), .A2(G868), .ZN(n581) );
  NAND2_X1 U654 ( .A1(n582), .A2(n581), .ZN(G284) );
  NAND2_X1 U655 ( .A1(G91), .A2(n641), .ZN(n584) );
  NAND2_X1 U656 ( .A1(G78), .A2(n634), .ZN(n583) );
  NAND2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n590) );
  NAND2_X1 U658 ( .A1(G53), .A2(n640), .ZN(n585) );
  XNOR2_X1 U659 ( .A(n585), .B(KEYINPUT68), .ZN(n588) );
  NAND2_X1 U660 ( .A1(G65), .A2(n637), .ZN(n586) );
  XOR2_X1 U661 ( .A(KEYINPUT67), .B(n586), .Z(n587) );
  NAND2_X1 U662 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U663 ( .A1(n590), .A2(n589), .ZN(n981) );
  XNOR2_X1 U664 ( .A(n981), .B(KEYINPUT69), .ZN(G299) );
  NAND2_X1 U665 ( .A1(G286), .A2(G868), .ZN(n592) );
  INV_X1 U666 ( .A(G868), .ZN(n657) );
  NAND2_X1 U667 ( .A1(G299), .A2(n657), .ZN(n591) );
  NAND2_X1 U668 ( .A1(n592), .A2(n591), .ZN(G297) );
  NAND2_X1 U669 ( .A1(n593), .A2(G559), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n594), .A2(n973), .ZN(n595) );
  XNOR2_X1 U671 ( .A(n595), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U672 ( .A1(G868), .A2(n980), .ZN(n596) );
  XNOR2_X1 U673 ( .A(KEYINPUT76), .B(n596), .ZN(n599) );
  NAND2_X1 U674 ( .A1(G868), .A2(n973), .ZN(n597) );
  NOR2_X1 U675 ( .A1(G559), .A2(n597), .ZN(n598) );
  NOR2_X1 U676 ( .A1(n599), .A2(n598), .ZN(G282) );
  NAND2_X1 U677 ( .A1(G111), .A2(n878), .ZN(n601) );
  NAND2_X1 U678 ( .A1(G135), .A2(n882), .ZN(n600) );
  NAND2_X1 U679 ( .A1(n601), .A2(n600), .ZN(n604) );
  NAND2_X1 U680 ( .A1(n879), .A2(G123), .ZN(n602) );
  XOR2_X1 U681 ( .A(KEYINPUT18), .B(n602), .Z(n603) );
  NOR2_X1 U682 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U683 ( .A1(n883), .A2(G99), .ZN(n605) );
  NAND2_X1 U684 ( .A1(n606), .A2(n605), .ZN(n931) );
  XNOR2_X1 U685 ( .A(n931), .B(G2096), .ZN(n607) );
  XNOR2_X1 U686 ( .A(n607), .B(KEYINPUT77), .ZN(n609) );
  INV_X1 U687 ( .A(G2100), .ZN(n608) );
  NAND2_X1 U688 ( .A1(n609), .A2(n608), .ZN(G156) );
  NAND2_X1 U689 ( .A1(G67), .A2(n637), .ZN(n611) );
  NAND2_X1 U690 ( .A1(G55), .A2(n640), .ZN(n610) );
  NAND2_X1 U691 ( .A1(n611), .A2(n610), .ZN(n614) );
  NAND2_X1 U692 ( .A1(n634), .A2(G80), .ZN(n612) );
  XOR2_X1 U693 ( .A(KEYINPUT78), .B(n612), .Z(n613) );
  NOR2_X1 U694 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U695 ( .A1(n641), .A2(G93), .ZN(n615) );
  NAND2_X1 U696 ( .A1(n616), .A2(n615), .ZN(n658) );
  NAND2_X1 U697 ( .A1(n973), .A2(G559), .ZN(n655) );
  XNOR2_X1 U698 ( .A(n980), .B(n655), .ZN(n617) );
  NOR2_X1 U699 ( .A1(n617), .A2(G860), .ZN(n618) );
  XNOR2_X1 U700 ( .A(n618), .B(KEYINPUT79), .ZN(n619) );
  XNOR2_X1 U701 ( .A(n658), .B(n619), .ZN(G145) );
  NAND2_X1 U702 ( .A1(G74), .A2(G651), .ZN(n620) );
  XNOR2_X1 U703 ( .A(n620), .B(KEYINPUT80), .ZN(n626) );
  NAND2_X1 U704 ( .A1(G49), .A2(n640), .ZN(n623) );
  NAND2_X1 U705 ( .A1(G87), .A2(n621), .ZN(n622) );
  NAND2_X1 U706 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U707 ( .A1(n637), .A2(n624), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n626), .A2(n625), .ZN(G288) );
  NAND2_X1 U709 ( .A1(G88), .A2(n641), .ZN(n628) );
  NAND2_X1 U710 ( .A1(G75), .A2(n634), .ZN(n627) );
  NAND2_X1 U711 ( .A1(n628), .A2(n627), .ZN(n631) );
  NAND2_X1 U712 ( .A1(G62), .A2(n637), .ZN(n629) );
  XNOR2_X1 U713 ( .A(KEYINPUT83), .B(n629), .ZN(n630) );
  NOR2_X1 U714 ( .A1(n631), .A2(n630), .ZN(n633) );
  NAND2_X1 U715 ( .A1(n640), .A2(G50), .ZN(n632) );
  NAND2_X1 U716 ( .A1(n633), .A2(n632), .ZN(G303) );
  INV_X1 U717 ( .A(G303), .ZN(G166) );
  NAND2_X1 U718 ( .A1(G73), .A2(n634), .ZN(n635) );
  XOR2_X1 U719 ( .A(KEYINPUT81), .B(n635), .Z(n636) );
  XNOR2_X1 U720 ( .A(n636), .B(KEYINPUT2), .ZN(n639) );
  NAND2_X1 U721 ( .A1(G61), .A2(n637), .ZN(n638) );
  NAND2_X1 U722 ( .A1(n639), .A2(n638), .ZN(n645) );
  NAND2_X1 U723 ( .A1(G48), .A2(n640), .ZN(n643) );
  NAND2_X1 U724 ( .A1(G86), .A2(n641), .ZN(n642) );
  NAND2_X1 U725 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U726 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U727 ( .A(KEYINPUT82), .B(n646), .Z(G305) );
  XNOR2_X1 U728 ( .A(KEYINPUT19), .B(KEYINPUT84), .ZN(n648) );
  XNOR2_X1 U729 ( .A(G290), .B(KEYINPUT85), .ZN(n647) );
  XNOR2_X1 U730 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U731 ( .A(n649), .B(G299), .ZN(n650) );
  XNOR2_X1 U732 ( .A(n650), .B(n658), .ZN(n651) );
  XNOR2_X1 U733 ( .A(G288), .B(n651), .ZN(n653) );
  XNOR2_X1 U734 ( .A(G166), .B(G305), .ZN(n652) );
  XNOR2_X1 U735 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U736 ( .A(n654), .B(n980), .ZN(n901) );
  XOR2_X1 U737 ( .A(n901), .B(n655), .Z(n656) );
  NAND2_X1 U738 ( .A1(G868), .A2(n656), .ZN(n660) );
  NAND2_X1 U739 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U740 ( .A1(n660), .A2(n659), .ZN(G295) );
  NAND2_X1 U741 ( .A1(G2078), .A2(G2084), .ZN(n661) );
  XOR2_X1 U742 ( .A(KEYINPUT20), .B(n661), .Z(n662) );
  NAND2_X1 U743 ( .A1(G2090), .A2(n662), .ZN(n663) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(n663), .ZN(n664) );
  NAND2_X1 U745 ( .A1(n664), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U746 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U747 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  NOR2_X1 U748 ( .A1(G220), .A2(G219), .ZN(n665) );
  XOR2_X1 U749 ( .A(KEYINPUT86), .B(n665), .Z(n666) );
  XNOR2_X1 U750 ( .A(n666), .B(KEYINPUT22), .ZN(n667) );
  NOR2_X1 U751 ( .A1(G218), .A2(n667), .ZN(n668) );
  NAND2_X1 U752 ( .A1(G96), .A2(n668), .ZN(n839) );
  NAND2_X1 U753 ( .A1(n839), .A2(G2106), .ZN(n674) );
  NAND2_X1 U754 ( .A1(G69), .A2(G120), .ZN(n669) );
  XOR2_X1 U755 ( .A(KEYINPUT87), .B(n669), .Z(n670) );
  NOR2_X1 U756 ( .A1(G237), .A2(n670), .ZN(n671) );
  XNOR2_X1 U757 ( .A(KEYINPUT88), .B(n671), .ZN(n672) );
  NAND2_X1 U758 ( .A1(n672), .A2(G108), .ZN(n838) );
  NAND2_X1 U759 ( .A1(G567), .A2(n838), .ZN(n673) );
  NAND2_X1 U760 ( .A1(n674), .A2(n673), .ZN(n840) );
  NAND2_X1 U761 ( .A1(G483), .A2(G661), .ZN(n675) );
  NOR2_X1 U762 ( .A1(n840), .A2(n675), .ZN(n837) );
  NAND2_X1 U763 ( .A1(n837), .A2(G36), .ZN(G176) );
  NAND2_X1 U764 ( .A1(G114), .A2(n878), .ZN(n677) );
  NAND2_X1 U765 ( .A1(G138), .A2(n882), .ZN(n676) );
  NAND2_X1 U766 ( .A1(n677), .A2(n676), .ZN(n681) );
  NAND2_X1 U767 ( .A1(G102), .A2(n883), .ZN(n679) );
  NAND2_X1 U768 ( .A1(G126), .A2(n879), .ZN(n678) );
  NAND2_X1 U769 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U770 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U771 ( .A(KEYINPUT89), .B(n682), .Z(G164) );
  AND2_X1 U772 ( .A1(G40), .A2(n683), .ZN(n684) );
  NAND2_X1 U773 ( .A1(n685), .A2(n684), .ZN(n686) );
  INV_X1 U774 ( .A(KEYINPUT94), .ZN(n687) );
  XNOR2_X1 U775 ( .A(n768), .B(n687), .ZN(n688) );
  NOR2_X1 U776 ( .A1(G164), .A2(G1384), .ZN(n767) );
  NAND2_X1 U777 ( .A1(n688), .A2(n767), .ZN(n689) );
  XNOR2_X2 U778 ( .A(n689), .B(KEYINPUT64), .ZN(n703) );
  NAND2_X1 U779 ( .A1(n703), .A2(G8), .ZN(n695) );
  INV_X1 U780 ( .A(KEYINPUT102), .ZN(n759) );
  NOR2_X1 U781 ( .A1(G1976), .A2(G288), .ZN(n988) );
  NAND2_X1 U782 ( .A1(n759), .A2(n988), .ZN(n692) );
  NAND2_X1 U783 ( .A1(n988), .A2(KEYINPUT33), .ZN(n690) );
  NAND2_X1 U784 ( .A1(n690), .A2(KEYINPUT102), .ZN(n691) );
  NAND2_X1 U785 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U786 ( .A1(n807), .A2(n693), .ZN(n766) );
  NOR2_X1 U787 ( .A1(n703), .A2(G2084), .ZN(n694) );
  XNOR2_X1 U788 ( .A(KEYINPUT96), .B(n694), .ZN(n751) );
  NOR2_X1 U789 ( .A1(G1966), .A2(n695), .ZN(n752) );
  INV_X1 U790 ( .A(KEYINPUT99), .ZN(n696) );
  XNOR2_X1 U791 ( .A(n697), .B(n696), .ZN(n698) );
  NAND2_X1 U792 ( .A1(n698), .A2(G8), .ZN(n699) );
  XNOR2_X1 U793 ( .A(n699), .B(n521), .ZN(n701) );
  XNOR2_X1 U794 ( .A(n702), .B(KEYINPUT101), .ZN(n708) );
  INV_X2 U795 ( .A(n704), .ZN(n724) );
  NOR2_X1 U796 ( .A1(G1961), .A2(n724), .ZN(n706) );
  XOR2_X1 U797 ( .A(KEYINPUT25), .B(G2078), .Z(n957) );
  NOR2_X1 U798 ( .A1(n737), .A2(n957), .ZN(n705) );
  NOR2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n734) );
  NAND2_X1 U800 ( .A1(n734), .A2(G301), .ZN(n707) );
  NAND2_X1 U801 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U802 ( .A(n709), .B(KEYINPUT31), .ZN(n750) );
  AND2_X1 U803 ( .A1(n724), .A2(G1996), .ZN(n710) );
  XNOR2_X1 U804 ( .A(n710), .B(KEYINPUT26), .ZN(n714) );
  NAND2_X1 U805 ( .A1(n737), .A2(G1341), .ZN(n712) );
  INV_X1 U806 ( .A(n980), .ZN(n711) );
  NAND2_X1 U807 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U808 ( .A1(n719), .A2(n973), .ZN(n718) );
  NAND2_X1 U809 ( .A1(G2067), .A2(n724), .ZN(n716) );
  NAND2_X1 U810 ( .A1(n737), .A2(G1348), .ZN(n715) );
  NAND2_X1 U811 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n721) );
  OR2_X1 U813 ( .A1(n719), .A2(n973), .ZN(n720) );
  NAND2_X1 U814 ( .A1(n721), .A2(n720), .ZN(n728) );
  NAND2_X1 U815 ( .A1(G2072), .A2(n724), .ZN(n723) );
  XOR2_X1 U816 ( .A(KEYINPUT97), .B(KEYINPUT27), .Z(n722) );
  XNOR2_X1 U817 ( .A(n723), .B(n722), .ZN(n726) );
  INV_X1 U818 ( .A(G1956), .ZN(n1001) );
  NOR2_X1 U819 ( .A1(n724), .A2(n1001), .ZN(n725) );
  NOR2_X1 U820 ( .A1(n726), .A2(n725), .ZN(n729) );
  NAND2_X1 U821 ( .A1(n729), .A2(n981), .ZN(n727) );
  NAND2_X1 U822 ( .A1(n728), .A2(n727), .ZN(n731) );
  NOR2_X1 U823 ( .A1(n729), .A2(n981), .ZN(n730) );
  NAND2_X1 U824 ( .A1(n731), .A2(n522), .ZN(n733) );
  XOR2_X1 U825 ( .A(KEYINPUT29), .B(KEYINPUT98), .Z(n732) );
  XNOR2_X1 U826 ( .A(n733), .B(n732), .ZN(n736) );
  OR2_X1 U827 ( .A1(n734), .A2(G301), .ZN(n735) );
  NAND2_X1 U828 ( .A1(n736), .A2(n735), .ZN(n749) );
  INV_X1 U829 ( .A(G8), .ZN(n742) );
  NOR2_X1 U830 ( .A1(G1971), .A2(n807), .ZN(n739) );
  NOR2_X1 U831 ( .A1(n737), .A2(G2090), .ZN(n738) );
  NOR2_X1 U832 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U833 ( .A1(n740), .A2(G303), .ZN(n741) );
  OR2_X1 U834 ( .A1(n742), .A2(n741), .ZN(n744) );
  AND2_X1 U835 ( .A1(n749), .A2(n744), .ZN(n743) );
  NAND2_X1 U836 ( .A1(n750), .A2(n743), .ZN(n747) );
  INV_X1 U837 ( .A(n744), .ZN(n745) );
  OR2_X1 U838 ( .A1(n745), .A2(G286), .ZN(n746) );
  NAND2_X1 U839 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U840 ( .A(n748), .B(KEYINPUT32), .ZN(n756) );
  NAND2_X1 U841 ( .A1(n750), .A2(n749), .ZN(n754) );
  AND2_X1 U842 ( .A1(n751), .A2(G8), .ZN(n753) );
  NAND2_X1 U843 ( .A1(n754), .A2(n523), .ZN(n755) );
  NAND2_X1 U844 ( .A1(n756), .A2(n755), .ZN(n802) );
  NOR2_X1 U845 ( .A1(G1971), .A2(G303), .ZN(n757) );
  NOR2_X1 U846 ( .A1(n757), .A2(n988), .ZN(n758) );
  NAND2_X1 U847 ( .A1(n802), .A2(n758), .ZN(n763) );
  OR2_X1 U848 ( .A1(n807), .A2(n759), .ZN(n761) );
  NAND2_X1 U849 ( .A1(G1976), .A2(G288), .ZN(n991) );
  NOR2_X1 U850 ( .A1(n764), .A2(KEYINPUT33), .ZN(n765) );
  NOR2_X1 U851 ( .A1(n766), .A2(n765), .ZN(n799) );
  XOR2_X1 U852 ( .A(G1981), .B(G305), .Z(n976) );
  NOR2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n828) );
  XNOR2_X1 U854 ( .A(G2067), .B(KEYINPUT37), .ZN(n825) );
  NAND2_X1 U855 ( .A1(G140), .A2(n882), .ZN(n770) );
  NAND2_X1 U856 ( .A1(G104), .A2(n883), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U858 ( .A(KEYINPUT34), .B(n771), .ZN(n777) );
  NAND2_X1 U859 ( .A1(n878), .A2(G116), .ZN(n772) );
  XOR2_X1 U860 ( .A(KEYINPUT91), .B(n772), .Z(n774) );
  NAND2_X1 U861 ( .A1(n879), .A2(G128), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U863 ( .A(KEYINPUT35), .B(n775), .Z(n776) );
  NOR2_X1 U864 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U865 ( .A(KEYINPUT36), .B(n778), .ZN(n898) );
  NOR2_X1 U866 ( .A1(n825), .A2(n898), .ZN(n938) );
  NAND2_X1 U867 ( .A1(n828), .A2(n938), .ZN(n823) );
  INV_X1 U868 ( .A(n823), .ZN(n796) );
  NAND2_X1 U869 ( .A1(G95), .A2(n883), .ZN(n780) );
  NAND2_X1 U870 ( .A1(G119), .A2(n879), .ZN(n779) );
  NAND2_X1 U871 ( .A1(n780), .A2(n779), .ZN(n783) );
  NAND2_X1 U872 ( .A1(n882), .A2(G131), .ZN(n781) );
  XOR2_X1 U873 ( .A(KEYINPUT92), .B(n781), .Z(n782) );
  NOR2_X1 U874 ( .A1(n783), .A2(n782), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n878), .A2(G107), .ZN(n784) );
  NAND2_X1 U876 ( .A1(n785), .A2(n784), .ZN(n893) );
  NAND2_X1 U877 ( .A1(G1991), .A2(n893), .ZN(n794) );
  NAND2_X1 U878 ( .A1(G117), .A2(n878), .ZN(n787) );
  NAND2_X1 U879 ( .A1(G141), .A2(n882), .ZN(n786) );
  NAND2_X1 U880 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n883), .A2(G105), .ZN(n788) );
  XOR2_X1 U882 ( .A(KEYINPUT38), .B(n788), .Z(n789) );
  NOR2_X1 U883 ( .A1(n790), .A2(n789), .ZN(n792) );
  NAND2_X1 U884 ( .A1(n879), .A2(G129), .ZN(n791) );
  NAND2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n889) );
  NAND2_X1 U886 ( .A1(G1996), .A2(n889), .ZN(n793) );
  NAND2_X1 U887 ( .A1(n794), .A2(n793), .ZN(n929) );
  NAND2_X1 U888 ( .A1(n828), .A2(n929), .ZN(n795) );
  XNOR2_X1 U889 ( .A(n795), .B(KEYINPUT93), .ZN(n820) );
  OR2_X1 U890 ( .A1(n796), .A2(n820), .ZN(n811) );
  INV_X1 U891 ( .A(n811), .ZN(n797) );
  AND2_X1 U892 ( .A1(n976), .A2(n797), .ZN(n798) );
  NAND2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n813) );
  NOR2_X1 U894 ( .A1(G2090), .A2(G303), .ZN(n800) );
  NAND2_X1 U895 ( .A1(G8), .A2(n800), .ZN(n801) );
  NAND2_X1 U896 ( .A1(n802), .A2(n801), .ZN(n803) );
  AND2_X1 U897 ( .A1(n807), .A2(n803), .ZN(n809) );
  NOR2_X1 U898 ( .A1(G1981), .A2(G305), .ZN(n804) );
  XNOR2_X1 U899 ( .A(n804), .B(KEYINPUT24), .ZN(n805) );
  XNOR2_X1 U900 ( .A(n805), .B(KEYINPUT95), .ZN(n806) );
  NOR2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n808) );
  NOR2_X1 U902 ( .A1(n809), .A2(n808), .ZN(n810) );
  OR2_X1 U903 ( .A1(n811), .A2(n810), .ZN(n812) );
  AND2_X1 U904 ( .A1(n813), .A2(n812), .ZN(n814) );
  XNOR2_X1 U905 ( .A(n814), .B(KEYINPUT103), .ZN(n816) );
  XNOR2_X1 U906 ( .A(G1986), .B(G290), .ZN(n985) );
  NAND2_X1 U907 ( .A1(n985), .A2(n828), .ZN(n815) );
  NAND2_X1 U908 ( .A1(n816), .A2(n815), .ZN(n831) );
  NOR2_X1 U909 ( .A1(G1996), .A2(n889), .ZN(n927) );
  NOR2_X1 U910 ( .A1(G1991), .A2(n893), .ZN(n930) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n817) );
  XNOR2_X1 U912 ( .A(KEYINPUT104), .B(n817), .ZN(n818) );
  NOR2_X1 U913 ( .A1(n930), .A2(n818), .ZN(n819) );
  NOR2_X1 U914 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U915 ( .A1(n927), .A2(n821), .ZN(n822) );
  XNOR2_X1 U916 ( .A(n822), .B(KEYINPUT39), .ZN(n824) );
  NAND2_X1 U917 ( .A1(n824), .A2(n823), .ZN(n826) );
  NAND2_X1 U918 ( .A1(n825), .A2(n898), .ZN(n943) );
  NAND2_X1 U919 ( .A1(n826), .A2(n943), .ZN(n827) );
  XOR2_X1 U920 ( .A(KEYINPUT105), .B(n827), .Z(n829) );
  NAND2_X1 U921 ( .A1(n829), .A2(n828), .ZN(n830) );
  NAND2_X1 U922 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U923 ( .A(KEYINPUT40), .B(n832), .ZN(G329) );
  NAND2_X1 U924 ( .A1(n833), .A2(G2106), .ZN(n834) );
  XOR2_X1 U925 ( .A(KEYINPUT107), .B(n834), .Z(G217) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U927 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U929 ( .A1(n837), .A2(n836), .ZN(G188) );
  XOR2_X1 U930 ( .A(G120), .B(KEYINPUT108), .Z(G236) );
  INV_X1 U932 ( .A(G108), .ZN(G238) );
  INV_X1 U933 ( .A(G69), .ZN(G235) );
  NOR2_X1 U934 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  INV_X1 U936 ( .A(n840), .ZN(G319) );
  XOR2_X1 U937 ( .A(KEYINPUT110), .B(KEYINPUT109), .Z(n842) );
  XNOR2_X1 U938 ( .A(G2678), .B(KEYINPUT43), .ZN(n841) );
  XNOR2_X1 U939 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U940 ( .A(KEYINPUT42), .B(G2090), .Z(n844) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2072), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U943 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U944 ( .A(G2096), .B(G2100), .ZN(n847) );
  XNOR2_X1 U945 ( .A(n848), .B(n847), .ZN(n850) );
  XOR2_X1 U946 ( .A(G2078), .B(G2084), .Z(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(G227) );
  XOR2_X1 U948 ( .A(G1981), .B(G1961), .Z(n852) );
  XNOR2_X1 U949 ( .A(G1986), .B(G1966), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U951 ( .A(n853), .B(KEYINPUT41), .Z(n855) );
  XNOR2_X1 U952 ( .A(G1996), .B(G1991), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U954 ( .A(G2474), .B(G1976), .Z(n857) );
  XNOR2_X1 U955 ( .A(G1956), .B(G1971), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n859), .B(n858), .ZN(G229) );
  NAND2_X1 U958 ( .A1(G112), .A2(n878), .ZN(n861) );
  NAND2_X1 U959 ( .A1(G100), .A2(n883), .ZN(n860) );
  NAND2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n867) );
  NAND2_X1 U961 ( .A1(n879), .A2(G124), .ZN(n862) );
  XNOR2_X1 U962 ( .A(n862), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U963 ( .A1(G136), .A2(n882), .ZN(n863) );
  NAND2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U965 ( .A(KEYINPUT111), .B(n865), .Z(n866) );
  NOR2_X1 U966 ( .A1(n867), .A2(n866), .ZN(G162) );
  XNOR2_X1 U967 ( .A(KEYINPUT48), .B(KEYINPUT112), .ZN(n869) );
  XNOR2_X1 U968 ( .A(n931), .B(KEYINPUT46), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U970 ( .A(G160), .B(n870), .ZN(n897) );
  NAND2_X1 U971 ( .A1(G139), .A2(n882), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G103), .A2(n883), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n877) );
  NAND2_X1 U974 ( .A1(G115), .A2(n878), .ZN(n874) );
  NAND2_X1 U975 ( .A1(G127), .A2(n879), .ZN(n873) );
  NAND2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U977 ( .A(KEYINPUT47), .B(n875), .Z(n876) );
  NOR2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n921) );
  NAND2_X1 U979 ( .A1(G118), .A2(n878), .ZN(n881) );
  NAND2_X1 U980 ( .A1(G130), .A2(n879), .ZN(n880) );
  NAND2_X1 U981 ( .A1(n881), .A2(n880), .ZN(n888) );
  NAND2_X1 U982 ( .A1(G142), .A2(n882), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G106), .A2(n883), .ZN(n884) );
  NAND2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n886) );
  XOR2_X1 U985 ( .A(n886), .B(KEYINPUT45), .Z(n887) );
  NOR2_X1 U986 ( .A1(n888), .A2(n887), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n890), .B(n889), .ZN(n891) );
  XNOR2_X1 U988 ( .A(n921), .B(n891), .ZN(n895) );
  XOR2_X1 U989 ( .A(G164), .B(G162), .Z(n892) );
  XNOR2_X1 U990 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n897), .B(n896), .ZN(n899) );
  XNOR2_X1 U993 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U994 ( .A1(G37), .A2(n900), .ZN(G395) );
  XNOR2_X1 U995 ( .A(n973), .B(G286), .ZN(n902) );
  XNOR2_X1 U996 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U997 ( .A(n903), .B(G171), .ZN(n904) );
  NOR2_X1 U998 ( .A1(G37), .A2(n904), .ZN(G397) );
  XOR2_X1 U999 ( .A(G2438), .B(KEYINPUT106), .Z(n906) );
  XNOR2_X1 U1000 ( .A(G2443), .B(G2430), .ZN(n905) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n907) );
  XOR2_X1 U1002 ( .A(n907), .B(G2435), .Z(n909) );
  XNOR2_X1 U1003 ( .A(G1348), .B(G1341), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(n909), .B(n908), .ZN(n913) );
  XOR2_X1 U1005 ( .A(G2451), .B(G2427), .Z(n911) );
  XNOR2_X1 U1006 ( .A(G2454), .B(G2446), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n912) );
  XOR2_X1 U1008 ( .A(n913), .B(n912), .Z(n914) );
  NAND2_X1 U1009 ( .A1(G14), .A2(n914), .ZN(n920) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n920), .ZN(n917) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n915) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n915), .ZN(n916) );
  NOR2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(n919) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1015 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G96), .ZN(G221) );
  INV_X1 U1018 ( .A(n920), .ZN(G401) );
  XNOR2_X1 U1019 ( .A(G2072), .B(n921), .ZN(n924) );
  XNOR2_X1 U1020 ( .A(G164), .B(G2078), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(n922), .B(KEYINPUT114), .ZN(n923) );
  NAND2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(n925), .B(KEYINPUT50), .ZN(n941) );
  XOR2_X1 U1024 ( .A(G2090), .B(G162), .Z(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1026 ( .A(KEYINPUT51), .B(n928), .Z(n936) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n932) );
  NAND2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n934) );
  XOR2_X1 U1029 ( .A(G160), .B(G2084), .Z(n933) );
  NOR2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(n939), .B(KEYINPUT113), .ZN(n940) );
  NOR2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n946) );
  XNOR2_X1 U1036 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n944) );
  XNOR2_X1 U1037 ( .A(n944), .B(KEYINPUT52), .ZN(n945) );
  XNOR2_X1 U1038 ( .A(n946), .B(n945), .ZN(n947) );
  INV_X1 U1039 ( .A(KEYINPUT55), .ZN(n969) );
  NAND2_X1 U1040 ( .A1(n947), .A2(n969), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n948), .A2(G29), .ZN(n1031) );
  XOR2_X1 U1042 ( .A(KEYINPUT118), .B(G34), .Z(n950) );
  XNOR2_X1 U1043 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(n950), .B(n949), .ZN(n951) );
  XNOR2_X1 U1045 ( .A(G2084), .B(n951), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(G2090), .B(G35), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n967) );
  XOR2_X1 U1048 ( .A(G1991), .B(G25), .Z(n954) );
  NAND2_X1 U1049 ( .A1(n954), .A2(G28), .ZN(n963) );
  XNOR2_X1 U1050 ( .A(G2067), .B(G26), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(G33), .B(G2072), .ZN(n955) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n961) );
  XNOR2_X1 U1053 ( .A(G1996), .B(G32), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(G27), .B(n957), .ZN(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(KEYINPUT117), .B(KEYINPUT53), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(n965), .B(n964), .ZN(n966) );
  NAND2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(n969), .B(n968), .ZN(n971) );
  INV_X1 U1062 ( .A(G29), .ZN(n970) );
  NAND2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1064 ( .A1(G11), .A2(n972), .ZN(n1029) );
  XNOR2_X1 U1065 ( .A(G16), .B(KEYINPUT56), .ZN(n999) );
  XOR2_X1 U1066 ( .A(G1348), .B(n973), .Z(n975) );
  XOR2_X1 U1067 ( .A(G171), .B(G1961), .Z(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n997) );
  XNOR2_X1 U1069 ( .A(G1966), .B(G168), .ZN(n977) );
  NAND2_X1 U1070 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(n978), .B(KEYINPUT120), .ZN(n979) );
  XNOR2_X1 U1072 ( .A(KEYINPUT57), .B(n979), .ZN(n987) );
  XOR2_X1 U1073 ( .A(n980), .B(G1341), .Z(n983) );
  XNOR2_X1 U1074 ( .A(n981), .B(G1956), .ZN(n982) );
  NAND2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n995) );
  XOR2_X1 U1078 ( .A(n988), .B(KEYINPUT121), .Z(n990) );
  XOR2_X1 U1079 ( .A(G166), .B(G1971), .Z(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(KEYINPUT122), .B(n993), .ZN(n994) );
  NOR2_X1 U1083 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1084 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1085 ( .A1(n999), .A2(n998), .ZN(n1027) );
  INV_X1 U1086 ( .A(G16), .ZN(n1025) );
  XOR2_X1 U1087 ( .A(G1961), .B(G5), .Z(n1014) );
  XNOR2_X1 U1088 ( .A(KEYINPUT59), .B(G1348), .ZN(n1000) );
  XNOR2_X1 U1089 ( .A(n1000), .B(G4), .ZN(n1007) );
  XOR2_X1 U1090 ( .A(G1341), .B(G19), .Z(n1003) );
  XNOR2_X1 U1091 ( .A(n1001), .B(G20), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(G6), .B(G1981), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  XOR2_X1 U1096 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n1008) );
  XNOR2_X1 U1097 ( .A(n1009), .B(n1008), .ZN(n1011) );
  XNOR2_X1 U1098 ( .A(G1966), .B(G21), .ZN(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1100 ( .A(KEYINPUT124), .B(n1012), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1022) );
  XOR2_X1 U1102 ( .A(G1986), .B(G24), .Z(n1018) );
  XNOR2_X1 U1103 ( .A(G1971), .B(G22), .ZN(n1016) );
  XNOR2_X1 U1104 ( .A(G23), .B(G1976), .ZN(n1015) );
  NOR2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1107 ( .A(KEYINPUT125), .B(n1019), .Z(n1020) );
  XNOR2_X1 U1108 ( .A(KEYINPUT58), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1110 ( .A(KEYINPUT61), .B(n1023), .ZN(n1024) );
  NAND2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1114 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1115 ( .A(n1032), .B(KEYINPUT62), .ZN(n1033) );
  XOR2_X1 U1116 ( .A(KEYINPUT126), .B(n1033), .Z(G311) );
  XNOR2_X1 U1117 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

