

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743;

  XNOR2_X1 U372 ( .A(n614), .B(KEYINPUT32), .ZN(n741) );
  NAND2_X1 U373 ( .A1(n616), .A2(n613), .ZN(n614) );
  INV_X1 U374 ( .A(n592), .ZN(n671) );
  NOR2_X1 U375 ( .A1(n699), .A2(G902), .ZN(n509) );
  OR2_X1 U376 ( .A1(n703), .A2(G902), .ZN(n427) );
  AND2_X2 U377 ( .A1(n596), .A2(n355), .ZN(n600) );
  NOR2_X2 U378 ( .A1(n618), .A2(KEYINPUT44), .ZN(n409) );
  XOR2_X2 U379 ( .A(KEYINPUT70), .B(G110), .Z(n499) );
  XNOR2_X2 U380 ( .A(n596), .B(KEYINPUT90), .ZN(n608) );
  OR2_X2 U381 ( .A1(n608), .A2(n435), .ZN(n429) );
  INV_X2 U382 ( .A(n664), .ZN(n510) );
  XNOR2_X2 U383 ( .A(n426), .B(n425), .ZN(n664) );
  NOR2_X1 U384 ( .A1(n592), .A2(n553), .ZN(n543) );
  XNOR2_X1 U385 ( .A(n380), .B(n515), .ZN(n715) );
  INV_X1 U386 ( .A(G953), .ZN(n710) );
  INV_X2 U387 ( .A(G122), .ZN(n371) );
  XNOR2_X2 U388 ( .A(n557), .B(KEYINPUT1), .ZN(n577) );
  NOR2_X1 U389 ( .A1(n407), .A2(n405), .ZN(n389) );
  AND2_X1 U390 ( .A1(n392), .A2(n390), .ZN(n723) );
  OR2_X1 U391 ( .A1(n560), .A2(n414), .ZN(n438) );
  AND2_X1 U392 ( .A1(n429), .A2(n434), .ZN(n428) );
  NOR2_X1 U393 ( .A1(n440), .A2(n368), .ZN(n566) );
  XNOR2_X1 U394 ( .A(n393), .B(n352), .ZN(n515) );
  XOR2_X1 U395 ( .A(G137), .B(G140), .Z(n500) );
  XNOR2_X1 U396 ( .A(n459), .B(n394), .ZN(n393) );
  XNOR2_X1 U397 ( .A(G119), .B(G116), .ZN(n459) );
  XNOR2_X1 U398 ( .A(n722), .B(n507), .ZN(n514) );
  INV_X1 U399 ( .A(G146), .ZN(n507) );
  INV_X1 U400 ( .A(KEYINPUT33), .ZN(n385) );
  INV_X1 U401 ( .A(KEYINPUT34), .ZN(n435) );
  XNOR2_X1 U402 ( .A(n446), .B(KEYINPUT67), .ZN(n506) );
  INV_X1 U403 ( .A(G131), .ZN(n446) );
  NOR2_X1 U404 ( .A1(n634), .A2(n637), .ZN(n656) );
  INV_X1 U405 ( .A(KEYINPUT65), .ZN(n425) );
  NAND2_X1 U406 ( .A1(n661), .A2(n662), .ZN(n426) );
  XNOR2_X1 U407 ( .A(n522), .B(G472), .ZN(n402) );
  NOR2_X1 U408 ( .A1(n402), .A2(G902), .ZN(n398) );
  AND2_X1 U409 ( .A1(n622), .A2(n402), .ZN(n401) );
  NOR2_X1 U410 ( .A1(n419), .A2(n418), .ZN(n417) );
  OR2_X1 U411 ( .A1(n739), .A2(n576), .ZN(n418) );
  XNOR2_X1 U412 ( .A(KEYINPUT4), .B(KEYINPUT18), .ZN(n454) );
  XNOR2_X1 U413 ( .A(n499), .B(n383), .ZN(n382) );
  INV_X1 U414 ( .A(KEYINPUT17), .ZN(n383) );
  INV_X1 U415 ( .A(n463), .ZN(n455) );
  INV_X1 U416 ( .A(n542), .ZN(n441) );
  XNOR2_X1 U417 ( .A(n379), .B(n467), .ZN(n380) );
  XNOR2_X1 U418 ( .A(n475), .B(n458), .ZN(n379) );
  XOR2_X1 U419 ( .A(KEYINPUT16), .B(KEYINPUT71), .Z(n458) );
  XOR2_X1 U420 ( .A(KEYINPUT66), .B(KEYINPUT8), .Z(n477) );
  XNOR2_X1 U421 ( .A(n479), .B(n423), .ZN(n422) );
  XNOR2_X1 U422 ( .A(n480), .B(n424), .ZN(n423) );
  XNOR2_X1 U423 ( .A(G116), .B(G134), .ZN(n424) );
  XNOR2_X1 U424 ( .A(n472), .B(n471), .ZN(n701) );
  XNOR2_X1 U425 ( .A(n465), .B(n376), .ZN(n472) );
  XNOR2_X1 U426 ( .A(n421), .B(n420), .ZN(n676) );
  XNOR2_X1 U427 ( .A(n545), .B(KEYINPUT105), .ZN(n420) );
  OR2_X1 U428 ( .A1(n654), .A2(n655), .ZN(n421) );
  XNOR2_X1 U429 ( .A(n537), .B(KEYINPUT39), .ZN(n538) );
  AND2_X1 U430 ( .A1(n566), .A2(n651), .ZN(n539) );
  INV_X1 U431 ( .A(n609), .ZN(n434) );
  INV_X1 U432 ( .A(KEYINPUT22), .ZN(n599) );
  BUF_X1 U433 ( .A(n661), .Z(n378) );
  XNOR2_X1 U434 ( .A(n514), .B(n370), .ZN(n699) );
  XNOR2_X1 U435 ( .A(n505), .B(n354), .ZN(n370) );
  XNOR2_X1 U436 ( .A(G101), .B(KEYINPUT3), .ZN(n394) );
  XNOR2_X1 U437 ( .A(G134), .B(KEYINPUT4), .ZN(n444) );
  NAND2_X1 U438 ( .A1(G234), .A2(G237), .ZN(n525) );
  NOR2_X1 U439 ( .A1(G953), .A2(G237), .ZN(n516) );
  XNOR2_X1 U440 ( .A(n604), .B(n406), .ZN(n405) );
  INV_X1 U441 ( .A(KEYINPUT99), .ZN(n406) );
  XOR2_X1 U442 ( .A(G113), .B(G104), .Z(n467) );
  XNOR2_X1 U443 ( .A(n466), .B(n377), .ZN(n376) );
  INV_X1 U444 ( .A(G122), .ZN(n377) );
  XNOR2_X1 U445 ( .A(n445), .B(n442), .ZN(n722) );
  XNOR2_X1 U446 ( .A(n444), .B(n443), .ZN(n442) );
  XNOR2_X1 U447 ( .A(n478), .B(n506), .ZN(n445) );
  INV_X1 U448 ( .A(KEYINPUT68), .ZN(n443) );
  OR2_X1 U449 ( .A1(G237), .A2(G902), .ZN(n534) );
  XNOR2_X1 U450 ( .A(n448), .B(n447), .ZN(n605) );
  INV_X1 U451 ( .A(KEYINPUT73), .ZN(n447) );
  XNOR2_X1 U452 ( .A(n474), .B(n473), .ZN(n564) );
  NAND2_X1 U453 ( .A1(n400), .A2(n397), .ZN(n592) );
  NOR2_X1 U454 ( .A1(n401), .A2(n353), .ZN(n400) );
  NAND2_X1 U455 ( .A1(n399), .A2(n398), .ZN(n397) );
  NOR2_X1 U456 ( .A1(n565), .A2(n564), .ZN(n598) );
  XNOR2_X1 U457 ( .A(G113), .B(G137), .ZN(n511) );
  NOR2_X1 U458 ( .A1(n732), .A2(n391), .ZN(n390) );
  INV_X1 U459 ( .A(n647), .ZN(n391) );
  XNOR2_X1 U460 ( .A(G110), .B(KEYINPUT24), .ZN(n485) );
  XNOR2_X1 U461 ( .A(n502), .B(n501), .ZN(n503) );
  INV_X1 U462 ( .A(G107), .ZN(n501) );
  XNOR2_X1 U463 ( .A(G101), .B(G104), .ZN(n502) );
  XNOR2_X1 U464 ( .A(n455), .B(n452), .ZN(n456) );
  XNOR2_X1 U465 ( .A(n523), .B(n524), .ZN(n368) );
  OR2_X1 U466 ( .A1(n593), .A2(n441), .ZN(n440) );
  XNOR2_X1 U467 ( .A(n481), .B(n422), .ZN(n482) );
  NOR2_X1 U468 ( .A1(n676), .A2(n562), .ZN(n546) );
  NOR2_X1 U469 ( .A1(n648), .A2(n435), .ZN(n433) );
  NOR2_X1 U470 ( .A1(n562), .A2(n589), .ZN(n638) );
  XNOR2_X1 U471 ( .A(n412), .B(n411), .ZN(n629) );
  INV_X1 U472 ( .A(KEYINPUT95), .ZN(n411) );
  NAND2_X1 U473 ( .A1(n608), .A2(n413), .ZN(n412) );
  NOR2_X1 U474 ( .A1(n593), .A2(n671), .ZN(n413) );
  INV_X1 U475 ( .A(KEYINPUT60), .ZN(n366) );
  XNOR2_X1 U476 ( .A(n697), .B(n384), .ZN(n700) );
  XNOR2_X1 U477 ( .A(n699), .B(n698), .ZN(n384) );
  INV_X1 U478 ( .A(KEYINPUT56), .ZN(n364) );
  XOR2_X1 U479 ( .A(n496), .B(n495), .Z(n351) );
  XNOR2_X1 U480 ( .A(KEYINPUT69), .B(KEYINPUT87), .ZN(n352) );
  AND2_X1 U481 ( .A1(n402), .A2(G902), .ZN(n353) );
  AND2_X1 U482 ( .A1(G227), .A2(n710), .ZN(n354) );
  AND2_X1 U483 ( .A1(n598), .A2(n662), .ZN(n355) );
  XNOR2_X1 U484 ( .A(n701), .B(KEYINPUT59), .ZN(n356) );
  XOR2_X1 U485 ( .A(n624), .B(KEYINPUT118), .Z(n357) );
  XOR2_X1 U486 ( .A(n462), .B(n461), .Z(n358) );
  XOR2_X1 U487 ( .A(n622), .B(KEYINPUT62), .Z(n359) );
  NOR2_X1 U488 ( .A1(G952), .A2(n710), .ZN(n708) );
  INV_X1 U489 ( .A(n708), .ZN(n374) );
  XOR2_X1 U490 ( .A(G902), .B(KEYINPUT15), .Z(n532) );
  NAND2_X1 U491 ( .A1(n389), .A2(n388), .ZN(n387) );
  XNOR2_X1 U492 ( .A(n382), .B(n360), .ZN(n457) );
  XNOR2_X1 U493 ( .A(n478), .B(n454), .ZN(n360) );
  XNOR2_X1 U494 ( .A(n361), .B(KEYINPUT119), .ZN(G63) );
  NAND2_X1 U495 ( .A1(n369), .A2(n374), .ZN(n361) );
  XNOR2_X2 U496 ( .A(n688), .B(KEYINPUT2), .ZN(n362) );
  NAND2_X2 U497 ( .A1(n709), .A2(n723), .ZN(n688) );
  AND2_X4 U498 ( .A1(n362), .A2(n532), .ZN(n704) );
  XNOR2_X1 U499 ( .A(n363), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U500 ( .A1(n372), .A2(n374), .ZN(n363) );
  XNOR2_X1 U501 ( .A(n365), .B(n364), .ZN(G51) );
  NAND2_X1 U502 ( .A1(n373), .A2(n374), .ZN(n365) );
  XNOR2_X1 U503 ( .A(n367), .B(n366), .ZN(G60) );
  NAND2_X1 U504 ( .A1(n375), .A2(n374), .ZN(n367) );
  XNOR2_X1 U505 ( .A(n625), .B(n357), .ZN(n369) );
  XNOR2_X1 U506 ( .A(n702), .B(n356), .ZN(n375) );
  XNOR2_X1 U507 ( .A(n623), .B(n359), .ZN(n372) );
  XNOR2_X1 U508 ( .A(n621), .B(n358), .ZN(n373) );
  XNOR2_X1 U509 ( .A(n381), .B(n610), .ZN(n736) );
  XNOR2_X2 U510 ( .A(n371), .B(G107), .ZN(n475) );
  NOR2_X2 U511 ( .A1(n431), .A2(n433), .ZN(n381) );
  XNOR2_X2 U512 ( .A(n590), .B(KEYINPUT0), .ZN(n596) );
  XNOR2_X2 U513 ( .A(n387), .B(KEYINPUT45), .ZN(n709) );
  XNOR2_X2 U514 ( .A(n386), .B(n385), .ZN(n648) );
  NOR2_X2 U515 ( .A1(n606), .A2(n607), .ZN(n386) );
  XNOR2_X1 U516 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U517 ( .A(n404), .B(KEYINPUT84), .ZN(n388) );
  NAND2_X1 U518 ( .A1(n437), .A2(n436), .ZN(n392) );
  INV_X1 U519 ( .A(n515), .ZN(n520) );
  NAND2_X1 U520 ( .A1(n735), .A2(n395), .ZN(n569) );
  NAND2_X1 U521 ( .A1(n396), .A2(KEYINPUT47), .ZN(n395) );
  NAND2_X1 U522 ( .A1(n638), .A2(n563), .ZN(n396) );
  INV_X1 U523 ( .A(n622), .ZN(n399) );
  XNOR2_X2 U524 ( .A(n561), .B(n451), .ZN(n589) );
  XNOR2_X2 U525 ( .A(n403), .B(KEYINPUT86), .ZN(n561) );
  NAND2_X1 U526 ( .A1(n552), .A2(n650), .ZN(n403) );
  XNOR2_X1 U527 ( .A(n536), .B(n535), .ZN(n552) );
  NAND2_X1 U528 ( .A1(n736), .A2(KEYINPUT44), .ZN(n404) );
  NAND2_X1 U529 ( .A1(n408), .A2(n617), .ZN(n407) );
  NAND2_X1 U530 ( .A1(n410), .A2(n409), .ZN(n408) );
  INV_X1 U531 ( .A(n736), .ZN(n410) );
  XNOR2_X2 U532 ( .A(G143), .B(G128), .ZN(n478) );
  INV_X1 U533 ( .A(n560), .ZN(n416) );
  NAND2_X1 U534 ( .A1(n575), .A2(n415), .ZN(n414) );
  INV_X1 U535 ( .A(n575), .ZN(n419) );
  INV_X1 U536 ( .A(n739), .ZN(n415) );
  NAND2_X1 U537 ( .A1(n417), .A2(n416), .ZN(n436) );
  NOR2_X1 U538 ( .A1(n624), .A2(G902), .ZN(n484) );
  NOR2_X2 U539 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X2 U540 ( .A(n427), .B(n351), .ZN(n661) );
  NAND2_X1 U541 ( .A1(n648), .A2(n432), .ZN(n430) );
  NAND2_X1 U542 ( .A1(n430), .A2(n428), .ZN(n431) );
  AND2_X1 U543 ( .A1(n608), .A2(n435), .ZN(n432) );
  NAND2_X1 U544 ( .A1(n438), .A2(n576), .ZN(n437) );
  NOR2_X1 U545 ( .A1(n439), .A2(n734), .ZN(n550) );
  XNOR2_X1 U546 ( .A(n439), .B(n743), .ZN(G33) );
  XNOR2_X1 U547 ( .A(n549), .B(KEYINPUT40), .ZN(n439) );
  INV_X1 U548 ( .A(n577), .ZN(n665) );
  NAND2_X1 U549 ( .A1(n510), .A2(n577), .ZN(n448) );
  XNOR2_X1 U550 ( .A(n449), .B(n514), .ZN(n622) );
  XNOR2_X1 U551 ( .A(n521), .B(n513), .ZN(n449) );
  BUF_X1 U552 ( .A(n688), .Z(n691) );
  XNOR2_X1 U553 ( .A(n539), .B(n538), .ZN(n548) );
  XOR2_X1 U554 ( .A(n469), .B(n468), .Z(n450) );
  XOR2_X1 U555 ( .A(KEYINPUT19), .B(KEYINPUT64), .Z(n451) );
  AND2_X1 U556 ( .A1(G224), .A2(n710), .ZN(n452) );
  AND2_X1 U557 ( .A1(n491), .A2(G221), .ZN(n453) );
  INV_X1 U558 ( .A(G469), .ZN(n508) );
  XNOR2_X1 U559 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U560 ( .A(n470), .B(n450), .ZN(n471) );
  INV_X1 U561 ( .A(KEYINPUT83), .ZN(n537) );
  INV_X1 U562 ( .A(n552), .ZN(n581) );
  XNOR2_X1 U563 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n462) );
  XNOR2_X2 U564 ( .A(G146), .B(G125), .ZN(n463) );
  XNOR2_X1 U565 ( .A(n457), .B(n456), .ZN(n460) );
  XNOR2_X1 U566 ( .A(n715), .B(n460), .ZN(n533) );
  XNOR2_X1 U567 ( .A(n533), .B(KEYINPUT117), .ZN(n461) );
  XNOR2_X1 U568 ( .A(KEYINPUT13), .B(G475), .ZN(n474) );
  NAND2_X1 U569 ( .A1(G214), .A2(n516), .ZN(n464) );
  XNOR2_X1 U570 ( .A(KEYINPUT10), .B(n463), .ZN(n490) );
  XNOR2_X1 U571 ( .A(n464), .B(n490), .ZN(n465) );
  XNOR2_X1 U572 ( .A(G143), .B(n506), .ZN(n466) );
  XNOR2_X1 U573 ( .A(n467), .B(KEYINPUT96), .ZN(n470) );
  XOR2_X1 U574 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n469) );
  XNOR2_X1 U575 ( .A(G140), .B(KEYINPUT97), .ZN(n468) );
  NOR2_X1 U576 ( .A1(G902), .A2(n701), .ZN(n473) );
  INV_X1 U577 ( .A(n564), .ZN(n547) );
  XNOR2_X1 U578 ( .A(n475), .B(KEYINPUT7), .ZN(n483) );
  NAND2_X1 U579 ( .A1(G234), .A2(n710), .ZN(n476) );
  XNOR2_X1 U580 ( .A(n477), .B(n476), .ZN(n491) );
  NAND2_X1 U581 ( .A1(G217), .A2(n491), .ZN(n481) );
  XNOR2_X1 U582 ( .A(KEYINPUT9), .B(KEYINPUT98), .ZN(n480) );
  INV_X1 U583 ( .A(n478), .ZN(n479) );
  XNOR2_X1 U584 ( .A(n483), .B(n482), .ZN(n624) );
  XOR2_X1 U585 ( .A(n484), .B(G478), .Z(n565) );
  NAND2_X1 U586 ( .A1(n547), .A2(n565), .ZN(n644) );
  XOR2_X1 U587 ( .A(KEYINPUT91), .B(KEYINPUT81), .Z(n486) );
  XNOR2_X1 U588 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U589 ( .A(n487), .B(KEYINPUT23), .Z(n489) );
  XNOR2_X1 U590 ( .A(G119), .B(G128), .ZN(n488) );
  XNOR2_X1 U591 ( .A(n489), .B(n488), .ZN(n493) );
  XNOR2_X1 U592 ( .A(n490), .B(n500), .ZN(n721) );
  XNOR2_X1 U593 ( .A(n721), .B(n453), .ZN(n492) );
  XNOR2_X1 U594 ( .A(n492), .B(n493), .ZN(n703) );
  XOR2_X1 U595 ( .A(KEYINPUT25), .B(KEYINPUT75), .Z(n496) );
  INV_X1 U596 ( .A(n532), .ZN(n620) );
  NAND2_X1 U597 ( .A1(G234), .A2(n620), .ZN(n494) );
  XNOR2_X1 U598 ( .A(KEYINPUT20), .B(n494), .ZN(n497) );
  NAND2_X1 U599 ( .A1(G217), .A2(n497), .ZN(n495) );
  NAND2_X1 U600 ( .A1(G221), .A2(n497), .ZN(n498) );
  XOR2_X1 U601 ( .A(KEYINPUT21), .B(n498), .Z(n662) );
  XOR2_X1 U602 ( .A(n499), .B(n500), .Z(n504) );
  XNOR2_X2 U603 ( .A(n509), .B(n508), .ZN(n557) );
  NAND2_X1 U604 ( .A1(n510), .A2(n557), .ZN(n593) );
  XNOR2_X1 U605 ( .A(KEYINPUT30), .B(KEYINPUT102), .ZN(n524) );
  NAND2_X1 U606 ( .A1(G214), .A2(n534), .ZN(n650) );
  INV_X1 U607 ( .A(KEYINPUT94), .ZN(n522) );
  XOR2_X1 U608 ( .A(KEYINPUT5), .B(KEYINPUT93), .Z(n512) );
  XNOR2_X1 U609 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U610 ( .A(KEYINPUT74), .B(KEYINPUT92), .Z(n518) );
  NAND2_X1 U611 ( .A1(n516), .A2(G210), .ZN(n517) );
  XNOR2_X1 U612 ( .A(n518), .B(n517), .ZN(n519) );
  NAND2_X1 U613 ( .A1(n650), .A2(n671), .ZN(n523) );
  XNOR2_X1 U614 ( .A(n525), .B(KEYINPUT14), .ZN(n526) );
  NAND2_X1 U615 ( .A1(G952), .A2(n526), .ZN(n682) );
  NOR2_X1 U616 ( .A1(G953), .A2(n682), .ZN(n583) );
  NAND2_X1 U617 ( .A1(n526), .A2(G902), .ZN(n527) );
  XOR2_X1 U618 ( .A(KEYINPUT88), .B(n527), .Z(n584) );
  NAND2_X1 U619 ( .A1(G953), .A2(n584), .ZN(n528) );
  NOR2_X1 U620 ( .A1(G900), .A2(n528), .ZN(n529) );
  XOR2_X1 U621 ( .A(KEYINPUT101), .B(n529), .Z(n530) );
  NOR2_X1 U622 ( .A1(n583), .A2(n530), .ZN(n531) );
  XOR2_X1 U623 ( .A(KEYINPUT76), .B(n531), .Z(n542) );
  NOR2_X1 U624 ( .A1(n533), .A2(n532), .ZN(n536) );
  NAND2_X1 U625 ( .A1(G210), .A2(n534), .ZN(n535) );
  XNOR2_X1 U626 ( .A(KEYINPUT38), .B(n581), .ZN(n651) );
  OR2_X1 U627 ( .A1(n644), .A2(n548), .ZN(n540) );
  XNOR2_X1 U628 ( .A(n540), .B(KEYINPUT107), .ZN(n732) );
  XOR2_X1 U629 ( .A(KEYINPUT46), .B(KEYINPUT82), .Z(n551) );
  INV_X1 U630 ( .A(n662), .ZN(n597) );
  NOR2_X1 U631 ( .A1(n597), .A2(n661), .ZN(n541) );
  NAND2_X1 U632 ( .A1(n542), .A2(n541), .ZN(n553) );
  XNOR2_X1 U633 ( .A(KEYINPUT28), .B(n543), .ZN(n544) );
  NAND2_X1 U634 ( .A1(n544), .A2(n557), .ZN(n562) );
  INV_X1 U635 ( .A(n598), .ZN(n654) );
  NAND2_X1 U636 ( .A1(n651), .A2(n650), .ZN(n655) );
  XNOR2_X1 U637 ( .A(KEYINPUT41), .B(KEYINPUT104), .ZN(n545) );
  XNOR2_X1 U638 ( .A(n546), .B(KEYINPUT42), .ZN(n734) );
  NOR2_X1 U639 ( .A1(n547), .A2(n565), .ZN(n637) );
  INV_X1 U640 ( .A(n637), .ZN(n641) );
  NOR2_X1 U641 ( .A1(n641), .A2(n548), .ZN(n549) );
  XNOR2_X1 U642 ( .A(n551), .B(n550), .ZN(n560) );
  NOR2_X1 U643 ( .A1(n641), .A2(n553), .ZN(n554) );
  XOR2_X1 U644 ( .A(n592), .B(KEYINPUT6), .Z(n607) );
  INV_X1 U645 ( .A(n607), .ZN(n612) );
  NAND2_X1 U646 ( .A1(n554), .A2(n612), .ZN(n578) );
  NOR2_X1 U647 ( .A1(n561), .A2(n578), .ZN(n556) );
  XNOR2_X1 U648 ( .A(KEYINPUT36), .B(KEYINPUT85), .ZN(n555) );
  XNOR2_X1 U649 ( .A(n556), .B(n555), .ZN(n558) );
  NOR2_X1 U650 ( .A1(n558), .A2(n665), .ZN(n559) );
  XNOR2_X1 U651 ( .A(n559), .B(KEYINPUT106), .ZN(n739) );
  INV_X1 U652 ( .A(n644), .ZN(n634) );
  INV_X1 U653 ( .A(n656), .ZN(n563) );
  NAND2_X1 U654 ( .A1(n565), .A2(n564), .ZN(n609) );
  NOR2_X1 U655 ( .A1(n581), .A2(n609), .ZN(n567) );
  NAND2_X1 U656 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U657 ( .A(KEYINPUT103), .B(n568), .Z(n735) );
  XNOR2_X1 U658 ( .A(KEYINPUT79), .B(n569), .ZN(n574) );
  XOR2_X1 U659 ( .A(n656), .B(KEYINPUT80), .Z(n594) );
  INV_X1 U660 ( .A(n594), .ZN(n570) );
  NOR2_X1 U661 ( .A1(KEYINPUT47), .A2(n570), .ZN(n571) );
  XNOR2_X1 U662 ( .A(KEYINPUT72), .B(n571), .ZN(n572) );
  NAND2_X1 U663 ( .A1(n572), .A2(n638), .ZN(n573) );
  AND2_X1 U664 ( .A1(n573), .A2(n574), .ZN(n575) );
  INV_X1 U665 ( .A(KEYINPUT48), .ZN(n576) );
  NOR2_X1 U666 ( .A1(n577), .A2(n578), .ZN(n579) );
  NAND2_X1 U667 ( .A1(n579), .A2(n650), .ZN(n580) );
  XNOR2_X1 U668 ( .A(n580), .B(KEYINPUT43), .ZN(n582) );
  NAND2_X1 U669 ( .A1(n582), .A2(n581), .ZN(n647) );
  INV_X1 U670 ( .A(n583), .ZN(n586) );
  NOR2_X1 U671 ( .A1(G898), .A2(n710), .ZN(n717) );
  NAND2_X1 U672 ( .A1(n717), .A2(n584), .ZN(n585) );
  NAND2_X1 U673 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U674 ( .A(KEYINPUT89), .B(n587), .ZN(n588) );
  NOR2_X1 U675 ( .A1(n592), .A2(n605), .ZN(n673) );
  NAND2_X1 U676 ( .A1(n596), .A2(n673), .ZN(n591) );
  XOR2_X1 U677 ( .A(KEYINPUT31), .B(n591), .Z(n643) );
  NAND2_X1 U678 ( .A1(n643), .A2(n629), .ZN(n595) );
  NAND2_X1 U679 ( .A1(n595), .A2(n594), .ZN(n603) );
  XNOR2_X1 U680 ( .A(n600), .B(n599), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n665), .A2(n607), .ZN(n601) );
  NOR2_X1 U682 ( .A1(n611), .A2(n601), .ZN(n602) );
  NAND2_X1 U683 ( .A1(n602), .A2(n378), .ZN(n626) );
  NAND2_X1 U684 ( .A1(n603), .A2(n626), .ZN(n604) );
  XNOR2_X1 U685 ( .A(n605), .B(KEYINPUT100), .ZN(n606) );
  INV_X1 U686 ( .A(KEYINPUT35), .ZN(n610) );
  NOR2_X1 U687 ( .A1(n611), .A2(n378), .ZN(n616) );
  NOR2_X1 U688 ( .A1(n612), .A2(n665), .ZN(n613) );
  NOR2_X1 U689 ( .A1(n671), .A2(n577), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n616), .A2(n615), .ZN(n633) );
  NAND2_X1 U691 ( .A1(n741), .A2(n633), .ZN(n618) );
  NAND2_X1 U692 ( .A1(n618), .A2(KEYINPUT44), .ZN(n617) );
  INV_X1 U693 ( .A(KEYINPUT2), .ZN(n619) );
  NAND2_X1 U694 ( .A1(n704), .A2(G210), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n704), .A2(G472), .ZN(n623) );
  NAND2_X1 U696 ( .A1(n704), .A2(G478), .ZN(n625) );
  XNOR2_X1 U697 ( .A(G101), .B(n626), .ZN(G3) );
  NOR2_X1 U698 ( .A1(n641), .A2(n629), .ZN(n627) );
  XOR2_X1 U699 ( .A(KEYINPUT108), .B(n627), .Z(n628) );
  XNOR2_X1 U700 ( .A(G104), .B(n628), .ZN(G6) );
  NOR2_X1 U701 ( .A1(n644), .A2(n629), .ZN(n631) );
  XNOR2_X1 U702 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n630) );
  XNOR2_X1 U703 ( .A(n631), .B(n630), .ZN(n632) );
  XNOR2_X1 U704 ( .A(G107), .B(n632), .ZN(G9) );
  XNOR2_X1 U705 ( .A(G110), .B(n633), .ZN(G12) );
  XOR2_X1 U706 ( .A(G128), .B(KEYINPUT29), .Z(n636) );
  NAND2_X1 U707 ( .A1(n638), .A2(n634), .ZN(n635) );
  XNOR2_X1 U708 ( .A(n636), .B(n635), .ZN(G30) );
  XOR2_X1 U709 ( .A(G146), .B(KEYINPUT109), .Z(n640) );
  NAND2_X1 U710 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U711 ( .A(n640), .B(n639), .ZN(G48) );
  NOR2_X1 U712 ( .A1(n641), .A2(n643), .ZN(n642) );
  XOR2_X1 U713 ( .A(G113), .B(n642), .Z(G15) );
  NOR2_X1 U714 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U715 ( .A(KEYINPUT110), .B(n645), .Z(n646) );
  XNOR2_X1 U716 ( .A(G116), .B(n646), .ZN(G18) );
  XNOR2_X1 U717 ( .A(G140), .B(n647), .ZN(G42) );
  INV_X1 U718 ( .A(n648), .ZN(n660) );
  NOR2_X1 U719 ( .A1(n676), .A2(n660), .ZN(n649) );
  XOR2_X1 U720 ( .A(KEYINPUT115), .B(n649), .Z(n685) );
  NOR2_X1 U721 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U722 ( .A(KEYINPUT113), .B(n652), .Z(n653) );
  NOR2_X1 U723 ( .A1(n654), .A2(n653), .ZN(n658) );
  NOR2_X1 U724 ( .A1(n656), .A2(n655), .ZN(n657) );
  NOR2_X1 U725 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U726 ( .A1(n660), .A2(n659), .ZN(n679) );
  NOR2_X1 U727 ( .A1(n662), .A2(n378), .ZN(n663) );
  XNOR2_X1 U728 ( .A(KEYINPUT49), .B(n663), .ZN(n669) );
  XOR2_X1 U729 ( .A(KEYINPUT50), .B(KEYINPUT111), .Z(n667) );
  NAND2_X1 U730 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U731 ( .A(n667), .B(n666), .ZN(n668) );
  NAND2_X1 U732 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U733 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U734 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U735 ( .A(KEYINPUT51), .B(n674), .Z(n675) );
  NOR2_X1 U736 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U737 ( .A(n677), .B(KEYINPUT112), .ZN(n678) );
  NOR2_X1 U738 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U739 ( .A(n680), .B(KEYINPUT52), .ZN(n681) );
  NOR2_X1 U740 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U741 ( .A(KEYINPUT114), .B(n683), .ZN(n684) );
  NOR2_X1 U742 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U743 ( .A(n686), .B(KEYINPUT116), .ZN(n687) );
  NAND2_X1 U744 ( .A1(n687), .A2(n710), .ZN(n695) );
  XOR2_X1 U745 ( .A(KEYINPUT2), .B(KEYINPUT78), .Z(n689) );
  NAND2_X1 U746 ( .A1(n689), .A2(n691), .ZN(n690) );
  XNOR2_X1 U747 ( .A(n690), .B(KEYINPUT77), .ZN(n693) );
  NOR2_X1 U748 ( .A1(n691), .A2(n619), .ZN(n692) );
  NOR2_X1 U749 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U750 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U751 ( .A(n696), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U752 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n698) );
  NAND2_X1 U753 ( .A1(n704), .A2(G469), .ZN(n697) );
  NOR2_X1 U754 ( .A1(n708), .A2(n700), .ZN(G54) );
  NAND2_X1 U755 ( .A1(n704), .A2(G475), .ZN(n702) );
  XNOR2_X1 U756 ( .A(n703), .B(KEYINPUT120), .ZN(n706) );
  NAND2_X1 U757 ( .A1(G217), .A2(n704), .ZN(n705) );
  XNOR2_X1 U758 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U759 ( .A1(n708), .A2(n707), .ZN(G66) );
  NAND2_X1 U760 ( .A1(n710), .A2(n709), .ZN(n714) );
  NAND2_X1 U761 ( .A1(G953), .A2(G224), .ZN(n711) );
  XNOR2_X1 U762 ( .A(KEYINPUT61), .B(n711), .ZN(n712) );
  NAND2_X1 U763 ( .A1(n712), .A2(G898), .ZN(n713) );
  NAND2_X1 U764 ( .A1(n714), .A2(n713), .ZN(n719) );
  XNOR2_X1 U765 ( .A(n715), .B(G110), .ZN(n716) );
  NOR2_X1 U766 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U767 ( .A(n719), .B(n718), .ZN(n720) );
  XOR2_X1 U768 ( .A(KEYINPUT121), .B(n720), .Z(G69) );
  XOR2_X1 U769 ( .A(n721), .B(n722), .Z(n725) );
  XNOR2_X1 U770 ( .A(n723), .B(n725), .ZN(n724) );
  NOR2_X1 U771 ( .A1(G953), .A2(n724), .ZN(n730) );
  XNOR2_X1 U772 ( .A(G227), .B(n725), .ZN(n726) );
  NAND2_X1 U773 ( .A1(n726), .A2(G900), .ZN(n727) );
  NAND2_X1 U774 ( .A1(G953), .A2(n727), .ZN(n728) );
  XOR2_X1 U775 ( .A(KEYINPUT122), .B(n728), .Z(n729) );
  NOR2_X1 U776 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U777 ( .A(KEYINPUT123), .B(n731), .ZN(G72) );
  XOR2_X1 U778 ( .A(G134), .B(n732), .Z(G36) );
  XOR2_X1 U779 ( .A(G137), .B(KEYINPUT126), .Z(n733) );
  XNOR2_X1 U780 ( .A(n734), .B(n733), .ZN(G39) );
  XNOR2_X1 U781 ( .A(G143), .B(n735), .ZN(G45) );
  XNOR2_X1 U782 ( .A(G122), .B(KEYINPUT124), .ZN(n738) );
  BUF_X1 U783 ( .A(n736), .Z(n737) );
  XOR2_X1 U784 ( .A(n738), .B(n737), .Z(G24) );
  XNOR2_X1 U785 ( .A(G125), .B(KEYINPUT37), .ZN(n740) );
  XNOR2_X1 U786 ( .A(n740), .B(n739), .ZN(G27) );
  XOR2_X1 U787 ( .A(n741), .B(G119), .Z(n742) );
  XNOR2_X1 U788 ( .A(KEYINPUT125), .B(n742), .ZN(G21) );
  XNOR2_X1 U789 ( .A(G131), .B(KEYINPUT127), .ZN(n743) );
endmodule

