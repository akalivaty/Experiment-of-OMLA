

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U553 ( .A1(n726), .A2(n520), .ZN(n518) );
  XOR2_X1 U554 ( .A(KEYINPUT29), .B(n651), .Z(n519) );
  OR2_X1 U555 ( .A1(n725), .A2(n733), .ZN(n520) );
  NAND2_X1 U556 ( .A1(n737), .A2(n736), .ZN(n521) );
  OR2_X1 U557 ( .A1(KEYINPUT33), .A2(n692), .ZN(n522) );
  NOR2_X1 U558 ( .A1(n607), .A2(n606), .ZN(n608) );
  INV_X1 U559 ( .A(KEYINPUT31), .ZN(n662) );
  AND2_X1 U560 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U561 ( .A1(G2105), .A2(G2104), .ZN(n532) );
  NOR2_X1 U562 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U563 ( .A1(n544), .A2(n525), .ZN(n794) );
  INV_X1 U564 ( .A(G651), .ZN(n525) );
  NOR2_X1 U565 ( .A1(G543), .A2(n525), .ZN(n523) );
  XOR2_X1 U566 ( .A(KEYINPUT1), .B(n523), .Z(n797) );
  AND2_X1 U567 ( .A1(n797), .A2(G60), .ZN(n529) );
  NOR2_X1 U568 ( .A1(G651), .A2(G543), .ZN(n793) );
  NAND2_X1 U569 ( .A1(G85), .A2(n793), .ZN(n527) );
  XNOR2_X1 U570 ( .A(G543), .B(KEYINPUT0), .ZN(n524) );
  XNOR2_X1 U571 ( .A(n524), .B(KEYINPUT67), .ZN(n544) );
  NAND2_X1 U572 ( .A1(G72), .A2(n794), .ZN(n526) );
  NAND2_X1 U573 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U574 ( .A1(n529), .A2(n528), .ZN(n531) );
  NOR2_X2 U575 ( .A1(G651), .A2(n544), .ZN(n798) );
  NAND2_X1 U576 ( .A1(n798), .A2(G47), .ZN(n530) );
  NAND2_X1 U577 ( .A1(n531), .A2(n530), .ZN(G290) );
  XOR2_X2 U578 ( .A(KEYINPUT17), .B(n532), .Z(n874) );
  NAND2_X1 U579 ( .A1(n874), .A2(G138), .ZN(n533) );
  XNOR2_X1 U580 ( .A(n533), .B(KEYINPUT87), .ZN(n542) );
  INV_X1 U581 ( .A(G2104), .ZN(n536) );
  NOR2_X1 U582 ( .A1(G2105), .A2(n536), .ZN(n872) );
  NAND2_X1 U583 ( .A1(G102), .A2(n872), .ZN(n534) );
  XNOR2_X1 U584 ( .A(n534), .B(KEYINPUT86), .ZN(n540) );
  NAND2_X1 U585 ( .A1(G2104), .A2(G2105), .ZN(n535) );
  XNOR2_X1 U586 ( .A(n535), .B(KEYINPUT65), .ZN(n881) );
  NAND2_X1 U587 ( .A1(G114), .A2(n881), .ZN(n538) );
  AND2_X1 U588 ( .A1(n536), .A2(G2105), .ZN(n878) );
  NAND2_X1 U589 ( .A1(G126), .A2(n878), .ZN(n537) );
  AND2_X1 U590 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U591 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X2 U592 ( .A1(n542), .A2(n541), .ZN(G164) );
  NAND2_X1 U593 ( .A1(G74), .A2(G651), .ZN(n543) );
  XNOR2_X1 U594 ( .A(n543), .B(KEYINPUT80), .ZN(n549) );
  NAND2_X1 U595 ( .A1(G49), .A2(n798), .ZN(n546) );
  NAND2_X1 U596 ( .A1(G87), .A2(n544), .ZN(n545) );
  NAND2_X1 U597 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U598 ( .A1(n797), .A2(n547), .ZN(n548) );
  NAND2_X1 U599 ( .A1(n549), .A2(n548), .ZN(G288) );
  NAND2_X1 U600 ( .A1(G64), .A2(n797), .ZN(n551) );
  NAND2_X1 U601 ( .A1(G52), .A2(n798), .ZN(n550) );
  NAND2_X1 U602 ( .A1(n551), .A2(n550), .ZN(n557) );
  NAND2_X1 U603 ( .A1(G90), .A2(n793), .ZN(n553) );
  NAND2_X1 U604 ( .A1(G77), .A2(n794), .ZN(n552) );
  NAND2_X1 U605 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U606 ( .A(KEYINPUT9), .B(n554), .Z(n555) );
  XNOR2_X1 U607 ( .A(KEYINPUT68), .B(n555), .ZN(n556) );
  NOR2_X1 U608 ( .A1(n557), .A2(n556), .ZN(G171) );
  NAND2_X1 U609 ( .A1(G78), .A2(n794), .ZN(n558) );
  XNOR2_X1 U610 ( .A(n558), .B(KEYINPUT70), .ZN(n561) );
  NAND2_X1 U611 ( .A1(G91), .A2(n793), .ZN(n559) );
  XOR2_X1 U612 ( .A(KEYINPUT69), .B(n559), .Z(n560) );
  NAND2_X1 U613 ( .A1(n561), .A2(n560), .ZN(n564) );
  NAND2_X1 U614 ( .A1(G65), .A2(n797), .ZN(n562) );
  XNOR2_X1 U615 ( .A(KEYINPUT71), .B(n562), .ZN(n563) );
  NOR2_X1 U616 ( .A1(n564), .A2(n563), .ZN(n566) );
  NAND2_X1 U617 ( .A1(n798), .A2(G53), .ZN(n565) );
  NAND2_X1 U618 ( .A1(n566), .A2(n565), .ZN(G299) );
  NAND2_X1 U619 ( .A1(n793), .A2(G89), .ZN(n567) );
  XNOR2_X1 U620 ( .A(n567), .B(KEYINPUT4), .ZN(n569) );
  NAND2_X1 U621 ( .A1(G76), .A2(n794), .ZN(n568) );
  NAND2_X1 U622 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U623 ( .A(n570), .B(KEYINPUT5), .ZN(n576) );
  XNOR2_X1 U624 ( .A(KEYINPUT6), .B(KEYINPUT75), .ZN(n574) );
  NAND2_X1 U625 ( .A1(G63), .A2(n797), .ZN(n572) );
  NAND2_X1 U626 ( .A1(G51), .A2(n798), .ZN(n571) );
  NAND2_X1 U627 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U628 ( .A(n574), .B(n573), .ZN(n575) );
  NAND2_X1 U629 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U630 ( .A(KEYINPUT7), .B(n577), .ZN(G168) );
  XOR2_X1 U631 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U632 ( .A1(G88), .A2(n793), .ZN(n579) );
  NAND2_X1 U633 ( .A1(G75), .A2(n794), .ZN(n578) );
  NAND2_X1 U634 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U635 ( .A1(G62), .A2(n797), .ZN(n581) );
  NAND2_X1 U636 ( .A1(G50), .A2(n798), .ZN(n580) );
  NAND2_X1 U637 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U638 ( .A1(n583), .A2(n582), .ZN(G166) );
  INV_X1 U639 ( .A(G166), .ZN(G303) );
  XOR2_X1 U640 ( .A(KEYINPUT2), .B(KEYINPUT81), .Z(n585) );
  NAND2_X1 U641 ( .A1(G73), .A2(n794), .ZN(n584) );
  XNOR2_X1 U642 ( .A(n585), .B(n584), .ZN(n592) );
  NAND2_X1 U643 ( .A1(G86), .A2(n793), .ZN(n587) );
  NAND2_X1 U644 ( .A1(G61), .A2(n797), .ZN(n586) );
  NAND2_X1 U645 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U646 ( .A1(n798), .A2(G48), .ZN(n588) );
  XOR2_X1 U647 ( .A(KEYINPUT82), .B(n588), .Z(n589) );
  NOR2_X1 U648 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U649 ( .A1(n592), .A2(n591), .ZN(G305) );
  XNOR2_X1 U650 ( .A(G1986), .B(G290), .ZN(n966) );
  NOR2_X1 U651 ( .A1(G164), .A2(G1384), .ZN(n603) );
  NAND2_X1 U652 ( .A1(G137), .A2(n874), .ZN(n593) );
  XNOR2_X1 U653 ( .A(n593), .B(KEYINPUT66), .ZN(n596) );
  NAND2_X1 U654 ( .A1(G101), .A2(n872), .ZN(n594) );
  XOR2_X1 U655 ( .A(KEYINPUT23), .B(n594), .Z(n595) );
  NAND2_X1 U656 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U657 ( .A1(G113), .A2(n881), .ZN(n598) );
  NAND2_X1 U658 ( .A1(G125), .A2(n878), .ZN(n597) );
  NAND2_X1 U659 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U660 ( .A1(n600), .A2(n599), .ZN(n777) );
  AND2_X1 U661 ( .A1(n777), .A2(G40), .ZN(n602) );
  INV_X1 U662 ( .A(n602), .ZN(n601) );
  NOR2_X1 U663 ( .A1(n603), .A2(n601), .ZN(n752) );
  NAND2_X1 U664 ( .A1(n966), .A2(n752), .ZN(n740) );
  NAND2_X1 U665 ( .A1(n603), .A2(n602), .ZN(n668) );
  NAND2_X1 U666 ( .A1(G8), .A2(n668), .ZN(n733) );
  NAND2_X1 U667 ( .A1(G1976), .A2(G288), .ZN(n973) );
  INV_X1 U668 ( .A(n668), .ZN(n623) );
  XNOR2_X1 U669 ( .A(G2078), .B(KEYINPUT96), .ZN(n604) );
  XNOR2_X1 U670 ( .A(n604), .B(KEYINPUT25), .ZN(n952) );
  NAND2_X1 U671 ( .A1(n623), .A2(n952), .ZN(n605) );
  XNOR2_X1 U672 ( .A(n605), .B(KEYINPUT97), .ZN(n607) );
  INV_X1 U673 ( .A(n668), .ZN(n637) );
  NOR2_X1 U674 ( .A1(n637), .A2(G1961), .ZN(n606) );
  XOR2_X1 U675 ( .A(KEYINPUT98), .B(n608), .Z(n659) );
  NAND2_X1 U676 ( .A1(G171), .A2(n659), .ZN(n652) );
  INV_X1 U677 ( .A(G299), .ZN(n975) );
  NAND2_X1 U678 ( .A1(n637), .A2(G2072), .ZN(n609) );
  XNOR2_X1 U679 ( .A(n609), .B(KEYINPUT27), .ZN(n611) );
  INV_X1 U680 ( .A(G1956), .ZN(n991) );
  NOR2_X1 U681 ( .A1(n991), .A2(n637), .ZN(n610) );
  NOR2_X1 U682 ( .A1(n611), .A2(n610), .ZN(n614) );
  NOR2_X1 U683 ( .A1(n975), .A2(n614), .ZN(n613) );
  XNOR2_X1 U684 ( .A(KEYINPUT99), .B(KEYINPUT28), .ZN(n612) );
  XNOR2_X1 U685 ( .A(n613), .B(n612), .ZN(n650) );
  NAND2_X1 U686 ( .A1(n975), .A2(n614), .ZN(n648) );
  NAND2_X1 U687 ( .A1(G79), .A2(n794), .ZN(n616) );
  NAND2_X1 U688 ( .A1(G54), .A2(n798), .ZN(n615) );
  NAND2_X1 U689 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U690 ( .A(KEYINPUT74), .B(n617), .ZN(n621) );
  NAND2_X1 U691 ( .A1(G92), .A2(n793), .ZN(n619) );
  NAND2_X1 U692 ( .A1(G66), .A2(n797), .ZN(n618) );
  NAND2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U694 ( .A(KEYINPUT15), .B(n622), .Z(n969) );
  NAND2_X1 U695 ( .A1(G2067), .A2(n623), .ZN(n625) );
  NAND2_X1 U696 ( .A1(G1348), .A2(n668), .ZN(n624) );
  NAND2_X1 U697 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U698 ( .A(KEYINPUT101), .B(n626), .ZN(n644) );
  OR2_X1 U699 ( .A1(n969), .A2(n644), .ZN(n643) );
  NAND2_X1 U700 ( .A1(n793), .A2(G81), .ZN(n627) );
  XNOR2_X1 U701 ( .A(n627), .B(KEYINPUT12), .ZN(n629) );
  NAND2_X1 U702 ( .A1(G68), .A2(n794), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U704 ( .A(KEYINPUT13), .B(n630), .Z(n634) );
  NAND2_X1 U705 ( .A1(G56), .A2(n797), .ZN(n631) );
  XNOR2_X1 U706 ( .A(n631), .B(KEYINPUT14), .ZN(n632) );
  XNOR2_X1 U707 ( .A(n632), .B(KEYINPUT73), .ZN(n633) );
  NOR2_X1 U708 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U709 ( .A1(n798), .A2(G43), .ZN(n635) );
  NAND2_X1 U710 ( .A1(n636), .A2(n635), .ZN(n964) );
  XNOR2_X1 U711 ( .A(G1996), .B(KEYINPUT100), .ZN(n946) );
  NAND2_X1 U712 ( .A1(n946), .A2(n637), .ZN(n638) );
  XNOR2_X1 U713 ( .A(n638), .B(KEYINPUT26), .ZN(n640) );
  NAND2_X1 U714 ( .A1(n668), .A2(G1341), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U716 ( .A1(n964), .A2(n641), .ZN(n642) );
  NAND2_X1 U717 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U718 ( .A1(n644), .A2(n969), .ZN(n645) );
  AND2_X1 U719 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U720 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U721 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U722 ( .A1(n652), .A2(n519), .ZN(n665) );
  INV_X1 U723 ( .A(G8), .ZN(n655) );
  NOR2_X1 U724 ( .A1(n655), .A2(G1966), .ZN(n653) );
  AND2_X1 U725 ( .A1(n653), .A2(n668), .ZN(n654) );
  XNOR2_X1 U726 ( .A(n654), .B(KEYINPUT95), .ZN(n680) );
  NOR2_X1 U727 ( .A1(G2084), .A2(n668), .ZN(n676) );
  NOR2_X1 U728 ( .A1(n655), .A2(n676), .ZN(n656) );
  AND2_X1 U729 ( .A1(n680), .A2(n656), .ZN(n657) );
  XOR2_X1 U730 ( .A(KEYINPUT30), .B(n657), .Z(n658) );
  NOR2_X1 U731 ( .A1(G168), .A2(n658), .ZN(n661) );
  NOR2_X1 U732 ( .A1(G171), .A2(n659), .ZN(n660) );
  NOR2_X1 U733 ( .A1(n661), .A2(n660), .ZN(n663) );
  XNOR2_X1 U734 ( .A(n663), .B(n662), .ZN(n664) );
  NAND2_X1 U735 ( .A1(n665), .A2(n664), .ZN(n679) );
  AND2_X1 U736 ( .A1(G286), .A2(G8), .ZN(n666) );
  NAND2_X1 U737 ( .A1(n679), .A2(n666), .ZN(n674) );
  NOR2_X1 U738 ( .A1(G1971), .A2(n733), .ZN(n667) );
  XOR2_X1 U739 ( .A(KEYINPUT103), .B(n667), .Z(n670) );
  NOR2_X1 U740 ( .A1(G2090), .A2(n668), .ZN(n669) );
  NOR2_X1 U741 ( .A1(n670), .A2(n669), .ZN(n671) );
  NAND2_X1 U742 ( .A1(n671), .A2(G303), .ZN(n672) );
  OR2_X1 U743 ( .A1(n655), .A2(n672), .ZN(n673) );
  XNOR2_X1 U744 ( .A(n675), .B(KEYINPUT32), .ZN(n686) );
  NAND2_X1 U745 ( .A1(n676), .A2(G8), .ZN(n677) );
  XNOR2_X1 U746 ( .A(n677), .B(KEYINPUT94), .ZN(n684) );
  INV_X1 U747 ( .A(KEYINPUT102), .ZN(n678) );
  XNOR2_X1 U748 ( .A(n679), .B(n678), .ZN(n682) );
  INV_X1 U749 ( .A(n680), .ZN(n681) );
  NOR2_X1 U750 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U751 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U752 ( .A1(n686), .A2(n685), .ZN(n729) );
  NOR2_X1 U753 ( .A1(G1976), .A2(G288), .ZN(n724) );
  NOR2_X1 U754 ( .A1(G1971), .A2(G303), .ZN(n687) );
  NOR2_X1 U755 ( .A1(n724), .A2(n687), .ZN(n974) );
  NAND2_X1 U756 ( .A1(n729), .A2(n974), .ZN(n688) );
  NAND2_X1 U757 ( .A1(n973), .A2(n688), .ZN(n689) );
  XNOR2_X1 U758 ( .A(KEYINPUT104), .B(n689), .ZN(n690) );
  NOR2_X1 U759 ( .A1(n733), .A2(n690), .ZN(n691) );
  XNOR2_X1 U760 ( .A(n691), .B(KEYINPUT64), .ZN(n692) );
  XOR2_X1 U761 ( .A(G1981), .B(G305), .Z(n981) );
  XNOR2_X1 U762 ( .A(G2067), .B(KEYINPUT37), .ZN(n693) );
  XNOR2_X1 U763 ( .A(n693), .B(KEYINPUT88), .ZN(n749) );
  NAND2_X1 U764 ( .A1(n872), .A2(G104), .ZN(n694) );
  XOR2_X1 U765 ( .A(KEYINPUT89), .B(n694), .Z(n696) );
  NAND2_X1 U766 ( .A1(n874), .A2(G140), .ZN(n695) );
  NAND2_X1 U767 ( .A1(n696), .A2(n695), .ZN(n698) );
  XNOR2_X1 U768 ( .A(KEYINPUT34), .B(KEYINPUT90), .ZN(n697) );
  XNOR2_X1 U769 ( .A(n698), .B(n697), .ZN(n703) );
  NAND2_X1 U770 ( .A1(G116), .A2(n881), .ZN(n700) );
  NAND2_X1 U771 ( .A1(G128), .A2(n878), .ZN(n699) );
  NAND2_X1 U772 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U773 ( .A(KEYINPUT35), .B(n701), .Z(n702) );
  NOR2_X1 U774 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U775 ( .A(KEYINPUT36), .B(n704), .ZN(n899) );
  NOR2_X1 U776 ( .A1(n749), .A2(n899), .ZN(n924) );
  NAND2_X1 U777 ( .A1(n752), .A2(n924), .ZN(n747) );
  NAND2_X1 U778 ( .A1(G119), .A2(n878), .ZN(n711) );
  NAND2_X1 U779 ( .A1(G131), .A2(n874), .ZN(n706) );
  NAND2_X1 U780 ( .A1(G107), .A2(n881), .ZN(n705) );
  NAND2_X1 U781 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U782 ( .A1(G95), .A2(n872), .ZN(n707) );
  XNOR2_X1 U783 ( .A(KEYINPUT91), .B(n707), .ZN(n708) );
  NOR2_X1 U784 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U785 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U786 ( .A(n712), .B(KEYINPUT92), .ZN(n886) );
  NAND2_X1 U787 ( .A1(G1991), .A2(n886), .ZN(n721) );
  NAND2_X1 U788 ( .A1(G117), .A2(n881), .ZN(n714) );
  NAND2_X1 U789 ( .A1(G129), .A2(n878), .ZN(n713) );
  NAND2_X1 U790 ( .A1(n714), .A2(n713), .ZN(n717) );
  NAND2_X1 U791 ( .A1(n872), .A2(G105), .ZN(n715) );
  XOR2_X1 U792 ( .A(KEYINPUT38), .B(n715), .Z(n716) );
  NOR2_X1 U793 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U794 ( .A1(n874), .A2(G141), .ZN(n718) );
  NAND2_X1 U795 ( .A1(n719), .A2(n718), .ZN(n887) );
  NAND2_X1 U796 ( .A1(G1996), .A2(n887), .ZN(n720) );
  NAND2_X1 U797 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U798 ( .A(KEYINPUT93), .B(n722), .ZN(n929) );
  INV_X1 U799 ( .A(n929), .ZN(n723) );
  NAND2_X1 U800 ( .A1(n723), .A2(n752), .ZN(n741) );
  AND2_X1 U801 ( .A1(n747), .A2(n741), .ZN(n737) );
  AND2_X1 U802 ( .A1(n981), .A2(n737), .ZN(n726) );
  NAND2_X1 U803 ( .A1(n724), .A2(KEYINPUT33), .ZN(n725) );
  NAND2_X1 U804 ( .A1(n522), .A2(n518), .ZN(n738) );
  NOR2_X1 U805 ( .A1(G2090), .A2(G303), .ZN(n727) );
  NAND2_X1 U806 ( .A1(G8), .A2(n727), .ZN(n728) );
  NAND2_X1 U807 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U808 ( .A1(n730), .A2(n733), .ZN(n735) );
  NOR2_X1 U809 ( .A1(G1981), .A2(G305), .ZN(n731) );
  XOR2_X1 U810 ( .A(n731), .B(KEYINPUT24), .Z(n732) );
  OR2_X1 U811 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U812 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U813 ( .A1(n738), .A2(n521), .ZN(n739) );
  NAND2_X1 U814 ( .A1(n740), .A2(n739), .ZN(n755) );
  NOR2_X1 U815 ( .A1(G1996), .A2(n887), .ZN(n915) );
  INV_X1 U816 ( .A(n741), .ZN(n744) );
  NOR2_X1 U817 ( .A1(G1991), .A2(n886), .ZN(n920) );
  NOR2_X1 U818 ( .A1(G1986), .A2(G290), .ZN(n742) );
  NOR2_X1 U819 ( .A1(n920), .A2(n742), .ZN(n743) );
  NOR2_X1 U820 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U821 ( .A1(n915), .A2(n745), .ZN(n746) );
  XNOR2_X1 U822 ( .A(n746), .B(KEYINPUT39), .ZN(n748) );
  NAND2_X1 U823 ( .A1(n748), .A2(n747), .ZN(n750) );
  NAND2_X1 U824 ( .A1(n749), .A2(n899), .ZN(n917) );
  NAND2_X1 U825 ( .A1(n750), .A2(n917), .ZN(n751) );
  XOR2_X1 U826 ( .A(KEYINPUT105), .B(n751), .Z(n753) );
  NAND2_X1 U827 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U828 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U829 ( .A(n756), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U830 ( .A(G2443), .B(G2446), .Z(n758) );
  XNOR2_X1 U831 ( .A(G2427), .B(G2451), .ZN(n757) );
  XNOR2_X1 U832 ( .A(n758), .B(n757), .ZN(n764) );
  XOR2_X1 U833 ( .A(G2430), .B(G2454), .Z(n760) );
  XNOR2_X1 U834 ( .A(G1341), .B(G1348), .ZN(n759) );
  XNOR2_X1 U835 ( .A(n760), .B(n759), .ZN(n762) );
  XOR2_X1 U836 ( .A(G2435), .B(G2438), .Z(n761) );
  XNOR2_X1 U837 ( .A(n762), .B(n761), .ZN(n763) );
  XOR2_X1 U838 ( .A(n764), .B(n763), .Z(n765) );
  AND2_X1 U839 ( .A1(G14), .A2(n765), .ZN(G401) );
  AND2_X1 U840 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U841 ( .A1(G111), .A2(n881), .ZN(n774) );
  NAND2_X1 U842 ( .A1(G123), .A2(n878), .ZN(n766) );
  XNOR2_X1 U843 ( .A(n766), .B(KEYINPUT76), .ZN(n767) );
  XNOR2_X1 U844 ( .A(n767), .B(KEYINPUT18), .ZN(n769) );
  NAND2_X1 U845 ( .A1(G135), .A2(n874), .ZN(n768) );
  NAND2_X1 U846 ( .A1(n769), .A2(n768), .ZN(n772) );
  NAND2_X1 U847 ( .A1(G99), .A2(n872), .ZN(n770) );
  XNOR2_X1 U848 ( .A(KEYINPUT77), .B(n770), .ZN(n771) );
  NOR2_X1 U849 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U850 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U851 ( .A(n775), .B(KEYINPUT78), .ZN(n922) );
  XNOR2_X1 U852 ( .A(n922), .B(G2096), .ZN(n776) );
  OR2_X1 U853 ( .A1(G2100), .A2(n776), .ZN(G156) );
  BUF_X1 U854 ( .A(n777), .Z(G160) );
  INV_X1 U855 ( .A(G57), .ZN(G237) );
  INV_X1 U856 ( .A(G132), .ZN(G219) );
  INV_X1 U857 ( .A(G82), .ZN(G220) );
  INV_X1 U858 ( .A(G96), .ZN(G221) );
  NAND2_X1 U859 ( .A1(G7), .A2(G661), .ZN(n778) );
  XNOR2_X1 U860 ( .A(n778), .B(KEYINPUT72), .ZN(n779) );
  XNOR2_X1 U861 ( .A(KEYINPUT10), .B(n779), .ZN(G223) );
  INV_X1 U862 ( .A(G223), .ZN(n830) );
  NAND2_X1 U863 ( .A1(n830), .A2(G567), .ZN(n780) );
  XOR2_X1 U864 ( .A(KEYINPUT11), .B(n780), .Z(G234) );
  INV_X1 U865 ( .A(G860), .ZN(n792) );
  OR2_X1 U866 ( .A1(n964), .A2(n792), .ZN(G153) );
  INV_X1 U867 ( .A(G171), .ZN(G301) );
  NAND2_X1 U868 ( .A1(G868), .A2(G301), .ZN(n782) );
  OR2_X1 U869 ( .A1(n969), .A2(G868), .ZN(n781) );
  NAND2_X1 U870 ( .A1(n782), .A2(n781), .ZN(G284) );
  INV_X1 U871 ( .A(G868), .ZN(n783) );
  NOR2_X1 U872 ( .A1(G286), .A2(n783), .ZN(n785) );
  NOR2_X1 U873 ( .A1(G868), .A2(G299), .ZN(n784) );
  NOR2_X1 U874 ( .A1(n785), .A2(n784), .ZN(G297) );
  NAND2_X1 U875 ( .A1(n792), .A2(G559), .ZN(n786) );
  NAND2_X1 U876 ( .A1(n786), .A2(n969), .ZN(n787) );
  XNOR2_X1 U877 ( .A(n787), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U878 ( .A1(G868), .A2(n964), .ZN(n790) );
  NAND2_X1 U879 ( .A1(G868), .A2(n969), .ZN(n788) );
  NOR2_X1 U880 ( .A1(G559), .A2(n788), .ZN(n789) );
  NOR2_X1 U881 ( .A1(n790), .A2(n789), .ZN(G282) );
  NAND2_X1 U882 ( .A1(G559), .A2(n969), .ZN(n791) );
  XOR2_X1 U883 ( .A(n964), .B(n791), .Z(n811) );
  NAND2_X1 U884 ( .A1(n792), .A2(n811), .ZN(n804) );
  NAND2_X1 U885 ( .A1(G93), .A2(n793), .ZN(n796) );
  NAND2_X1 U886 ( .A1(G80), .A2(n794), .ZN(n795) );
  NAND2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n803) );
  NAND2_X1 U888 ( .A1(G67), .A2(n797), .ZN(n800) );
  NAND2_X1 U889 ( .A1(G55), .A2(n798), .ZN(n799) );
  NAND2_X1 U890 ( .A1(n800), .A2(n799), .ZN(n801) );
  XOR2_X1 U891 ( .A(KEYINPUT79), .B(n801), .Z(n802) );
  NOR2_X1 U892 ( .A1(n803), .A2(n802), .ZN(n813) );
  XOR2_X1 U893 ( .A(n804), .B(n813), .Z(G145) );
  XOR2_X1 U894 ( .A(KEYINPUT83), .B(KEYINPUT19), .Z(n805) );
  XNOR2_X1 U895 ( .A(G288), .B(n805), .ZN(n806) );
  XNOR2_X1 U896 ( .A(G166), .B(n806), .ZN(n808) );
  XNOR2_X1 U897 ( .A(G290), .B(n975), .ZN(n807) );
  XNOR2_X1 U898 ( .A(n808), .B(n807), .ZN(n809) );
  XOR2_X1 U899 ( .A(n813), .B(n809), .Z(n810) );
  XNOR2_X1 U900 ( .A(G305), .B(n810), .ZN(n902) );
  XNOR2_X1 U901 ( .A(n811), .B(n902), .ZN(n812) );
  NAND2_X1 U902 ( .A1(n812), .A2(G868), .ZN(n815) );
  OR2_X1 U903 ( .A1(G868), .A2(n813), .ZN(n814) );
  NAND2_X1 U904 ( .A1(n815), .A2(n814), .ZN(G295) );
  NAND2_X1 U905 ( .A1(G2084), .A2(G2078), .ZN(n816) );
  XOR2_X1 U906 ( .A(KEYINPUT20), .B(n816), .Z(n817) );
  NAND2_X1 U907 ( .A1(G2090), .A2(n817), .ZN(n818) );
  XNOR2_X1 U908 ( .A(KEYINPUT21), .B(n818), .ZN(n819) );
  NAND2_X1 U909 ( .A1(n819), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U910 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U911 ( .A1(G220), .A2(G219), .ZN(n820) );
  XOR2_X1 U912 ( .A(KEYINPUT22), .B(n820), .Z(n821) );
  NOR2_X1 U913 ( .A1(G218), .A2(n821), .ZN(n822) );
  XOR2_X1 U914 ( .A(KEYINPUT84), .B(n822), .Z(n823) );
  NOR2_X1 U915 ( .A1(G221), .A2(n823), .ZN(n824) );
  XNOR2_X1 U916 ( .A(KEYINPUT85), .B(n824), .ZN(n835) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n835), .ZN(n828) );
  NAND2_X1 U918 ( .A1(G69), .A2(G120), .ZN(n825) );
  NOR2_X1 U919 ( .A1(G237), .A2(n825), .ZN(n826) );
  NAND2_X1 U920 ( .A1(G108), .A2(n826), .ZN(n834) );
  NAND2_X1 U921 ( .A1(G567), .A2(n834), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n828), .A2(n827), .ZN(n856) );
  NAND2_X1 U923 ( .A1(G661), .A2(G483), .ZN(n829) );
  NOR2_X1 U924 ( .A1(n856), .A2(n829), .ZN(n833) );
  NAND2_X1 U925 ( .A1(n833), .A2(G36), .ZN(G176) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n830), .ZN(G217) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U928 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U930 ( .A1(n833), .A2(n832), .ZN(G188) );
  INV_X1 U932 ( .A(G120), .ZN(G236) );
  INV_X1 U933 ( .A(G69), .ZN(G235) );
  NOR2_X1 U934 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  XOR2_X1 U936 ( .A(KEYINPUT43), .B(KEYINPUT108), .Z(n837) );
  XNOR2_X1 U937 ( .A(KEYINPUT42), .B(G2678), .ZN(n836) );
  XNOR2_X1 U938 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U939 ( .A(KEYINPUT107), .B(G2090), .Z(n839) );
  XNOR2_X1 U940 ( .A(G2067), .B(G2072), .ZN(n838) );
  XNOR2_X1 U941 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U942 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U943 ( .A(G2096), .B(G2100), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n845) );
  XOR2_X1 U945 ( .A(G2084), .B(G2078), .Z(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(G227) );
  XOR2_X1 U947 ( .A(G1976), .B(G1971), .Z(n847) );
  XNOR2_X1 U948 ( .A(G1986), .B(G1956), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U950 ( .A(G1981), .B(G1966), .Z(n849) );
  XNOR2_X1 U951 ( .A(G1996), .B(G1991), .ZN(n848) );
  XNOR2_X1 U952 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U953 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U954 ( .A(KEYINPUT109), .B(G2474), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n855) );
  XOR2_X1 U956 ( .A(G1961), .B(KEYINPUT41), .Z(n854) );
  XNOR2_X1 U957 ( .A(n855), .B(n854), .ZN(G229) );
  XOR2_X1 U958 ( .A(KEYINPUT106), .B(n856), .Z(G319) );
  NAND2_X1 U959 ( .A1(G124), .A2(n878), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n857), .B(KEYINPUT44), .ZN(n859) );
  NAND2_X1 U961 ( .A1(n881), .A2(G112), .ZN(n858) );
  NAND2_X1 U962 ( .A1(n859), .A2(n858), .ZN(n863) );
  NAND2_X1 U963 ( .A1(G100), .A2(n872), .ZN(n861) );
  NAND2_X1 U964 ( .A1(G136), .A2(n874), .ZN(n860) );
  NAND2_X1 U965 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U966 ( .A1(n863), .A2(n862), .ZN(G162) );
  NAND2_X1 U967 ( .A1(G103), .A2(n872), .ZN(n865) );
  NAND2_X1 U968 ( .A1(G139), .A2(n874), .ZN(n864) );
  NAND2_X1 U969 ( .A1(n865), .A2(n864), .ZN(n871) );
  NAND2_X1 U970 ( .A1(n878), .A2(G127), .ZN(n866) );
  XOR2_X1 U971 ( .A(KEYINPUT113), .B(n866), .Z(n868) );
  NAND2_X1 U972 ( .A1(n881), .A2(G115), .ZN(n867) );
  NAND2_X1 U973 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U974 ( .A(KEYINPUT47), .B(n869), .Z(n870) );
  NOR2_X1 U975 ( .A1(n871), .A2(n870), .ZN(n930) );
  NAND2_X1 U976 ( .A1(n872), .A2(G106), .ZN(n873) );
  XOR2_X1 U977 ( .A(KEYINPUT111), .B(n873), .Z(n876) );
  NAND2_X1 U978 ( .A1(n874), .A2(G142), .ZN(n875) );
  NAND2_X1 U979 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U980 ( .A(n877), .B(KEYINPUT45), .ZN(n880) );
  NAND2_X1 U981 ( .A1(G130), .A2(n878), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n884) );
  NAND2_X1 U983 ( .A1(n881), .A2(G118), .ZN(n882) );
  XOR2_X1 U984 ( .A(KEYINPUT110), .B(n882), .Z(n883) );
  NOR2_X1 U985 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U986 ( .A(n930), .B(n885), .ZN(n897) );
  XNOR2_X1 U987 ( .A(n887), .B(n886), .ZN(n889) );
  XNOR2_X1 U988 ( .A(G164), .B(G160), .ZN(n888) );
  XNOR2_X1 U989 ( .A(n889), .B(n888), .ZN(n893) );
  XOR2_X1 U990 ( .A(KEYINPUT114), .B(KEYINPUT112), .Z(n891) );
  XNOR2_X1 U991 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n890) );
  XNOR2_X1 U992 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U993 ( .A(n893), .B(n892), .Z(n895) );
  XNOR2_X1 U994 ( .A(n922), .B(G162), .ZN(n894) );
  XNOR2_X1 U995 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U996 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U997 ( .A(n899), .B(n898), .Z(n900) );
  NOR2_X1 U998 ( .A1(G37), .A2(n900), .ZN(n901) );
  XOR2_X1 U999 ( .A(KEYINPUT115), .B(n901), .Z(G395) );
  XNOR2_X1 U1000 ( .A(n964), .B(n902), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(G171), .B(n969), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(n904), .B(n903), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n905), .B(G286), .ZN(n906) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n906), .ZN(G397) );
  NOR2_X1 U1005 ( .A1(G227), .A2(G229), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n907), .B(KEYINPUT49), .ZN(n911) );
  INV_X1 U1007 ( .A(G319), .ZN(n908) );
  NOR2_X1 U1008 ( .A1(n908), .A2(G401), .ZN(n909) );
  XOR2_X1 U1009 ( .A(KEYINPUT116), .B(n909), .Z(n910) );
  NOR2_X1 U1010 ( .A1(n911), .A2(n910), .ZN(n913) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1012 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1015 ( .A(KEYINPUT55), .B(KEYINPUT118), .ZN(n960) );
  XOR2_X1 U1016 ( .A(G2090), .B(G162), .Z(n914) );
  NOR2_X1 U1017 ( .A1(n915), .A2(n914), .ZN(n916) );
  XOR2_X1 U1018 ( .A(KEYINPUT51), .B(n916), .Z(n918) );
  NAND2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n927) );
  XOR2_X1 U1020 ( .A(G160), .B(G2084), .Z(n919) );
  NOR2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1024 ( .A(KEYINPUT117), .B(n925), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n935) );
  XOR2_X1 U1027 ( .A(G2072), .B(n930), .Z(n932) );
  XOR2_X1 U1028 ( .A(G164), .B(G2078), .Z(n931) );
  NOR2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1030 ( .A(KEYINPUT50), .B(n933), .Z(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1032 ( .A(KEYINPUT52), .B(n936), .Z(n937) );
  NOR2_X1 U1033 ( .A1(n960), .A2(n937), .ZN(n938) );
  XNOR2_X1 U1034 ( .A(KEYINPUT119), .B(n938), .ZN(n939) );
  NAND2_X1 U1035 ( .A1(n939), .A2(G29), .ZN(n1021) );
  XOR2_X1 U1036 ( .A(G2090), .B(G35), .Z(n942) );
  XOR2_X1 U1037 ( .A(G34), .B(KEYINPUT54), .Z(n940) );
  XNOR2_X1 U1038 ( .A(n940), .B(G2084), .ZN(n941) );
  NAND2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n958) );
  XNOR2_X1 U1040 ( .A(G1991), .B(G25), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(G33), .B(G2072), .ZN(n943) );
  NOR2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n951) );
  XOR2_X1 U1043 ( .A(G2067), .B(G26), .Z(n945) );
  NAND2_X1 U1044 ( .A1(n945), .A2(G28), .ZN(n949) );
  XNOR2_X1 U1045 ( .A(G32), .B(n946), .ZN(n947) );
  XNOR2_X1 U1046 ( .A(KEYINPUT120), .B(n947), .ZN(n948) );
  NOR2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n954) );
  XOR2_X1 U1049 ( .A(G27), .B(n952), .Z(n953) );
  NOR2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1051 ( .A(KEYINPUT53), .B(n955), .Z(n956) );
  XNOR2_X1 U1052 ( .A(n956), .B(KEYINPUT121), .ZN(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1054 ( .A(n960), .B(n959), .Z(n961) );
  NOR2_X1 U1055 ( .A1(G29), .A2(n961), .ZN(n962) );
  XOR2_X1 U1056 ( .A(KEYINPUT122), .B(n962), .Z(n963) );
  NAND2_X1 U1057 ( .A1(G11), .A2(n963), .ZN(n1019) );
  XNOR2_X1 U1058 ( .A(G16), .B(KEYINPUT56), .ZN(n990) );
  XNOR2_X1 U1059 ( .A(G171), .B(G1961), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(G1341), .B(n964), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n972) );
  XOR2_X1 U1063 ( .A(G1348), .B(n969), .Z(n970) );
  XNOR2_X1 U1064 ( .A(KEYINPUT124), .B(n970), .ZN(n971) );
  NOR2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n988) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n979) );
  XNOR2_X1 U1067 ( .A(n975), .B(G1956), .ZN(n977) );
  NAND2_X1 U1068 ( .A1(G1971), .A2(G303), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n980) );
  XNOR2_X1 U1071 ( .A(n980), .B(KEYINPUT125), .ZN(n986) );
  XNOR2_X1 U1072 ( .A(G1966), .B(G168), .ZN(n982) );
  NAND2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(n983), .B(KEYINPUT123), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(n984), .B(KEYINPUT57), .ZN(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  NAND2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n1017) );
  INV_X1 U1079 ( .A(G16), .ZN(n1015) );
  XNOR2_X1 U1080 ( .A(G20), .B(n991), .ZN(n995) );
  XNOR2_X1 U1081 ( .A(G1341), .B(G19), .ZN(n993) );
  XNOR2_X1 U1082 ( .A(G1981), .B(G6), .ZN(n992) );
  NOR2_X1 U1083 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n998) );
  XOR2_X1 U1085 ( .A(KEYINPUT59), .B(G1348), .Z(n996) );
  XNOR2_X1 U1086 ( .A(G4), .B(n996), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1088 ( .A(KEYINPUT60), .B(n999), .Z(n1001) );
  XNOR2_X1 U1089 ( .A(G1961), .B(G5), .ZN(n1000) );
  NOR2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1011) );
  XNOR2_X1 U1091 ( .A(G1966), .B(KEYINPUT126), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(n1002), .B(G21), .ZN(n1009) );
  XNOR2_X1 U1093 ( .A(G1971), .B(G22), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(G23), .B(G1976), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XOR2_X1 U1096 ( .A(G1986), .B(G24), .Z(n1005) );
  NAND2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1098 ( .A(KEYINPUT58), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(n1012), .B(KEYINPUT127), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(KEYINPUT61), .B(n1013), .ZN(n1014) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1105 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1022), .Z(G311) );
  INV_X1 U1108 ( .A(G311), .ZN(G150) );
endmodule

