//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1308, new_n1309, new_n1310, new_n1311;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G50), .ZN(new_n204));
  INV_X1    g0004(.A(new_n204), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G77), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(KEYINPUT64), .ZN(new_n209));
  INV_X1    g0009(.A(KEYINPUT64), .ZN(new_n210));
  NAND3_X1  g0010(.A1(new_n210), .A2(G1), .A3(G13), .ZN(new_n211));
  AND2_X1   g0011(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n203), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT0), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n219), .A2(G13), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n220), .B(G250), .C1(G257), .C2(G264), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n217), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G68), .A2(G238), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT65), .Z(new_n228));
  AOI211_X1 g0028(.A(new_n226), .B(new_n228), .C1(G77), .C2(G244), .ZN(new_n229));
  INV_X1    g0029(.A(new_n219), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT1), .Z(new_n232));
  AOI211_X1 g0032(.A(new_n222), .B(new_n232), .C1(new_n218), .C2(new_n221), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n235), .B(new_n236), .Z(new_n237));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND2_X1  g0048(.A1(new_n230), .A2(G33), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n212), .A2(KEYINPUT68), .A3(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  OAI211_X1 g0051(.A(new_n209), .B(new_n211), .C1(new_n251), .C2(new_n219), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT68), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n251), .A2(G20), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n257), .A2(G77), .B1(new_n258), .B2(G50), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(new_n213), .B2(G68), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n256), .A2(new_n260), .ZN(new_n261));
  XOR2_X1   g0061(.A(new_n261), .B(KEYINPUT11), .Z(new_n262));
  NOR2_X1   g0062(.A1(new_n213), .A2(G1), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G13), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G68), .ZN(new_n265));
  OR2_X1    g0065(.A1(new_n265), .A2(KEYINPUT77), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT12), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n267), .B1(new_n265), .B2(KEYINPUT77), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(new_n268), .ZN(new_n270));
  INV_X1    g0070(.A(new_n252), .ZN(new_n271));
  INV_X1    g0071(.A(new_n263), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n269), .B(new_n270), .C1(new_n202), .C2(new_n273), .ZN(new_n274));
  OR2_X1    g0074(.A1(new_n274), .A2(KEYINPUT78), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(KEYINPUT78), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n262), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n279), .A2(new_n280), .A3(G226), .A4(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT73), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT3), .B(G33), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n285), .A2(KEYINPUT73), .A3(G226), .A4(new_n281), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT74), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n279), .A2(new_n280), .A3(G232), .A4(G1698), .ZN(new_n289));
  INV_X1    g0089(.A(G97), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n251), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  AND2_X1   g0092(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  AND3_X1   g0093(.A1(new_n287), .A2(new_n288), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n288), .B1(new_n287), .B2(new_n293), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT67), .ZN(new_n296));
  NAND2_X1  g0096(.A1(G33), .A2(G41), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  AOI211_X1 g0098(.A(new_n296), .B(new_n298), .C1(new_n209), .C2(new_n211), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n209), .A2(new_n211), .ZN(new_n300));
  AOI21_X1  g0100(.A(KEYINPUT67), .B1(new_n300), .B2(new_n297), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n294), .A2(new_n295), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G1), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(G41), .B2(G45), .ZN(new_n305));
  INV_X1    g0105(.A(G274), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n297), .A2(G1), .A3(G13), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n308), .A2(new_n305), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n307), .B1(new_n309), .B2(G238), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT13), .B1(new_n303), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n287), .A2(new_n293), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT74), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n296), .B1(new_n212), .B2(new_n298), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n300), .A2(KEYINPUT67), .A3(new_n297), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n287), .A2(new_n288), .A3(new_n293), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n314), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT13), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n319), .A2(new_n320), .A3(new_n310), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n312), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT75), .B1(new_n322), .B2(G200), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT75), .ZN(new_n324));
  INV_X1    g0124(.A(G200), .ZN(new_n325));
  AOI211_X1 g0125(.A(new_n324), .B(new_n325), .C1(new_n312), .C2(new_n321), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n277), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G190), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n321), .A2(KEYINPUT76), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n320), .B1(new_n319), .B2(new_n310), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n312), .A2(KEYINPUT76), .A3(new_n321), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n328), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT79), .B1(new_n327), .B2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n321), .ZN(new_n335));
  OAI21_X1  g0135(.A(G200), .B1(new_n335), .B2(new_n330), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n324), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n322), .A2(KEYINPUT75), .A3(G200), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n312), .B1(KEYINPUT76), .B2(new_n321), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n329), .A2(new_n330), .ZN(new_n341));
  OAI21_X1  g0141(.A(G190), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT79), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n339), .A2(new_n342), .A3(new_n343), .A4(new_n277), .ZN(new_n344));
  AND2_X1   g0144(.A1(new_n334), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n285), .A2(G1698), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n346), .B(KEYINPUT66), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n279), .A2(new_n280), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n347), .A2(G238), .B1(G107), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n285), .A2(G232), .A3(new_n281), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n307), .B1(new_n351), .B2(new_n317), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n309), .A2(G244), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G179), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n352), .A2(new_n353), .ZN(new_n357));
  INV_X1    g0157(.A(G169), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT15), .B(G87), .ZN(new_n360));
  INV_X1    g0160(.A(new_n360), .ZN(new_n361));
  XOR2_X1   g0161(.A(KEYINPUT8), .B(G58), .Z(new_n362));
  AOI22_X1  g0162(.A1(new_n361), .A2(new_n257), .B1(new_n362), .B2(new_n258), .ZN(new_n363));
  INV_X1    g0163(.A(G77), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n363), .B1(new_n213), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n252), .ZN(new_n366));
  INV_X1    g0166(.A(new_n264), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(new_n364), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n366), .B(new_n368), .C1(new_n364), .C2(new_n273), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n356), .A2(new_n359), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(G58), .A2(G68), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n213), .B1(new_n203), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G159), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n374), .A2(G20), .A3(G33), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT80), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(new_n372), .ZN(new_n377));
  NOR2_X1   g0177(.A1(G58), .A2(G68), .ZN(new_n378));
  OAI21_X1  g0178(.A(G20), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n375), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT80), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT7), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n384), .B1(new_n285), .B2(G20), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n348), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n202), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n271), .B1(new_n388), .B2(KEYINPUT16), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT81), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n278), .B2(G33), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n251), .A2(KEYINPUT81), .A3(KEYINPUT3), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(new_n279), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n393), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT82), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n393), .A2(KEYINPUT82), .A3(KEYINPUT7), .A4(new_n213), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(new_n385), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n383), .B1(new_n398), .B2(G68), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n389), .B1(new_n399), .B2(KEYINPUT16), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n285), .B1(G223), .B2(G1698), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n281), .A2(G226), .ZN(new_n402));
  INV_X1    g0202(.A(G87), .ZN(new_n403));
  OAI22_X1  g0203(.A1(new_n401), .A2(new_n402), .B1(new_n251), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n317), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n307), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n309), .A2(G232), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n405), .A2(G190), .A3(new_n406), .A4(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(G200), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n362), .A2(new_n264), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n263), .B1(new_n250), .B2(new_n254), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n411), .B1(new_n412), .B2(new_n362), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n400), .A2(new_n408), .A3(new_n410), .A4(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT17), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n415), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n400), .A2(new_n413), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n409), .A2(G169), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n355), .B2(new_n409), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT18), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  AND3_X1   g0221(.A1(new_n418), .A2(KEYINPUT18), .A3(new_n420), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n416), .B(new_n417), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n371), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n369), .B1(new_n354), .B2(G190), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n357), .A2(G200), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n345), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT10), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n347), .A2(G223), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n348), .A2(G77), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n285), .A2(G222), .A3(new_n281), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n433), .A2(new_n317), .B1(G226), .B2(new_n309), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n406), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(G200), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(G190), .A3(new_n406), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G50), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n264), .A2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n412), .B2(new_n439), .ZN(new_n441));
  XNOR2_X1  g0241(.A(new_n441), .B(KEYINPUT70), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n362), .A2(new_n257), .B1(G150), .B2(new_n258), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n443), .B(KEYINPUT69), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n204), .A2(new_n213), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n256), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(KEYINPUT9), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT9), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n442), .A2(new_n449), .A3(new_n446), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n429), .B1(new_n438), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n448), .A2(KEYINPUT71), .A3(new_n450), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n453), .A2(new_n429), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT72), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT71), .ZN(new_n456));
  INV_X1    g0256(.A(new_n450), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n449), .B1(new_n442), .B2(new_n446), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n454), .A2(new_n455), .A3(new_n438), .A4(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n459), .A2(new_n438), .A3(new_n453), .A4(new_n429), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT72), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n452), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n435), .A2(new_n358), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n464), .B(new_n447), .C1(G179), .C2(new_n435), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(G179), .B1(new_n340), .B2(new_n341), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n322), .A2(G169), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT14), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT14), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n322), .A2(new_n470), .A3(G169), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n467), .A2(new_n469), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(new_n277), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NOR4_X1   g0275(.A1(new_n428), .A2(new_n463), .A3(new_n466), .A4(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  XOR2_X1   g0277(.A(KEYINPUT85), .B(KEYINPUT19), .Z(new_n478));
  INV_X1    g0278(.A(new_n257), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n478), .B1(new_n290), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n285), .A2(new_n213), .A3(G68), .ZN(new_n481));
  XNOR2_X1  g0281(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n482));
  AOI21_X1  g0282(.A(G20), .B1(new_n482), .B2(new_n291), .ZN(new_n483));
  NOR3_X1   g0283(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n480), .B(new_n481), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(new_n252), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n367), .B1(new_n304), .B2(G33), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n255), .A2(G87), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n367), .A2(new_n360), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n486), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(G45), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(G1), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G274), .ZN(new_n493));
  OAI211_X1 g0293(.A(new_n308), .B(G250), .C1(G1), .C2(new_n491), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n279), .A2(new_n280), .A3(G244), .A4(G1698), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G116), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT84), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n285), .A2(new_n498), .A3(G238), .A4(new_n281), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n279), .A2(new_n280), .A3(G238), .A4(new_n281), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT84), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n497), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n493), .B(new_n494), .C1(new_n502), .C2(new_n302), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n490), .B1(new_n504), .B2(G190), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(G200), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n485), .A2(new_n252), .B1(new_n367), .B2(new_n360), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n255), .A2(new_n361), .A3(new_n487), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n503), .A2(new_n358), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n504), .A2(new_n355), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n505), .A2(new_n506), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g0311(.A1(KEYINPUT5), .A2(G41), .ZN(new_n512));
  NOR2_X1   g0312(.A1(KEYINPUT5), .A2(G41), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n492), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AND3_X1   g0314(.A1(new_n514), .A2(G257), .A3(new_n308), .ZN(new_n515));
  OR2_X1    g0315(.A1(new_n514), .A2(new_n306), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n279), .A2(new_n280), .A3(G244), .A4(new_n281), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT4), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n285), .A2(KEYINPUT4), .A3(G244), .A4(new_n281), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n285), .A2(G250), .A3(G1698), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G283), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT83), .ZN(new_n524));
  XNOR2_X1  g0324(.A(new_n523), .B(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n520), .A2(new_n521), .A3(new_n522), .A4(new_n525), .ZN(new_n526));
  AOI211_X1 g0326(.A(new_n515), .B(new_n517), .C1(new_n317), .C2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n355), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n317), .A2(new_n526), .ZN(new_n529));
  INV_X1    g0329(.A(new_n515), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(new_n516), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n358), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n398), .A2(G107), .B1(G77), .B2(new_n258), .ZN(new_n533));
  INV_X1    g0333(.A(G107), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(KEYINPUT6), .A3(G97), .ZN(new_n535));
  XOR2_X1   g0335(.A(G97), .B(G107), .Z(new_n536));
  OAI21_X1  g0336(.A(new_n535), .B1(new_n536), .B2(KEYINPUT6), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G20), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n271), .B1(new_n533), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n264), .A2(G97), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n255), .A2(new_n487), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n540), .B1(new_n542), .B2(G97), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n528), .B(new_n532), .C1(new_n539), .C2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n533), .A2(new_n538), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n252), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n529), .A2(new_n328), .A3(new_n516), .A4(new_n530), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n527), .B2(G200), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(new_n543), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n511), .A2(new_n545), .A3(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n496), .A2(G20), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n279), .A2(new_n280), .A3(new_n213), .A4(G87), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT22), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT22), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n285), .A2(new_n555), .A3(new_n213), .A4(G87), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n552), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT86), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n213), .A2(G107), .ZN(new_n559));
  XNOR2_X1  g0359(.A(new_n559), .B(KEYINPUT23), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n558), .B1(new_n557), .B2(new_n560), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n561), .A2(new_n562), .A3(KEYINPUT24), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT24), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n554), .A2(new_n556), .ZN(new_n565));
  INV_X1    g0365(.A(new_n552), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n566), .A3(new_n560), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT86), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n557), .A2(new_n558), .A3(new_n560), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n564), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n252), .B1(new_n563), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT87), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n367), .A2(new_n534), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT25), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g0376(.A(new_n576), .B(KEYINPUT88), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n574), .A2(new_n575), .ZN(new_n578));
  XNOR2_X1  g0378(.A(new_n578), .B(KEYINPUT89), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n577), .A2(new_n579), .B1(G107), .B2(new_n542), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT24), .B1(new_n561), .B2(new_n562), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n568), .A2(new_n564), .A3(new_n569), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n583), .A2(KEYINPUT87), .A3(new_n252), .ZN(new_n584));
  AND3_X1   g0384(.A1(new_n573), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n285), .B1(G250), .B2(G1698), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n281), .A2(G257), .ZN(new_n587));
  INV_X1    g0387(.A(G294), .ZN(new_n588));
  OAI22_X1  g0388(.A1(new_n586), .A2(new_n587), .B1(new_n251), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n317), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n514), .A2(new_n308), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(G264), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n593), .A2(new_n517), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n328), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(G200), .B2(new_n594), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n551), .B1(new_n585), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(G20), .B1(new_n251), .B2(G97), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n525), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(G116), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(G20), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n252), .A3(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT20), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n599), .A2(KEYINPUT20), .A3(new_n252), .A4(new_n601), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n367), .A2(new_n600), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n487), .A2(G116), .A3(new_n271), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n281), .A2(G257), .ZN(new_n610));
  NAND2_X1  g0410(.A1(G264), .A2(G1698), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n285), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  OAI221_X1 g0412(.A(new_n612), .B1(G303), .B2(new_n285), .C1(new_n299), .C2(new_n301), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n591), .A2(G270), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n516), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n609), .A2(G169), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT21), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n615), .A2(new_n355), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n609), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n609), .A2(new_n615), .A3(KEYINPUT21), .A4(G169), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n618), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n609), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n615), .A2(G200), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n624), .B(new_n625), .C1(new_n328), .C2(new_n615), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n573), .A2(new_n580), .A3(new_n584), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT90), .ZN(new_n629));
  INV_X1    g0429(.A(new_n594), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n358), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n594), .A2(new_n355), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n628), .A2(new_n629), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n629), .B1(new_n628), .B2(new_n634), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n597), .B(new_n627), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n477), .A2(new_n637), .ZN(G372));
  NAND3_X1  g0438(.A1(new_n339), .A2(new_n342), .A3(new_n277), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n474), .B1(new_n640), .B2(new_n370), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n414), .B(KEYINPUT17), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n418), .A2(new_n420), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(KEYINPUT92), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT92), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n418), .A2(new_n645), .A3(new_n420), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n644), .A2(KEYINPUT18), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT18), .ZN(new_n648));
  AND3_X1   g0448(.A1(new_n418), .A2(new_n645), .A3(new_n420), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n645), .B1(new_n418), .B2(new_n420), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n641), .A2(new_n642), .B1(new_n647), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n465), .B1(new_n652), .B2(new_n463), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n628), .A2(new_n634), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n623), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n597), .A2(new_n656), .A3(KEYINPUT91), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT91), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n545), .A2(new_n550), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n573), .A2(new_n596), .A3(new_n580), .A4(new_n584), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(new_n660), .A3(new_n511), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n622), .B1(new_n628), .B2(new_n634), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n658), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n545), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n664), .A2(KEYINPUT26), .A3(new_n511), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT26), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n505), .A2(new_n506), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n509), .A2(new_n510), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n666), .B1(new_n669), .B2(new_n545), .ZN(new_n670));
  AOI22_X1  g0470(.A1(new_n665), .A2(new_n670), .B1(new_n510), .B2(new_n509), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n657), .A2(new_n663), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n654), .B1(new_n477), .B2(new_n673), .ZN(G369));
  INV_X1    g0474(.A(G13), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G20), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n304), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n624), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n622), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n627), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n686), .A2(new_n684), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n685), .B1(new_n687), .B2(KEYINPUT93), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n685), .A2(KEYINPUT93), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  OAI221_X1 g0491(.A(new_n660), .B1(new_n585), .B2(new_n683), .C1(new_n635), .C2(new_n636), .ZN(new_n692));
  INV_X1    g0492(.A(new_n655), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n682), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n693), .A2(new_n683), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n622), .A2(new_n683), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n698), .B1(new_n692), .B2(new_n699), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n697), .A2(new_n700), .ZN(G399));
  INV_X1    g0501(.A(new_n220), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(G41), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n484), .A2(new_n600), .ZN(new_n704));
  NOR3_X1   g0504(.A1(new_n703), .A2(new_n704), .A3(new_n304), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n216), .B2(new_n703), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT94), .ZN(new_n707));
  XOR2_X1   g0507(.A(new_n707), .B(KEYINPUT28), .Z(new_n708));
  INV_X1    g0508(.A(KEYINPUT29), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n672), .A2(new_n709), .A3(new_n683), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n623), .B1(new_n635), .B2(new_n636), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n659), .A2(new_n667), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n711), .A2(new_n660), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n682), .B1(new_n713), .B2(new_n671), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n710), .B1(new_n714), .B2(new_n709), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n615), .A2(new_n593), .A3(new_n355), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(new_n504), .A3(new_n527), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT30), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n504), .A2(new_n527), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n721), .A2(new_n630), .A3(new_n355), .A4(new_n615), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n717), .A2(KEYINPUT30), .A3(new_n504), .A4(new_n527), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n720), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n725));
  AOI21_X1  g0525(.A(KEYINPUT31), .B1(new_n724), .B2(new_n682), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n637), .B2(new_n682), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G330), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n716), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n708), .B1(new_n731), .B2(G1), .ZN(G364));
  INV_X1    g0532(.A(new_n703), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n676), .A2(G45), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(G1), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n702), .A2(new_n285), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n216), .A2(new_n491), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n736), .B(new_n737), .C1(new_n244), .C2(new_n491), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(G116), .B2(new_n220), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n702), .A2(new_n348), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n739), .B1(G355), .B2(new_n740), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT95), .Z(new_n742));
  AOI21_X1  g0542(.A(new_n212), .B1(G20), .B2(new_n358), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G13), .A2(G33), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n735), .B1(new_n742), .B2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n743), .ZN(new_n749));
  NOR4_X1   g0549(.A1(new_n213), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n750), .A2(KEYINPUT96), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(KEYINPUT96), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n374), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT32), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n213), .A2(new_n328), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n355), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G58), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n328), .A2(G179), .A3(G200), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n213), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n763), .A2(KEYINPUT97), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(KEYINPUT97), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n290), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n325), .A2(G179), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n756), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n213), .A2(G190), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n757), .A2(new_n771), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n770), .A2(new_n403), .B1(new_n772), .B2(new_n364), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n771), .A2(new_n769), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n355), .A2(new_n325), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n756), .A2(new_n775), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n285), .B1(new_n774), .B2(new_n534), .C1(new_n439), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n775), .A2(new_n771), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI211_X1 g0579(.A(new_n773), .B(new_n777), .C1(G68), .C2(new_n779), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n755), .A2(new_n760), .A3(new_n768), .A4(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G311), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n772), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G283), .ZN(new_n784));
  INV_X1    g0584(.A(G326), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n348), .B1(new_n774), .B2(new_n784), .C1(new_n785), .C2(new_n776), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n783), .B(new_n786), .C1(G294), .C2(new_n763), .ZN(new_n787));
  XNOR2_X1  g0587(.A(new_n770), .B(KEYINPUT98), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G303), .ZN(new_n790));
  XNOR2_X1  g0590(.A(KEYINPUT33), .B(G317), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n779), .A2(new_n791), .B1(new_n759), .B2(G322), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT99), .ZN(new_n793));
  INV_X1    g0593(.A(new_n753), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G329), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n787), .A2(new_n790), .A3(new_n793), .A4(new_n795), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n781), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n746), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n748), .B1(new_n749), .B2(new_n797), .C1(new_n690), .C2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n691), .A2(new_n735), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n690), .A2(G330), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(G396));
  NAND2_X1  g0602(.A1(new_n672), .A2(new_n683), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n371), .A2(new_n683), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n425), .A2(new_n426), .B1(new_n369), .B2(new_n682), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n371), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  MUX2_X1   g0607(.A(new_n682), .B(new_n805), .S(new_n370), .Z(new_n808));
  NAND3_X1  g0608(.A1(new_n672), .A2(new_n683), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n729), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n807), .A2(G330), .A3(new_n728), .A4(new_n809), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n735), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT100), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n743), .A2(new_n744), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n364), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G143), .A2(new_n759), .B1(new_n779), .B2(G150), .ZN(new_n818));
  INV_X1    g0618(.A(new_n776), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(G137), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n818), .B(new_n820), .C1(new_n374), .C2(new_n772), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT34), .Z(new_n822));
  NOR2_X1   g0622(.A1(new_n774), .A2(new_n202), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n794), .A2(G132), .B1(G58), .B2(new_n763), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n439), .B2(new_n788), .ZN(new_n825));
  NOR4_X1   g0625(.A1(new_n822), .A2(new_n348), .A3(new_n823), .A4(new_n825), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n753), .A2(new_n782), .B1(new_n788), .B2(new_n534), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G283), .A2(new_n779), .B1(new_n759), .B2(G294), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n285), .B1(new_n819), .B2(G303), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n828), .B(new_n829), .C1(new_n600), .C2(new_n772), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n774), .A2(new_n403), .ZN(new_n831));
  NOR4_X1   g0631(.A1(new_n767), .A2(new_n827), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n743), .B1(new_n826), .B2(new_n832), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n817), .B(new_n833), .C1(new_n808), .C2(new_n745), .ZN(new_n834));
  INV_X1    g0634(.A(new_n735), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n814), .A2(new_n815), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n835), .B1(new_n811), .B2(new_n812), .ZN(new_n838));
  INV_X1    g0638(.A(new_n836), .ZN(new_n839));
  OAI21_X1  g0639(.A(KEYINPUT100), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n837), .A2(new_n840), .ZN(G384));
  AND3_X1   g0641(.A1(new_n467), .A2(new_n469), .A3(new_n471), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n334), .A2(new_n842), .A3(new_n344), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n277), .A2(new_n683), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n844), .B1(new_n472), .B2(new_n473), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n639), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n806), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n388), .A2(KEYINPUT16), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT16), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n850), .B1(new_n383), .B2(new_n387), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n849), .A2(new_n256), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(new_n413), .ZN(new_n853));
  INV_X1    g0653(.A(new_n680), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n423), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT104), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(new_n418), .B2(new_n854), .ZN(new_n859));
  AOI211_X1 g0659(.A(KEYINPUT104), .B(new_n680), .C1(new_n400), .C2(new_n413), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n643), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n414), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n853), .B1(new_n420), .B2(new_n854), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n864), .A2(new_n414), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n861), .A2(new_n863), .B1(new_n865), .B2(new_n862), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n857), .A2(new_n866), .A3(KEYINPUT105), .A4(KEYINPUT38), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT38), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n862), .B1(new_n864), .B2(new_n414), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n418), .A2(new_n420), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n418), .A2(new_n854), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT104), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n418), .A2(new_n858), .A3(new_n854), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n863), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n869), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n643), .A2(new_n648), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n418), .A2(KEYINPUT18), .A3(new_n420), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n855), .B1(new_n642), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n868), .B1(new_n876), .B2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT105), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n857), .A2(new_n866), .A3(KEYINPUT38), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n848), .A2(new_n728), .A3(new_n867), .A4(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT40), .ZN(new_n886));
  INV_X1    g0686(.A(new_n728), .ZN(new_n887));
  AOI22_X1  g0687(.A1(new_n843), .A2(new_n844), .B1(new_n639), .B2(new_n846), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n887), .A2(new_n888), .A3(new_n806), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n414), .B1(new_n649), .B2(new_n650), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n859), .A2(new_n860), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT106), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n874), .A2(new_n893), .A3(new_n875), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT106), .B1(new_n861), .B2(new_n863), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n891), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n651), .A2(new_n647), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n897), .B1(new_n898), .B2(new_n642), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n868), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n886), .B1(new_n900), .B2(new_n883), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n885), .A2(new_n886), .B1(new_n889), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n476), .A2(new_n728), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n902), .B(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(G330), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n898), .A2(new_n854), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT103), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n804), .B(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n888), .B1(new_n809), .B2(new_n908), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n884), .A2(new_n867), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n906), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n884), .A2(new_n867), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(KEYINPUT39), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n474), .A2(new_n682), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT39), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n898), .A2(new_n642), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n891), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n892), .A2(new_n894), .A3(new_n895), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT38), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n883), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n915), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n913), .A2(new_n914), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n911), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n653), .B1(new_n476), .B2(new_n715), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n923), .B(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n905), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n304), .B2(new_n676), .ZN(new_n927));
  XOR2_X1   g0727(.A(new_n537), .B(KEYINPUT101), .Z(new_n928));
  AOI21_X1  g0728(.A(new_n600), .B1(new_n928), .B2(KEYINPUT35), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n929), .B(new_n214), .C1(KEYINPUT35), .C2(new_n928), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT102), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT36), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n372), .A2(G77), .ZN(new_n933));
  OAI22_X1  g0733(.A1(new_n215), .A2(new_n933), .B1(G50), .B2(new_n202), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(G1), .A3(new_n675), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n927), .A2(new_n932), .A3(new_n935), .ZN(G367));
  INV_X1    g0736(.A(KEYINPUT42), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n682), .B1(new_n539), .B2(new_n544), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n659), .A2(new_n938), .ZN(new_n939));
  OR3_X1    g0739(.A1(new_n692), .A2(new_n699), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(KEYINPUT109), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n940), .A2(KEYINPUT109), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n937), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n943), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n945), .A2(KEYINPUT42), .A3(new_n941), .ZN(new_n946));
  INV_X1    g0746(.A(new_n636), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n628), .A2(new_n629), .A3(new_n634), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n545), .B1(new_n949), .B2(new_n939), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n683), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n944), .A2(new_n946), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n490), .A2(new_n682), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n511), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n668), .B2(new_n953), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT107), .Z(new_n956));
  XOR2_X1   g0756(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n959));
  AND3_X1   g0759(.A1(new_n952), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n958), .B1(new_n952), .B2(new_n959), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT110), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n664), .A2(new_n682), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n939), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n697), .A2(new_n964), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n960), .A2(new_n961), .B1(new_n962), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n962), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n962), .B(new_n965), .C1(new_n960), .C2(new_n961), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n703), .B(KEYINPUT41), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(KEYINPUT111), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n700), .A2(new_n939), .A3(new_n963), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT44), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n973), .B(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n697), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n698), .B(new_n964), .C1(new_n692), .C2(new_n699), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT45), .Z(new_n978));
  AND3_X1   g0778(.A1(new_n975), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n976), .B1(new_n975), .B2(new_n978), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n972), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n696), .A2(new_n699), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n692), .B2(new_n699), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(new_n691), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n984), .A2(new_n730), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n975), .A2(new_n978), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n697), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(KEYINPUT111), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n981), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n971), .B1(new_n989), .B2(new_n731), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n734), .A2(G1), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n968), .B(new_n969), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  INV_X1    g0792(.A(new_n736), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n747), .B1(new_n220), .B2(new_n360), .C1(new_n240), .C2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n835), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT112), .Z(new_n996));
  AND2_X1   g0796(.A1(new_n794), .A2(G137), .ZN(new_n997));
  INV_X1    g0797(.A(new_n774), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n348), .B1(new_n998), .B2(G77), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n439), .B2(new_n772), .C1(new_n201), .C2(new_n770), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n766), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(G68), .ZN(new_n1002));
  INV_X1    g0802(.A(G143), .ZN(new_n1003));
  INV_X1    g0803(.A(G150), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1002), .B1(new_n1003), .B2(new_n776), .C1(new_n1004), .C2(new_n758), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n997), .B(new_n1000), .C1(new_n1005), .C2(KEYINPUT114), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(KEYINPUT114), .B2(new_n1005), .C1(new_n374), .C2(new_n778), .ZN(new_n1007));
  INV_X1    g0807(.A(G317), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n753), .A2(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(G294), .A2(new_n779), .B1(new_n759), .B2(G303), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n290), .B2(new_n774), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n770), .ZN(new_n1012));
  AOI21_X1  g0812(.A(KEYINPUT46), .B1(new_n1012), .B2(G116), .ZN(new_n1013));
  NOR3_X1   g0813(.A1(new_n1011), .A2(new_n285), .A3(new_n1013), .ZN(new_n1014));
  OAI22_X1  g0814(.A1(new_n762), .A2(new_n534), .B1(new_n772), .B2(new_n784), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT113), .Z(new_n1016));
  NAND2_X1  g0816(.A1(new_n819), .A2(G311), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n789), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1007), .B1(new_n1009), .B2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT47), .Z(new_n1021));
  OAI221_X1 g0821(.A(new_n996), .B1(new_n955), .B2(new_n798), .C1(new_n1021), .C2(new_n749), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n992), .A2(new_n1022), .ZN(G387));
  AOI22_X1  g0823(.A1(G311), .A2(new_n779), .B1(new_n759), .B2(G317), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n819), .A2(G322), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n772), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(G303), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1024), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT48), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n784), .B2(new_n762), .C1(new_n588), .C2(new_n770), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT49), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1033), .B(new_n348), .C1(new_n785), .C2(new_n753), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1032), .B(new_n1034), .C1(G116), .C2(new_n998), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n285), .B1(new_n772), .B2(new_n202), .C1(new_n290), .C2(new_n774), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G77), .A2(new_n1012), .B1(new_n779), .B2(new_n362), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n439), .B2(new_n758), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(KEYINPUT115), .B(G150), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1036), .B(new_n1038), .C1(new_n794), .C2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1001), .A2(new_n361), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(new_n374), .C2(new_n776), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT116), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n743), .B1(new_n1035), .B2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n993), .B1(new_n237), .B2(G45), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n704), .B2(new_n740), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n362), .A2(new_n439), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n704), .B1(new_n1047), .B2(KEYINPUT50), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1048), .B(new_n491), .C1(KEYINPUT50), .C2(new_n1047), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(G68), .B2(G77), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n1046), .A2(new_n1050), .B1(G107), .B2(new_n220), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n735), .B1(new_n1051), .B2(new_n747), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1044), .B(new_n1052), .C1(new_n695), .C2(new_n798), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n991), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n984), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n703), .B1(new_n1055), .B2(new_n731), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1053), .B1(new_n1054), .B2(new_n984), .C1(new_n1056), .C2(new_n985), .ZN(G393));
  NAND3_X1  g0857(.A1(new_n975), .A2(new_n976), .A3(new_n978), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n987), .A2(new_n991), .A3(new_n1058), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n747), .B1(new_n290), .B2(new_n220), .C1(new_n247), .C2(new_n993), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT117), .Z(new_n1061));
  NOR2_X1   g0861(.A1(new_n766), .A2(new_n364), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n362), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n1063), .A2(new_n772), .B1(new_n202), .B2(new_n770), .ZN(new_n1064));
  NOR4_X1   g0864(.A1(new_n1062), .A2(new_n348), .A3(new_n831), .A4(new_n1064), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G150), .A2(new_n819), .B1(new_n759), .B2(G159), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n1066), .A2(KEYINPUT51), .B1(new_n753), .B2(new_n1003), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(KEYINPUT51), .B2(new_n1066), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1065), .B(new_n1068), .C1(new_n439), .C2(new_n778), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n794), .A2(G322), .B1(G107), .B2(new_n998), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n776), .A2(new_n1008), .B1(new_n758), .B2(new_n782), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT52), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n285), .B1(new_n1012), .B2(G283), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1070), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n762), .A2(new_n600), .B1(new_n772), .B2(new_n588), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(G303), .B2(new_n779), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT118), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1069), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1061), .B1(new_n1078), .B2(new_n743), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n835), .B(new_n1079), .C1(new_n964), .C2(new_n798), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1059), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n987), .A2(new_n1058), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n730), .B2(new_n984), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n989), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1081), .B1(new_n1084), .B2(new_n703), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(G390));
  NOR3_X1   g0886(.A1(new_n463), .A2(new_n466), .A3(new_n475), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n428), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1087), .A2(new_n1088), .A3(G330), .A4(new_n728), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n845), .A2(new_n847), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1090), .A2(G330), .A3(new_n728), .A4(new_n808), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n804), .B(KEYINPUT103), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n714), .B2(new_n808), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n728), .A2(G330), .A3(new_n808), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n888), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1091), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1096), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1091), .A2(new_n1095), .B1(new_n809), .B2(new_n908), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n924), .B(new_n1089), .C1(new_n1097), .C2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT39), .B1(new_n900), .B2(new_n883), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n915), .B1(new_n884), .B2(new_n867), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n1100), .A2(new_n1101), .B1(new_n909), .B2(new_n914), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n914), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n900), .A2(new_n883), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1103), .B(new_n1104), .C1(new_n1093), .C2(new_n888), .ZN(new_n1105));
  AND3_X1   g0905(.A1(new_n1102), .A2(new_n1105), .A3(new_n1091), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1091), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1099), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1091), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n809), .A2(new_n908), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n1090), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1111), .A2(new_n1103), .B1(new_n913), .B2(new_n921), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1103), .B1(new_n919), .B2(new_n920), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n713), .A2(new_n671), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1114), .A2(new_n683), .A3(new_n808), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n908), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1113), .B1(new_n1116), .B2(new_n1090), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1109), .B1(new_n1112), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1102), .A2(new_n1105), .A3(new_n1091), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n476), .A2(new_n715), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1120), .A2(new_n654), .A3(new_n1089), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1091), .A2(new_n1095), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n1110), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n1096), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n1118), .A2(new_n1119), .A3(new_n1121), .A4(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1108), .A2(new_n1125), .A3(new_n703), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n744), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1062), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G107), .A2(new_n779), .B1(new_n759), .B2(G116), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1129), .B1(new_n784), .B2(new_n776), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n1130), .A2(new_n285), .A3(new_n823), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1026), .A2(G97), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(G294), .A2(new_n794), .B1(new_n789), .B2(G87), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1128), .A2(new_n1131), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(G132), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n285), .B1(new_n758), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n819), .A2(G128), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n779), .A2(G137), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT54), .B(G143), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1137), .B(new_n1138), .C1(new_n772), .C2(new_n1139), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1136), .B(new_n1140), .C1(G50), .C2(new_n998), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n794), .A2(G125), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(new_n374), .C2(new_n766), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1012), .A2(new_n1039), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT53), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1134), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1146), .A2(new_n743), .B1(new_n1063), .B2(new_n816), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1127), .A2(new_n835), .A3(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1148), .B1(new_n1149), .B2(new_n991), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1126), .A2(new_n1150), .ZN(G378));
  NAND3_X1  g0951(.A1(new_n1090), .A2(new_n728), .A3(new_n808), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n886), .B1(new_n1152), .B2(new_n912), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1104), .A2(KEYINPUT40), .A3(new_n728), .A4(new_n848), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(G330), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1155), .A2(new_n922), .A3(new_n911), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n923), .A2(new_n902), .A3(G330), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n463), .A2(new_n466), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT55), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1159), .B(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n447), .A2(new_n854), .ZN(new_n1162));
  XOR2_X1   g0962(.A(new_n1162), .B(KEYINPUT56), .Z(new_n1163));
  XOR2_X1   g0963(.A(new_n1161), .B(new_n1163), .Z(new_n1164));
  NAND2_X1  g0964(.A1(new_n1158), .A2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1161), .B(new_n1163), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1166), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1054), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n744), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1002), .B1(new_n600), .B2(new_n776), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT120), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G97), .A2(new_n779), .B1(new_n998), .B2(G58), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n534), .B2(new_n758), .ZN(new_n1173));
  INV_X1    g0973(.A(G41), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1174), .B(new_n348), .C1(new_n770), .C2(new_n364), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT119), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1173), .B(new_n1176), .C1(new_n794), .C2(G283), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1171), .B(new_n1177), .C1(new_n360), .C2(new_n772), .ZN(new_n1178));
  XOR2_X1   g0978(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n1179));
  OR2_X1    g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G128), .A2(new_n759), .B1(new_n779), .B2(G132), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n819), .A2(G125), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(new_n770), .C2(new_n1139), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n766), .A2(new_n1004), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1183), .B(new_n1184), .C1(G137), .C2(new_n1026), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(new_n1185), .B(KEYINPUT59), .ZN(new_n1186));
  AOI21_X1  g0986(.A(G41), .B1(new_n794), .B2(G124), .ZN(new_n1187));
  AOI21_X1  g0987(.A(G33), .B1(new_n998), .B2(G159), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1174), .B1(new_n278), .B2(new_n251), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n439), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1180), .A2(new_n1189), .A3(new_n1190), .A4(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n1193), .A2(new_n743), .B1(new_n439), .B2(new_n816), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1169), .A2(new_n835), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1168), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1125), .A2(new_n1121), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n1166), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1166), .B1(new_n1157), .B2(new_n1156), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1198), .B(KEYINPUT57), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n703), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1165), .A2(new_n1167), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT57), .B1(new_n1203), .B2(new_n1198), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1197), .B1(new_n1202), .B2(new_n1204), .ZN(G375));
  AOI21_X1  g1005(.A(new_n1054), .B1(new_n1123), .B2(new_n1096), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n888), .A2(new_n744), .ZN(new_n1207));
  AOI22_X1  g1007(.A1(G128), .A2(new_n794), .B1(new_n789), .B2(G159), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n285), .B1(new_n774), .B2(new_n201), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n776), .A2(new_n1135), .B1(new_n778), .B2(new_n1139), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1209), .B(new_n1210), .C1(G137), .C2(new_n759), .ZN(new_n1211));
  AND2_X1   g1011(.A1(new_n1208), .A2(new_n1211), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n439), .B2(new_n766), .C1(new_n1004), .C2(new_n772), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n758), .A2(new_n784), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G303), .A2(new_n794), .B1(new_n789), .B2(G97), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n348), .B1(new_n774), .B2(new_n364), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n776), .A2(new_n588), .B1(new_n778), .B2(new_n600), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1216), .B(new_n1217), .C1(G107), .C2(new_n1026), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1041), .A2(new_n1215), .A3(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1213), .B1(new_n1214), .B2(new_n1219), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n1220), .A2(new_n743), .B1(new_n202), .B2(new_n816), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1207), .A2(new_n835), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  OR3_X1    g1023(.A1(new_n1206), .A2(KEYINPUT122), .A3(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(KEYINPUT122), .B1(new_n1206), .B2(new_n1223), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n924), .A2(new_n1089), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1229), .A2(new_n970), .A3(new_n1099), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n1226), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(G381));
  AOI22_X1  g1032(.A1(new_n1165), .A2(new_n1167), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n733), .B1(new_n1233), .B2(KEYINPUT57), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT57), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1198), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1234), .A2(new_n1238), .ZN(new_n1239));
  NOR3_X1   g1039(.A1(G378), .A2(new_n1168), .A3(new_n1196), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1241), .A2(G384), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(G393), .A2(G396), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n992), .A2(new_n1085), .A3(new_n1022), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1242), .A2(new_n1231), .A3(new_n1243), .A4(new_n1245), .ZN(G407));
  OAI211_X1 g1046(.A(G407), .B(G213), .C1(G343), .C2(new_n1241), .ZN(G409));
  XNOR2_X1  g1047(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n1248));
  AND2_X1   g1048(.A1(new_n681), .A2(G213), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1233), .A2(new_n970), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1249), .B1(new_n1240), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(G378), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1195), .B1(new_n1236), .B2(new_n1054), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n1234), .B2(new_n1238), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1251), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT60), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1229), .A2(new_n1256), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1227), .A2(KEYINPUT60), .A3(new_n1228), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1257), .A2(new_n703), .A3(new_n1099), .A4(new_n1258), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n837), .A2(new_n840), .A3(KEYINPUT123), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(new_n1226), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1249), .A2(G2897), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1258), .A2(new_n703), .A3(new_n1099), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n1264), .A2(new_n1257), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT123), .B1(new_n837), .B2(new_n840), .ZN(new_n1266));
  OR2_X1    g1066(.A1(new_n1260), .A2(new_n1266), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1261), .B(new_n1263), .C1(new_n1265), .C2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1259), .A2(new_n1226), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1260), .A2(new_n1266), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1263), .B1(new_n1272), .B2(new_n1261), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1269), .A2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1248), .B1(new_n1255), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(G375), .A2(G378), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1272), .A2(new_n1261), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1276), .A2(new_n1251), .A3(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT62), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1279), .A2(KEYINPUT125), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1276), .A2(new_n1251), .A3(new_n1277), .A4(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1275), .A2(new_n1281), .A3(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT126), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  XOR2_X1   g1086(.A(G393), .B(G396), .Z(new_n1287));
  AOI21_X1  g1087(.A(new_n1085), .B1(new_n992), .B2(new_n1022), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1287), .B1(new_n1245), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(G387), .A2(G390), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1287), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(new_n1291), .A3(new_n1244), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1289), .A2(new_n1292), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1275), .A2(new_n1281), .A3(KEYINPUT126), .A4(new_n1283), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1286), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  AND2_X1   g1095(.A1(new_n1255), .A2(new_n1274), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT63), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1278), .B1(new_n1296), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1293), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT61), .ZN(new_n1300));
  OR2_X1    g1100(.A1(new_n1278), .A2(new_n1297), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .A4(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1295), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(KEYINPUT127), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT127), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1295), .A2(new_n1302), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1304), .A2(new_n1306), .ZN(G405));
  NAND2_X1  g1107(.A1(new_n1299), .A2(new_n1277), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1293), .A2(new_n1272), .A3(new_n1261), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1276), .A2(new_n1241), .ZN(new_n1311));
  XNOR2_X1  g1111(.A(new_n1310), .B(new_n1311), .ZN(G402));
endmodule


