// Benchmark "locked_c2670" written by ABC on Sat Dec 16 10:59:06 2023

module locked_c2670 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6,
    G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26,
    G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48,
    G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64,
    G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80,
    G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96,
    G99, G100, G101, G102, G103, G104, G105, G106, G107, G108, G111, G112,
    G113, G114, G115, G116, G117, G118, G119, G120, G123, G124, G125, G126,
    G127, G128, G129, G130, G131, G132, G135, G136, G137, G138, G139, G140,
    G141, G142, G169, G174, G177, G178, G179, G180, G181, G182, G183, G184,
    G185, G186, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198,
    G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210,
    G211, G212, G213, G214, G215, G239, G240, G241, G242, G243, G244, G245,
    G246, G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
    G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272, G273,
    G274, G275, G276, G277, G278, G279, G452, G483, G543, G559, G567, G651,
    G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966,
    G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078,
    G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435,
    G2438, G2443, G2446, G2451, G2454, G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3,
    G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22, G23, G24,
    G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40, G43, G44,
    G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60, G61, G62,
    G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76, G77, G78,
    G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92, G93, G94,
    G95, G96, G99, G100, G101, G102, G103, G104, G105, G106, G107, G108,
    G111, G112, G113, G114, G115, G116, G117, G118, G119, G120, G123, G124,
    G125, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G138,
    G139, G140, G141, G142, G169, G174, G177, G178, G179, G180, G181, G182,
    G183, G184, G185, G186, G189, G190, G191, G192, G193, G194, G195, G196,
    G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208,
    G209, G210, G211, G212, G213, G214, G215, G239, G240, G241, G242, G243,
    G244, G245, G246, G247, G248, G249, G250, G251, G252, G253, G254, G255,
    G256, G257, G262, G263, G264, G265, G266, G267, G268, G269, G270, G271,
    G272, G273, G274, G275, G276, G277, G278, G279, G452, G483, G543, G559,
    G567, G651, G661, G860, G868, G1083, G1341, G1348, G1384, G1956, G1961,
    G1966, G1971, G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072,
    G2078, G2084, G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430,
    G2435, G2438, G2443, G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n382, new_n386, new_n387, new_n388, new_n389, new_n392, new_n393,
    new_n394, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n409,
    new_n410, new_n411, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n439, new_n440,
    new_n441, new_n442, new_n443, new_n444, new_n445, new_n446, new_n447,
    new_n449, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n468, new_n469, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n484,
    new_n485, new_n486, new_n487, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n495, new_n496, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n513, new_n516, new_n517, new_n519, new_n520,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n579, new_n580, new_n581, new_n582,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n595, new_n596,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n606, new_n607, new_n608, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n930, new_n931;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n382));
  XOR2_X1   g021(.A(new_n382), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n386));
  XOR2_X1   g025(.A(new_n386), .B(KEYINPUT2), .Z(new_n387));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n388));
  INV_X1    g027(.A(new_n388), .ZN(new_n389));
  NOR2_X1   g028(.A1(new_n387), .A2(new_n389), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n387), .A2(G2106), .ZN(new_n392));
  NAND2_X1  g031(.A1(new_n389), .A2(G567), .ZN(new_n393));
  NAND2_X1  g032(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g033(.A(new_n394), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n396));
  INV_X1    g035(.A(G2104), .ZN(new_n397));
  NAND2_X1  g036(.A1(new_n397), .A2(KEYINPUT3), .ZN(new_n398));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n399));
  NAND2_X1  g038(.A1(new_n399), .A2(G2104), .ZN(new_n400));
  NAND3_X1  g039(.A1(new_n398), .A2(new_n400), .A3(G125), .ZN(new_n401));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n402));
  AOI21_X1  g041(.A(new_n396), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND4_X1  g042(.A1(new_n398), .A2(new_n400), .A3(G137), .A4(new_n396), .ZN(new_n404));
  NOR2_X1   g043(.A1(new_n397), .A2(G2105), .ZN(new_n405));
  NAND2_X1  g044(.A1(new_n405), .A2(G101), .ZN(new_n406));
  NAND2_X1  g045(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g046(.A1(new_n403), .A2(new_n407), .ZN(G160));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n409));
  MUX2_X1   g048(.A(G136), .B(G124), .S(G2105), .Z(new_n410));
  MUX2_X1   g049(.A(G100), .B(G112), .S(G2105), .Z(new_n411));
  AOI22_X1  g050(.A1(new_n409), .A2(new_n410), .B1(new_n411), .B2(G2104), .ZN(G162));
  NAND2_X1  g051(.A1(G114), .A2(G2105), .ZN(new_n413));
  INV_X1    g052(.A(G102), .ZN(new_n414));
  OAI21_X1  g053(.A(new_n413), .B1(new_n414), .B2(G2105), .ZN(new_n415));
  NAND2_X1  g054(.A1(new_n415), .A2(G2104), .ZN(new_n416));
  NAND4_X1  g055(.A1(new_n398), .A2(new_n400), .A3(G126), .A4(G2105), .ZN(new_n417));
  NAND2_X1  g056(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g057(.A1(new_n398), .A2(new_n400), .A3(G138), .A4(new_n396), .ZN(new_n419));
  NAND2_X1  g058(.A1(new_n419), .A2(KEYINPUT4), .ZN(new_n420));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n421));
  NAND4_X1  g060(.A1(new_n409), .A2(new_n421), .A3(G138), .A4(new_n396), .ZN(new_n422));
  AOI21_X1  g061(.A(new_n418), .B1(new_n420), .B2(new_n422), .ZN(G164));
  INV_X1    g062(.A(G543), .ZN(new_n424));
  NAND2_X1  g063(.A1(new_n424), .A2(KEYINPUT5), .ZN(new_n425));
  INV_X1    g064(.A(KEYINPUT5), .ZN(new_n426));
  NAND2_X1  g065(.A1(new_n426), .A2(G543), .ZN(new_n427));
  AND2_X1   g066(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  AOI22_X1  g067(.A1(new_n428), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n429));
  INV_X1    g068(.A(G651), .ZN(new_n430));
  NOR2_X1   g069(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI22_X1  g070(.A1(new_n428), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n432));
  NAND2_X1  g071(.A1(new_n430), .A2(KEYINPUT6), .ZN(new_n433));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n434));
  NAND2_X1  g073(.A1(new_n434), .A2(G651), .ZN(new_n435));
  NAND2_X1  g074(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g075(.A1(new_n432), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g076(.A1(new_n431), .A2(new_n437), .ZN(G166));
  NAND3_X1  g077(.A1(new_n428), .A2(G63), .A3(G651), .ZN(new_n439));
  NAND3_X1  g078(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n440));
  XNOR2_X1  g079(.A(new_n440), .B(KEYINPUT7), .ZN(new_n441));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n442));
  NAND3_X1  g081(.A1(new_n442), .A2(G51), .A3(G543), .ZN(new_n443));
  NAND3_X1  g082(.A1(new_n439), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g083(.A1(new_n425), .A2(new_n427), .ZN(new_n445));
  NOR2_X1   g084(.A1(new_n445), .A2(new_n436), .ZN(new_n446));
  AND2_X1   g085(.A1(new_n446), .A2(G89), .ZN(new_n447));
  NOR2_X1   g086(.A1(new_n444), .A2(new_n447), .ZN(G168));
  NAND2_X1  g087(.A1(G77), .A2(G543), .ZN(new_n449));
  INV_X1    g088(.A(G64), .ZN(new_n450));
  OAI21_X1  g089(.A(new_n449), .B1(new_n445), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g090(.A1(new_n451), .A2(G651), .ZN(new_n452));
  NAND2_X1  g091(.A1(G52), .A2(G543), .ZN(new_n453));
  INV_X1    g092(.A(G90), .ZN(new_n454));
  OAI21_X1  g093(.A(new_n453), .B1(new_n445), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g094(.A1(new_n455), .A2(new_n442), .ZN(new_n456));
  NAND2_X1  g095(.A1(new_n452), .A2(new_n456), .ZN(G301));
  INV_X1    g096(.A(G301), .ZN(G171));
  AOI22_X1  g097(.A1(new_n428), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n459));
  OR2_X1    g098(.A1(new_n459), .A2(new_n430), .ZN(new_n460));
  AOI22_X1  g099(.A1(new_n428), .A2(G81), .B1(G43), .B2(G543), .ZN(new_n461));
  OR2_X1    g100(.A1(new_n461), .A2(new_n436), .ZN(new_n462));
  NAND2_X1  g101(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g102(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g103(.A1(new_n464), .A2(G860), .ZN(G153));
  AND3_X1   g104(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n466));
  NAND2_X1  g105(.A1(new_n466), .A2(G36), .ZN(G176));
  NAND2_X1  g106(.A1(G1), .A2(G3), .ZN(new_n468));
  XNOR2_X1  g107(.A(new_n468), .B(KEYINPUT8), .ZN(new_n469));
  NAND2_X1  g108(.A1(new_n466), .A2(new_n469), .ZN(G188));
  NAND2_X1  g109(.A1(G53), .A2(G543), .ZN(new_n471));
  OAI21_X1  g110(.A(KEYINPUT9), .B1(new_n436), .B2(new_n471), .ZN(new_n472));
  INV_X1    g111(.A(KEYINPUT9), .ZN(new_n473));
  NAND4_X1  g112(.A1(new_n442), .A2(new_n473), .A3(G53), .A4(G543), .ZN(new_n474));
  NAND2_X1  g113(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g114(.A1(G78), .A2(G543), .ZN(new_n476));
  INV_X1    g115(.A(G65), .ZN(new_n477));
  OAI21_X1  g116(.A(new_n476), .B1(new_n445), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g117(.A1(new_n478), .A2(G651), .ZN(new_n479));
  NAND2_X1  g118(.A1(new_n446), .A2(G91), .ZN(new_n480));
  NAND3_X1  g119(.A1(new_n475), .A2(new_n479), .A3(new_n480), .ZN(G299));
  INV_X1    g120(.A(G168), .ZN(G286));
  OR2_X1    g121(.A1(new_n431), .A2(new_n437), .ZN(G303));
  AOI22_X1  g122(.A1(new_n428), .A2(G87), .B1(G49), .B2(G543), .ZN(new_n484));
  NOR2_X1   g123(.A1(new_n484), .A2(new_n436), .ZN(new_n485));
  INV_X1    g124(.A(G74), .ZN(new_n486));
  AOI21_X1  g125(.A(new_n430), .B1(new_n445), .B2(new_n486), .ZN(new_n487));
  OR2_X1    g126(.A1(new_n485), .A2(new_n487), .ZN(G288));
  AOI22_X1  g127(.A1(new_n428), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n489));
  NOR2_X1   g128(.A1(new_n489), .A2(new_n430), .ZN(new_n490));
  AOI22_X1  g129(.A1(new_n428), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n491));
  NOR2_X1   g130(.A1(new_n491), .A2(new_n436), .ZN(new_n492));
  NOR2_X1   g131(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g132(.A(new_n493), .ZN(G305));
  AOI22_X1  g133(.A1(new_n428), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n495));
  AOI22_X1  g134(.A1(new_n428), .A2(G85), .B1(G47), .B2(G543), .ZN(new_n496));
  OAI22_X1  g135(.A1(new_n430), .A2(new_n495), .B1(new_n496), .B2(new_n436), .ZN(G290));
  INV_X1    g136(.A(KEYINPUT10), .ZN(new_n498));
  NAND2_X1  g137(.A1(new_n428), .A2(new_n442), .ZN(new_n499));
  INV_X1    g138(.A(G92), .ZN(new_n500));
  OAI21_X1  g139(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g140(.A1(new_n446), .A2(KEYINPUT10), .A3(G92), .ZN(new_n502));
  NAND2_X1  g141(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g142(.A1(G79), .A2(G543), .ZN(new_n504));
  INV_X1    g143(.A(G66), .ZN(new_n505));
  OAI21_X1  g144(.A(new_n504), .B1(new_n445), .B2(new_n505), .ZN(new_n506));
  AND2_X1   g145(.A1(G54), .A2(G543), .ZN(new_n507));
  AOI22_X1  g146(.A1(new_n506), .A2(G651), .B1(new_n442), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g147(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g148(.A1(new_n509), .A2(G868), .ZN(new_n510));
  AOI21_X1  g149(.A(new_n510), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g150(.A(new_n510), .B1(G868), .B2(G171), .ZN(G321));
  NOR2_X1   g151(.A1(G299), .A2(G868), .ZN(new_n513));
  AOI21_X1  g152(.A(new_n513), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g153(.A(new_n513), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g154(.A(new_n509), .ZN(new_n516));
  INV_X1    g155(.A(G559), .ZN(new_n517));
  OAI21_X1  g156(.A(new_n516), .B1(new_n517), .B2(G860), .ZN(G148));
  NOR2_X1   g157(.A1(new_n463), .A2(G868), .ZN(new_n519));
  NOR2_X1   g158(.A1(new_n509), .A2(G559), .ZN(new_n520));
  AOI21_X1  g159(.A(new_n519), .B1(G868), .B2(new_n520), .ZN(G323));
  XNOR2_X1  g160(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g161(.A1(new_n409), .A2(new_n405), .ZN(new_n523));
  XNOR2_X1  g162(.A(new_n523), .B(KEYINPUT12), .ZN(new_n524));
  XNOR2_X1  g163(.A(new_n524), .B(G2100), .ZN(new_n525));
  XNOR2_X1  g164(.A(new_n525), .B(KEYINPUT13), .ZN(new_n526));
  MUX2_X1   g165(.A(G135), .B(G123), .S(G2105), .Z(new_n527));
  NAND2_X1  g166(.A1(new_n527), .A2(new_n409), .ZN(new_n528));
  MUX2_X1   g167(.A(G99), .B(G111), .S(G2105), .Z(new_n529));
  NAND2_X1  g168(.A1(new_n529), .A2(G2104), .ZN(new_n530));
  NAND2_X1  g169(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  XOR2_X1   g170(.A(new_n531), .B(G2096), .Z(new_n532));
  NAND2_X1  g171(.A1(new_n526), .A2(new_n532), .ZN(G156));
  XOR2_X1   g172(.A(G2427), .B(G2430), .Z(new_n534));
  XNOR2_X1  g173(.A(new_n534), .B(KEYINPUT15), .ZN(new_n535));
  XNOR2_X1  g174(.A(G2435), .B(G2438), .ZN(new_n536));
  NAND3_X1  g175(.A1(new_n535), .A2(KEYINPUT14), .A3(new_n536), .ZN(new_n537));
  INV_X1    g176(.A(new_n536), .ZN(new_n538));
  NAND2_X1  g177(.A1(new_n538), .A2(KEYINPUT14), .ZN(new_n539));
  OAI21_X1  g178(.A(new_n537), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  XNOR2_X1  g179(.A(G2443), .B(G2446), .ZN(new_n541));
  XNOR2_X1  g180(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XNOR2_X1  g181(.A(G2451), .B(G2454), .ZN(new_n543));
  XNOR2_X1  g182(.A(new_n543), .B(KEYINPUT16), .ZN(new_n544));
  XOR2_X1   g183(.A(G1341), .B(G1348), .Z(new_n545));
  XOR2_X1   g184(.A(new_n544), .B(new_n545), .Z(new_n546));
  XNOR2_X1  g185(.A(new_n542), .B(new_n546), .ZN(new_n547));
  AND2_X1   g186(.A1(new_n547), .A2(G14), .ZN(G401));
  XOR2_X1   g187(.A(G2084), .B(G2090), .Z(new_n549));
  XNOR2_X1  g188(.A(G2072), .B(G2078), .ZN(new_n550));
  XNOR2_X1  g189(.A(G2067), .B(G2678), .ZN(new_n551));
  NAND3_X1  g190(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  XNOR2_X1  g191(.A(new_n552), .B(KEYINPUT18), .ZN(new_n553));
  XOR2_X1   g192(.A(new_n550), .B(KEYINPUT17), .Z(new_n554));
  INV_X1    g193(.A(new_n549), .ZN(new_n555));
  AND3_X1   g194(.A1(new_n554), .A2(new_n555), .A3(new_n551), .ZN(new_n556));
  MUX2_X1   g195(.A(new_n550), .B(new_n554), .S(new_n549), .Z(new_n557));
  INV_X1    g196(.A(new_n551), .ZN(new_n558));
  AOI211_X1 g197(.A(new_n553), .B(new_n556), .C1(new_n557), .C2(new_n558), .ZN(new_n559));
  XNOR2_X1  g198(.A(G2096), .B(G2100), .ZN(new_n560));
  XNOR2_X1  g199(.A(new_n559), .B(new_n560), .ZN(G227));
  XOR2_X1   g200(.A(G1971), .B(G1976), .Z(new_n562));
  XNOR2_X1  g201(.A(new_n562), .B(KEYINPUT19), .ZN(new_n563));
  XOR2_X1   g202(.A(G1961), .B(G1966), .Z(new_n564));
  NAND2_X1  g203(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g204(.A(G1956), .B(G2474), .ZN(new_n566));
  NOR2_X1   g205(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  XOR2_X1   g206(.A(new_n567), .B(KEYINPUT20), .Z(new_n568));
  NAND2_X1  g207(.A1(new_n565), .A2(new_n566), .ZN(new_n569));
  NOR2_X1   g208(.A1(new_n563), .A2(new_n564), .ZN(new_n570));
  XOR2_X1   g209(.A(new_n569), .B(new_n570), .Z(new_n571));
  NAND2_X1  g210(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g211(.A(G1981), .B(G1986), .ZN(new_n573));
  XNOR2_X1  g212(.A(new_n573), .B(KEYINPUT21), .ZN(new_n574));
  XOR2_X1   g213(.A(G1991), .B(G1996), .Z(new_n575));
  XNOR2_X1  g214(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XOR2_X1   g215(.A(new_n576), .B(KEYINPUT22), .Z(new_n577));
  XNOR2_X1  g216(.A(new_n572), .B(new_n577), .ZN(G229));
  NOR2_X1   g217(.A1(G4), .A2(G16), .ZN(new_n579));
  AOI21_X1  g218(.A(new_n579), .B1(new_n516), .B2(G16), .ZN(new_n580));
  XNOR2_X1  g219(.A(new_n580), .B(G1348), .ZN(new_n581));
  INV_X1    g220(.A(G16), .ZN(new_n582));
  NAND2_X1  g221(.A1(new_n582), .A2(G20), .ZN(new_n583));
  XNOR2_X1  g222(.A(new_n583), .B(KEYINPUT23), .ZN(new_n584));
  INV_X1    g223(.A(G299), .ZN(new_n585));
  OAI21_X1  g224(.A(new_n584), .B1(new_n585), .B2(new_n582), .ZN(new_n586));
  XNOR2_X1  g225(.A(new_n586), .B(G1956), .ZN(new_n587));
  NOR2_X1   g226(.A1(new_n581), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g227(.A1(G5), .A2(G16), .ZN(new_n589));
  AOI21_X1  g228(.A(new_n589), .B1(G171), .B2(G16), .ZN(new_n590));
  NAND2_X1  g229(.A1(new_n590), .A2(G1961), .ZN(new_n591));
  OR2_X1    g230(.A1(new_n590), .A2(G1961), .ZN(new_n592));
  INV_X1    g231(.A(G29), .ZN(new_n593));
  NAND2_X1  g232(.A1(new_n593), .A2(G26), .ZN(new_n594));
  XNOR2_X1  g233(.A(new_n594), .B(KEYINPUT28), .ZN(new_n595));
  MUX2_X1   g234(.A(G140), .B(G128), .S(G2105), .Z(new_n596));
  MUX2_X1   g235(.A(G104), .B(G116), .S(G2105), .Z(new_n597));
  AOI22_X1  g236(.A1(new_n409), .A2(new_n596), .B1(new_n597), .B2(G2104), .ZN(new_n598));
  OAI21_X1  g237(.A(new_n595), .B1(new_n598), .B2(new_n593), .ZN(new_n599));
  INV_X1    g238(.A(G2067), .ZN(new_n600));
  XNOR2_X1  g239(.A(new_n599), .B(new_n600), .ZN(new_n601));
  NAND4_X1  g240(.A1(new_n588), .A2(new_n591), .A3(new_n592), .A4(new_n601), .ZN(new_n602));
  NAND3_X1  g241(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n603));
  XOR2_X1   g242(.A(new_n603), .B(KEYINPUT26), .Z(new_n604));
  AND2_X1   g243(.A1(G129), .A2(G2105), .ZN(new_n605));
  AOI22_X1  g244(.A1(new_n409), .A2(new_n605), .B1(G105), .B2(new_n405), .ZN(new_n606));
  NAND3_X1  g245(.A1(new_n409), .A2(G141), .A3(new_n396), .ZN(new_n607));
  NAND3_X1  g246(.A1(new_n604), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  MUX2_X1   g247(.A(G32), .B(new_n608), .S(G29), .Z(new_n609));
  XNOR2_X1  g248(.A(new_n609), .B(G1996), .ZN(new_n610));
  XNOR2_X1  g249(.A(new_n610), .B(KEYINPUT27), .ZN(new_n611));
  NOR2_X1   g250(.A1(G29), .A2(G35), .ZN(new_n612));
  AOI21_X1  g251(.A(new_n612), .B1(G162), .B2(G29), .ZN(new_n613));
  XOR2_X1   g252(.A(new_n613), .B(KEYINPUT29), .Z(new_n614));
  INV_X1    g253(.A(G2090), .ZN(new_n615));
  NAND2_X1  g254(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OR2_X1    g255(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g256(.A1(new_n405), .A2(G103), .ZN(new_n618));
  INV_X1    g257(.A(KEYINPUT25), .ZN(new_n619));
  XNOR2_X1  g258(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND3_X1  g259(.A1(new_n409), .A2(G139), .A3(new_n396), .ZN(new_n621));
  AOI22_X1  g260(.A1(new_n409), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n622));
  OAI211_X1 g261(.A(new_n620), .B(new_n621), .C1(new_n396), .C2(new_n622), .ZN(new_n623));
  MUX2_X1   g262(.A(G33), .B(new_n623), .S(G29), .Z(new_n624));
  XOR2_X1   g263(.A(new_n624), .B(G2072), .Z(new_n625));
  NAND4_X1  g264(.A1(new_n611), .A2(new_n616), .A3(new_n617), .A4(new_n625), .ZN(new_n626));
  NOR2_X1   g265(.A1(G16), .A2(G19), .ZN(new_n627));
  AOI21_X1  g266(.A(new_n627), .B1(new_n464), .B2(G16), .ZN(new_n628));
  XOR2_X1   g267(.A(new_n628), .B(G1341), .Z(new_n629));
  OR2_X1    g268(.A1(KEYINPUT24), .A2(G34), .ZN(new_n630));
  NAND2_X1  g269(.A1(KEYINPUT24), .A2(G34), .ZN(new_n631));
  AOI21_X1  g270(.A(G29), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g271(.A(new_n632), .B1(G160), .B2(G29), .ZN(new_n633));
  XNOR2_X1  g272(.A(new_n633), .B(G2084), .ZN(new_n634));
  INV_X1    g273(.A(G1966), .ZN(new_n635));
  NAND2_X1  g274(.A1(G168), .A2(G16), .ZN(new_n636));
  OAI21_X1  g275(.A(new_n636), .B1(G16), .B2(G21), .ZN(new_n637));
  AOI21_X1  g276(.A(new_n634), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g277(.A1(new_n530), .A2(new_n528), .A3(G29), .ZN(new_n639));
  AND2_X1   g278(.A1(KEYINPUT30), .A2(G28), .ZN(new_n640));
  NOR2_X1   g279(.A1(KEYINPUT30), .A2(G28), .ZN(new_n641));
  OAI21_X1  g280(.A(new_n593), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g281(.A(KEYINPUT31), .ZN(new_n643));
  OR2_X1    g282(.A1(new_n643), .A2(G11), .ZN(new_n644));
  NAND2_X1  g283(.A1(new_n643), .A2(G11), .ZN(new_n645));
  NAND4_X1  g284(.A1(new_n639), .A2(new_n642), .A3(new_n644), .A4(new_n645), .ZN(new_n646));
  NOR2_X1   g285(.A1(G27), .A2(G29), .ZN(new_n647));
  AOI21_X1  g286(.A(new_n647), .B1(G164), .B2(G29), .ZN(new_n648));
  AOI21_X1  g287(.A(new_n646), .B1(new_n648), .B2(G2078), .ZN(new_n649));
  NAND3_X1  g288(.A1(new_n629), .A2(new_n638), .A3(new_n649), .ZN(new_n650));
  OAI22_X1  g289(.A1(new_n637), .A2(new_n635), .B1(new_n648), .B2(G2078), .ZN(new_n651));
  NOR4_X1   g290(.A1(new_n602), .A2(new_n626), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  INV_X1    g291(.A(new_n652), .ZN(new_n653));
  INV_X1    g292(.A(KEYINPUT36), .ZN(new_n654));
  NOR2_X1   g293(.A1(G6), .A2(G16), .ZN(new_n655));
  AOI21_X1  g294(.A(new_n655), .B1(new_n493), .B2(G16), .ZN(new_n656));
  XNOR2_X1  g295(.A(new_n656), .B(KEYINPUT32), .ZN(new_n657));
  INV_X1    g296(.A(G1981), .ZN(new_n658));
  XNOR2_X1  g297(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NOR2_X1   g298(.A1(G16), .A2(G23), .ZN(new_n660));
  NOR2_X1   g299(.A1(new_n485), .A2(new_n487), .ZN(new_n661));
  AOI21_X1  g300(.A(new_n660), .B1(new_n661), .B2(G16), .ZN(new_n662));
  XNOR2_X1  g301(.A(new_n662), .B(G1976), .ZN(new_n663));
  XNOR2_X1  g302(.A(new_n663), .B(KEYINPUT33), .ZN(new_n664));
  NOR2_X1   g303(.A1(G16), .A2(G22), .ZN(new_n665));
  AOI21_X1  g304(.A(new_n665), .B1(G166), .B2(G16), .ZN(new_n666));
  INV_X1    g305(.A(G1971), .ZN(new_n667));
  XNOR2_X1  g306(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NAND3_X1  g307(.A1(new_n659), .A2(new_n664), .A3(new_n668), .ZN(new_n669));
  OR2_X1    g308(.A1(new_n669), .A2(KEYINPUT34), .ZN(new_n670));
  MUX2_X1   g309(.A(G24), .B(G290), .S(G16), .Z(new_n671));
  OR2_X1    g310(.A1(new_n671), .A2(G1986), .ZN(new_n672));
  NAND2_X1  g311(.A1(new_n671), .A2(G1986), .ZN(new_n673));
  MUX2_X1   g312(.A(G131), .B(G119), .S(G2105), .Z(new_n674));
  NAND2_X1  g313(.A1(new_n674), .A2(new_n409), .ZN(new_n675));
  AND2_X1   g314(.A1(G107), .A2(G2105), .ZN(new_n676));
  AOI21_X1  g315(.A(new_n676), .B1(G95), .B2(new_n396), .ZN(new_n677));
  OAI21_X1  g316(.A(new_n675), .B1(new_n397), .B2(new_n677), .ZN(new_n678));
  MUX2_X1   g317(.A(G25), .B(new_n678), .S(G29), .Z(new_n679));
  XOR2_X1   g318(.A(KEYINPUT35), .B(G1991), .Z(new_n680));
  XNOR2_X1  g319(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND3_X1  g320(.A1(new_n672), .A2(new_n673), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g321(.A(new_n682), .B1(new_n669), .B2(KEYINPUT34), .ZN(new_n683));
  AOI21_X1  g322(.A(new_n654), .B1(new_n670), .B2(new_n683), .ZN(new_n684));
  INV_X1    g323(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g324(.A1(new_n670), .A2(new_n654), .A3(new_n683), .ZN(new_n686));
  AOI21_X1  g325(.A(new_n653), .B1(new_n685), .B2(new_n686), .ZN(G311));
  INV_X1    g326(.A(new_n686), .ZN(new_n688));
  OAI21_X1  g327(.A(new_n652), .B1(new_n688), .B2(new_n684), .ZN(G150));
  NOR2_X1   g328(.A1(new_n509), .A2(new_n517), .ZN(new_n690));
  XNOR2_X1  g329(.A(new_n690), .B(new_n463), .ZN(new_n691));
  XNOR2_X1  g330(.A(new_n691), .B(KEYINPUT38), .ZN(new_n692));
  AOI22_X1  g331(.A1(new_n428), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n693));
  NOR2_X1   g332(.A1(new_n693), .A2(new_n430), .ZN(new_n694));
  AOI22_X1  g333(.A1(new_n428), .A2(G93), .B1(G55), .B2(G543), .ZN(new_n695));
  NOR2_X1   g334(.A1(new_n695), .A2(new_n436), .ZN(new_n696));
  NOR2_X1   g335(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g336(.A(new_n692), .B(new_n697), .ZN(new_n698));
  INV_X1    g337(.A(KEYINPUT39), .ZN(new_n699));
  OR2_X1    g338(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g339(.A(G860), .ZN(new_n701));
  NAND2_X1  g340(.A1(new_n698), .A2(new_n699), .ZN(new_n702));
  NAND3_X1  g341(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NOR2_X1   g342(.A1(new_n697), .A2(new_n701), .ZN(new_n704));
  XNOR2_X1  g343(.A(new_n704), .B(KEYINPUT37), .ZN(new_n705));
  NAND2_X1  g344(.A1(new_n703), .A2(new_n705), .ZN(G145));
  NAND2_X1  g345(.A1(new_n420), .A2(new_n422), .ZN(new_n707));
  AND2_X1   g346(.A1(new_n416), .A2(new_n417), .ZN(new_n708));
  NAND2_X1  g347(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g348(.A(new_n623), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g349(.A(new_n608), .B(new_n598), .ZN(new_n711));
  XNOR2_X1  g350(.A(new_n710), .B(new_n711), .ZN(new_n712));
  MUX2_X1   g351(.A(G106), .B(G118), .S(G2105), .Z(new_n713));
  MUX2_X1   g352(.A(G142), .B(G130), .S(G2105), .Z(new_n714));
  AOI22_X1  g353(.A1(G2104), .A2(new_n713), .B1(new_n714), .B2(new_n409), .ZN(new_n715));
  XOR2_X1   g354(.A(new_n678), .B(new_n715), .Z(new_n716));
  XNOR2_X1  g355(.A(new_n712), .B(new_n716), .ZN(new_n717));
  XNOR2_X1  g356(.A(new_n524), .B(new_n531), .ZN(new_n718));
  XNOR2_X1  g357(.A(G160), .B(G162), .ZN(new_n719));
  XNOR2_X1  g358(.A(new_n718), .B(new_n719), .ZN(new_n720));
  XNOR2_X1  g359(.A(new_n717), .B(new_n720), .ZN(new_n721));
  INV_X1    g360(.A(G37), .ZN(new_n722));
  NAND2_X1  g361(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g362(.A(new_n723), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g363(.A(new_n493), .B(G290), .Z(new_n725));
  XNOR2_X1  g364(.A(G166), .B(new_n661), .ZN(new_n726));
  XNOR2_X1  g365(.A(new_n725), .B(new_n726), .ZN(new_n727));
  INV_X1    g366(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g367(.A1(new_n509), .A2(new_n585), .ZN(new_n729));
  NAND3_X1  g368(.A1(new_n503), .A2(G299), .A3(new_n508), .ZN(new_n730));
  NAND2_X1  g369(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g370(.A(KEYINPUT41), .ZN(new_n732));
  NAND2_X1  g371(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g372(.A(new_n463), .B(new_n697), .ZN(new_n734));
  NAND3_X1  g373(.A1(new_n729), .A2(new_n730), .A3(KEYINPUT41), .ZN(new_n735));
  NAND3_X1  g374(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  INV_X1    g375(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g376(.A1(new_n734), .A2(new_n731), .ZN(new_n738));
  OAI22_X1  g377(.A1(new_n737), .A2(new_n738), .B1(G559), .B2(new_n509), .ZN(new_n739));
  INV_X1    g378(.A(KEYINPUT42), .ZN(new_n740));
  INV_X1    g379(.A(new_n735), .ZN(new_n741));
  AOI21_X1  g380(.A(KEYINPUT41), .B1(new_n729), .B2(new_n730), .ZN(new_n742));
  NOR3_X1   g381(.A1(new_n741), .A2(new_n734), .A3(new_n742), .ZN(new_n743));
  INV_X1    g382(.A(new_n731), .ZN(new_n744));
  NAND2_X1  g383(.A1(new_n744), .A2(new_n734), .ZN(new_n745));
  INV_X1    g384(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g385(.A(new_n520), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  AND3_X1   g386(.A1(new_n739), .A2(new_n740), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g387(.A(new_n740), .B1(new_n739), .B2(new_n747), .ZN(new_n749));
  OAI21_X1  g388(.A(new_n728), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g389(.A1(new_n750), .A2(G868), .ZN(new_n751));
  NOR3_X1   g390(.A1(new_n748), .A2(new_n749), .A3(new_n728), .ZN(new_n752));
  OAI22_X1  g391(.A1(new_n751), .A2(new_n752), .B1(G868), .B2(new_n697), .ZN(G295));
  OAI22_X1  g392(.A1(new_n751), .A2(new_n752), .B1(G868), .B2(new_n697), .ZN(G331));
  XNOR2_X1  g393(.A(G168), .B(G171), .ZN(new_n755));
  INV_X1    g394(.A(new_n738), .ZN(new_n756));
  AOI21_X1  g395(.A(new_n755), .B1(new_n756), .B2(new_n736), .ZN(new_n757));
  INV_X1    g396(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g397(.A(new_n755), .B1(new_n743), .B2(new_n746), .ZN(new_n759));
  NAND3_X1  g398(.A1(new_n758), .A2(new_n728), .A3(new_n759), .ZN(new_n760));
  INV_X1    g399(.A(new_n755), .ZN(new_n761));
  INV_X1    g400(.A(new_n734), .ZN(new_n762));
  NAND3_X1  g401(.A1(new_n762), .A2(new_n733), .A3(new_n735), .ZN(new_n763));
  AOI21_X1  g402(.A(new_n761), .B1(new_n763), .B2(new_n745), .ZN(new_n764));
  OAI21_X1  g403(.A(new_n727), .B1(new_n764), .B2(new_n757), .ZN(new_n765));
  NAND3_X1  g404(.A1(new_n760), .A2(new_n765), .A3(new_n722), .ZN(new_n766));
  NAND2_X1  g405(.A1(new_n766), .A2(KEYINPUT43), .ZN(new_n767));
  INV_X1    g406(.A(KEYINPUT44), .ZN(new_n768));
  INV_X1    g407(.A(KEYINPUT43), .ZN(new_n769));
  NAND4_X1  g408(.A1(new_n760), .A2(new_n765), .A3(new_n769), .A4(new_n722), .ZN(new_n770));
  AND3_X1   g409(.A1(new_n767), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g410(.A(new_n768), .B1(new_n767), .B2(new_n770), .ZN(new_n772));
  NOR2_X1   g411(.A1(new_n771), .A2(new_n772), .ZN(G397));
  INV_X1    g412(.A(G40), .ZN(new_n774));
  NOR3_X1   g413(.A1(new_n403), .A2(new_n407), .A3(new_n774), .ZN(new_n775));
  INV_X1    g414(.A(G1384), .ZN(new_n776));
  AOI21_X1  g415(.A(KEYINPUT45), .B1(new_n709), .B2(new_n776), .ZN(new_n777));
  INV_X1    g416(.A(KEYINPUT45), .ZN(new_n778));
  AOI211_X1 g417(.A(new_n778), .B(G1384), .C1(new_n707), .C2(new_n708), .ZN(new_n779));
  OAI21_X1  g418(.A(new_n775), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  INV_X1    g419(.A(new_n780), .ZN(new_n781));
  NAND3_X1  g420(.A1(new_n775), .A2(new_n709), .A3(new_n776), .ZN(new_n782));
  NAND3_X1  g421(.A1(new_n781), .A2(new_n600), .A3(new_n782), .ZN(new_n783));
  INV_X1    g422(.A(new_n782), .ZN(new_n784));
  NOR3_X1   g423(.A1(new_n780), .A2(new_n598), .A3(new_n784), .ZN(new_n785));
  NOR2_X1   g424(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  INV_X1    g425(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g426(.A1(new_n781), .A2(new_n608), .A3(new_n782), .ZN(new_n788));
  NOR3_X1   g427(.A1(new_n780), .A2(G1996), .A3(new_n784), .ZN(new_n789));
  OR2_X1    g428(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g429(.A1(new_n783), .A2(new_n785), .ZN(new_n791));
  NAND2_X1  g430(.A1(new_n788), .A2(new_n789), .ZN(new_n792));
  AND4_X1   g431(.A1(new_n787), .A2(new_n790), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  NAND3_X1  g432(.A1(new_n781), .A2(new_n678), .A3(new_n782), .ZN(new_n794));
  AND4_X1   g433(.A1(new_n680), .A2(new_n794), .A3(new_n782), .A4(new_n781), .ZN(new_n795));
  AOI21_X1  g434(.A(new_n786), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  NAND3_X1  g435(.A1(new_n781), .A2(new_n680), .A3(new_n782), .ZN(new_n797));
  XNOR2_X1  g436(.A(new_n797), .B(new_n794), .ZN(new_n798));
  NAND3_X1  g437(.A1(new_n781), .A2(G290), .A3(new_n782), .ZN(new_n799));
  NOR3_X1   g438(.A1(new_n780), .A2(G1986), .A3(new_n784), .ZN(new_n800));
  NAND2_X1  g439(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g440(.A(new_n801), .B(KEYINPUT48), .ZN(new_n802));
  NAND3_X1  g441(.A1(new_n793), .A2(new_n798), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g442(.A1(new_n796), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g443(.A1(new_n787), .A2(new_n791), .A3(new_n788), .ZN(new_n805));
  XNOR2_X1  g444(.A(new_n789), .B(KEYINPUT46), .ZN(new_n806));
  OAI21_X1  g445(.A(KEYINPUT47), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OR3_X1    g446(.A1(new_n805), .A2(KEYINPUT47), .A3(new_n806), .ZN(new_n808));
  AOI21_X1  g447(.A(new_n804), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g448(.A(new_n778), .B1(G164), .B2(G1384), .ZN(new_n810));
  NAND3_X1  g449(.A1(new_n709), .A2(KEYINPUT45), .A3(new_n776), .ZN(new_n811));
  NAND3_X1  g450(.A1(new_n810), .A2(new_n811), .A3(new_n775), .ZN(new_n812));
  NAND2_X1  g451(.A1(new_n812), .A2(new_n667), .ZN(new_n813));
  INV_X1    g452(.A(KEYINPUT50), .ZN(new_n814));
  OAI21_X1  g453(.A(new_n814), .B1(G164), .B2(G1384), .ZN(new_n815));
  NAND3_X1  g454(.A1(new_n709), .A2(KEYINPUT50), .A3(new_n776), .ZN(new_n816));
  NAND2_X1  g455(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g456(.A1(new_n817), .A2(new_n775), .ZN(new_n818));
  OAI21_X1  g457(.A(new_n813), .B1(new_n818), .B2(G2090), .ZN(new_n819));
  AOI21_X1  g458(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n820));
  NAND3_X1  g459(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n821));
  INV_X1    g460(.A(new_n821), .ZN(new_n822));
  OAI211_X1 g461(.A(new_n819), .B(G8), .C1(new_n820), .C2(new_n822), .ZN(new_n823));
  AND2_X1   g462(.A1(new_n782), .A2(G8), .ZN(new_n824));
  INV_X1    g463(.A(KEYINPUT52), .ZN(new_n825));
  NOR2_X1   g464(.A1(G288), .A2(G1976), .ZN(new_n826));
  INV_X1    g465(.A(G1976), .ZN(new_n827));
  NOR2_X1   g466(.A1(new_n661), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g467(.A(new_n824), .B(new_n825), .C1(new_n826), .C2(new_n828), .ZN(new_n829));
  XOR2_X1   g468(.A(KEYINPUT49), .B(G1981), .Z(new_n830));
  NAND2_X1  g469(.A1(new_n493), .A2(new_n830), .ZN(new_n831));
  INV_X1    g470(.A(new_n830), .ZN(new_n832));
  OAI21_X1  g471(.A(new_n832), .B1(new_n490), .B2(new_n492), .ZN(new_n833));
  NAND2_X1  g472(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g473(.A1(new_n834), .A2(new_n824), .ZN(new_n835));
  NAND2_X1  g474(.A1(new_n782), .A2(G8), .ZN(new_n836));
  AOI21_X1  g475(.A(new_n836), .B1(G1976), .B2(new_n661), .ZN(new_n837));
  OAI211_X1 g476(.A(new_n829), .B(new_n835), .C1(new_n825), .C2(new_n837), .ZN(new_n838));
  NOR2_X1   g477(.A1(new_n823), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g478(.A1(new_n826), .A2(new_n833), .A3(new_n831), .ZN(new_n840));
  NAND2_X1  g479(.A1(new_n493), .A2(new_n658), .ZN(new_n841));
  AOI21_X1  g480(.A(new_n836), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g481(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g482(.A1(new_n819), .A2(G8), .ZN(new_n844));
  NOR2_X1   g483(.A1(new_n822), .A2(new_n820), .ZN(new_n845));
  NAND2_X1  g484(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AND2_X1   g485(.A1(new_n846), .A2(new_n823), .ZN(new_n847));
  NAND2_X1  g486(.A1(new_n812), .A2(new_n635), .ZN(new_n848));
  INV_X1    g487(.A(G2084), .ZN(new_n849));
  NOR3_X1   g488(.A1(G164), .A2(new_n814), .A3(G1384), .ZN(new_n850));
  AOI21_X1  g489(.A(KEYINPUT50), .B1(new_n709), .B2(new_n776), .ZN(new_n851));
  OAI211_X1 g490(.A(new_n849), .B(new_n775), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NAND2_X1  g491(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g492(.A1(new_n853), .A2(G8), .A3(G168), .ZN(new_n854));
  NOR2_X1   g493(.A1(new_n838), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g494(.A(KEYINPUT63), .B1(new_n847), .B2(new_n855), .ZN(new_n856));
  AND4_X1   g495(.A1(KEYINPUT63), .A2(new_n855), .A3(new_n823), .A4(new_n846), .ZN(new_n857));
  OAI21_X1  g496(.A(new_n843), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g497(.A(G8), .ZN(new_n859));
  AOI21_X1  g498(.A(new_n859), .B1(new_n848), .B2(new_n852), .ZN(new_n860));
  NOR2_X1   g499(.A1(G168), .A2(new_n859), .ZN(new_n861));
  NOR3_X1   g500(.A1(new_n860), .A2(KEYINPUT51), .A3(new_n861), .ZN(new_n862));
  INV_X1    g501(.A(new_n862), .ZN(new_n863));
  NAND4_X1  g502(.A1(new_n848), .A2(new_n852), .A3(G8), .A4(G286), .ZN(new_n864));
  AND2_X1   g503(.A1(new_n854), .A2(new_n864), .ZN(new_n865));
  INV_X1    g504(.A(KEYINPUT51), .ZN(new_n866));
  OAI211_X1 g505(.A(new_n863), .B(KEYINPUT62), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  INV_X1    g506(.A(G1961), .ZN(new_n868));
  NAND2_X1  g507(.A1(new_n818), .A2(new_n868), .ZN(new_n869));
  INV_X1    g508(.A(G2078), .ZN(new_n870));
  NAND4_X1  g509(.A1(new_n810), .A2(new_n811), .A3(new_n870), .A4(new_n775), .ZN(new_n871));
  AND2_X1   g510(.A1(new_n871), .A2(KEYINPUT53), .ZN(new_n872));
  NOR2_X1   g511(.A1(new_n871), .A2(KEYINPUT53), .ZN(new_n873));
  OAI21_X1  g512(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g513(.A1(new_n874), .A2(G171), .ZN(new_n875));
  NOR2_X1   g514(.A1(new_n875), .A2(new_n838), .ZN(new_n876));
  INV_X1    g515(.A(KEYINPUT62), .ZN(new_n877));
  AOI21_X1  g516(.A(new_n866), .B1(new_n854), .B2(new_n864), .ZN(new_n878));
  OAI21_X1  g517(.A(new_n877), .B1(new_n878), .B2(new_n862), .ZN(new_n879));
  NAND3_X1  g518(.A1(new_n867), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  XNOR2_X1  g519(.A(G299), .B(KEYINPUT57), .ZN(new_n881));
  AOI21_X1  g520(.A(G1956), .B1(new_n817), .B2(new_n775), .ZN(new_n882));
  XNOR2_X1  g521(.A(KEYINPUT56), .B(G2072), .ZN(new_n883));
  AND4_X1   g522(.A1(new_n775), .A2(new_n810), .A3(new_n811), .A4(new_n883), .ZN(new_n884));
  OAI21_X1  g523(.A(new_n881), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  XOR2_X1   g524(.A(G299), .B(KEYINPUT57), .Z(new_n886));
  NAND4_X1  g525(.A1(new_n810), .A2(new_n811), .A3(new_n775), .A4(new_n883), .ZN(new_n887));
  INV_X1    g526(.A(new_n775), .ZN(new_n888));
  AOI21_X1  g527(.A(new_n888), .B1(new_n815), .B2(new_n816), .ZN(new_n889));
  OAI211_X1 g528(.A(new_n886), .B(new_n887), .C1(G1956), .C2(new_n889), .ZN(new_n890));
  OAI22_X1  g529(.A1(new_n889), .A2(G1348), .B1(G2067), .B2(new_n782), .ZN(new_n891));
  NAND4_X1  g530(.A1(new_n885), .A2(new_n890), .A3(new_n516), .A4(new_n891), .ZN(new_n892));
  NAND2_X1  g531(.A1(new_n892), .A2(new_n885), .ZN(new_n893));
  AND3_X1   g532(.A1(new_n885), .A2(KEYINPUT61), .A3(new_n890), .ZN(new_n894));
  AOI21_X1  g533(.A(KEYINPUT61), .B1(new_n885), .B2(new_n890), .ZN(new_n895));
  INV_X1    g534(.A(KEYINPUT59), .ZN(new_n896));
  INV_X1    g535(.A(G1996), .ZN(new_n897));
  NAND4_X1  g536(.A1(new_n810), .A2(new_n811), .A3(new_n897), .A4(new_n775), .ZN(new_n898));
  XOR2_X1   g537(.A(KEYINPUT58), .B(G1341), .Z(new_n899));
  NAND2_X1  g538(.A1(new_n782), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g539(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g540(.A(new_n896), .B1(new_n901), .B2(new_n464), .ZN(new_n902));
  AOI211_X1 g541(.A(KEYINPUT59), .B(new_n463), .C1(new_n898), .C2(new_n900), .ZN(new_n903));
  NOR2_X1   g542(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NOR3_X1   g543(.A1(new_n894), .A2(new_n895), .A3(new_n904), .ZN(new_n905));
  NOR3_X1   g544(.A1(new_n891), .A2(KEYINPUT60), .A3(new_n509), .ZN(new_n906));
  XNOR2_X1  g545(.A(new_n891), .B(new_n516), .ZN(new_n907));
  AOI21_X1  g546(.A(new_n906), .B1(new_n907), .B2(KEYINPUT60), .ZN(new_n908));
  AOI21_X1  g547(.A(new_n893), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  NOR2_X1   g548(.A1(new_n878), .A2(new_n862), .ZN(new_n910));
  INV_X1    g549(.A(KEYINPUT54), .ZN(new_n911));
  NOR2_X1   g550(.A1(new_n777), .A2(new_n779), .ZN(new_n912));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n913));
  NAND4_X1  g552(.A1(new_n912), .A2(new_n913), .A3(new_n870), .A4(new_n775), .ZN(new_n914));
  NAND2_X1  g553(.A1(new_n871), .A2(KEYINPUT53), .ZN(new_n915));
  AOI221_X4 g554(.A(G171), .B1(new_n818), .B2(new_n868), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  NAND2_X1  g555(.A1(new_n914), .A2(new_n915), .ZN(new_n917));
  AOI21_X1  g556(.A(G301), .B1(new_n917), .B2(new_n869), .ZN(new_n918));
  OAI21_X1  g557(.A(new_n911), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g558(.A1(new_n917), .A2(G301), .A3(new_n869), .ZN(new_n920));
  NAND3_X1  g559(.A1(new_n875), .A2(new_n920), .A3(KEYINPUT54), .ZN(new_n921));
  INV_X1    g560(.A(new_n838), .ZN(new_n922));
  NAND4_X1  g561(.A1(new_n910), .A2(new_n919), .A3(new_n921), .A4(new_n922), .ZN(new_n923));
  OAI21_X1  g562(.A(new_n880), .B1(new_n909), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g563(.A(new_n858), .B1(new_n924), .B2(new_n847), .ZN(new_n925));
  OR2_X1    g564(.A1(new_n799), .A2(new_n800), .ZN(new_n926));
  NAND4_X1  g565(.A1(new_n793), .A2(new_n798), .A3(new_n801), .A4(new_n926), .ZN(new_n927));
  OAI21_X1  g566(.A(new_n809), .B1(new_n925), .B2(new_n927), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g567(.A1(new_n767), .A2(new_n770), .ZN(new_n930));
  NOR4_X1   g568(.A1(G401), .A2(G229), .A3(new_n394), .A4(G227), .ZN(new_n931));
  NAND3_X1  g569(.A1(new_n930), .A2(new_n723), .A3(new_n931), .ZN(G225));
  INV_X1    g570(.A(G225), .ZN(G308));
endmodule


