//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n553, new_n554, new_n555, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n611,
    new_n612, new_n614, new_n615, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192, new_n1193, new_n1194;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT67), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  OR4_X1    g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  AND2_X1   g033(.A1(new_n458), .A2(KEYINPUT68), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n454), .A2(G567), .ZN(new_n460));
  OAI21_X1  g035(.A(new_n460), .B1(new_n458), .B2(KEYINPUT68), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  XOR2_X1   g037(.A(new_n462), .B(KEYINPUT69), .Z(G319));
  INV_X1    g038(.A(KEYINPUT70), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n470), .A2(KEYINPUT70), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n467), .A2(new_n472), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n469), .A2(G2105), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n477), .A2(G137), .B1(G101), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n482), .B1(new_n470), .B2(new_n471), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n482), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n487), .B1(G136), .B2(new_n477), .ZN(new_n488));
  XNOR2_X1  g063(.A(new_n488), .B(KEYINPUT71), .ZN(G162));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  AND3_X1   g065(.A1(new_n490), .A2(new_n482), .A3(G138), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n467), .A2(new_n472), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(KEYINPUT73), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT73), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n467), .A2(new_n472), .A3(new_n494), .A4(new_n491), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n490), .B1(new_n477), .B2(G138), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  OR2_X1    g074(.A1(G102), .A2(G2105), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n500), .B(G2104), .C1(G114), .C2(new_n482), .ZN(new_n501));
  OAI211_X1 g076(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT72), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT72), .B1(new_n501), .B2(new_n502), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n499), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XOR2_X1   g087(.A(KEYINPUT5), .B(G543), .Z(new_n513));
  AND2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  XOR2_X1   g092(.A(KEYINPUT74), .B(G88), .Z(new_n518));
  INV_X1    g093(.A(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n517), .A2(new_n518), .B1(new_n520), .B2(G50), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n512), .A2(new_n521), .ZN(G166));
  NAND2_X1  g097(.A1(new_n513), .A2(KEYINPUT75), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT75), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n509), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G63), .ZN(new_n527));
  NOR3_X1   g102(.A1(new_n526), .A2(new_n527), .A3(new_n511), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n520), .A2(G51), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  INV_X1    g106(.A(G89), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n509), .B1(new_n515), .B2(new_n514), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n529), .B(new_n531), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n528), .A2(new_n534), .ZN(G168));
  NAND3_X1  g110(.A1(new_n523), .A2(G64), .A3(new_n525), .ZN(new_n536));
  NAND2_X1  g111(.A1(G77), .A2(G543), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n511), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n517), .A2(G90), .B1(new_n520), .B2(G52), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n538), .A2(new_n540), .ZN(G171));
  OR2_X1    g116(.A1(new_n514), .A2(new_n515), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n543), .A2(new_n544), .B1(new_n533), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(G68), .A2(G543), .ZN(new_n547));
  INV_X1    g122(.A(G56), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n526), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n546), .B1(new_n549), .B2(G651), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT76), .ZN(G188));
  NAND2_X1  g131(.A1(new_n520), .A2(G53), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT77), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n513), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n562), .A2(G651), .B1(new_n517), .B2(G91), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n558), .A2(new_n563), .ZN(G299));
  OAI21_X1  g139(.A(KEYINPUT78), .B1(new_n538), .B2(new_n540), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NOR3_X1   g141(.A1(new_n538), .A2(new_n540), .A3(KEYINPUT78), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n566), .A2(new_n567), .ZN(G301));
  INV_X1    g143(.A(G168), .ZN(G286));
  OAI21_X1  g144(.A(new_n521), .B1(new_n511), .B2(new_n510), .ZN(G303));
  NAND3_X1  g145(.A1(new_n542), .A2(G49), .A3(G543), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT79), .ZN(new_n572));
  INV_X1    g147(.A(G74), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n509), .A2(new_n524), .ZN(new_n574));
  OR2_X1    g149(.A1(KEYINPUT5), .A2(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(KEYINPUT5), .A2(G543), .ZN(new_n576));
  AOI21_X1  g151(.A(KEYINPUT75), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n573), .B1(new_n574), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(G651), .B1(G87), .B2(new_n517), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n572), .A2(new_n579), .ZN(G288));
  INV_X1    g155(.A(G86), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT80), .B1(new_n533), .B2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT80), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n542), .A2(new_n583), .A3(G86), .A4(new_n509), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(G73), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n513), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(new_n520), .B2(G48), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n585), .A2(new_n589), .ZN(G305));
  AOI22_X1  g165(.A1(new_n517), .A2(G85), .B1(new_n520), .B2(G47), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT81), .ZN(new_n592));
  NAND2_X1  g167(.A1(G72), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G60), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n526), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(G290));
  AND3_X1   g172(.A1(new_n542), .A2(G92), .A3(new_n509), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT10), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n513), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(new_n520), .B2(G54), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n604), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G301), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G284));
  AOI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G321));
  MUX2_X1   g183(.A(G299), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g184(.A(G299), .B(G286), .S(G868), .Z(G280));
  INV_X1    g185(.A(new_n604), .ZN(new_n611));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G860), .ZN(G148));
  NAND2_X1  g188(.A1(new_n611), .A2(new_n612), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g191(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n617));
  XNOR2_X1  g192(.A(G323), .B(new_n617), .ZN(G282));
  AND2_X1   g193(.A1(new_n467), .A2(new_n472), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(new_n478), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT12), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  INV_X1    g197(.A(G2100), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n477), .A2(G135), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n483), .A2(G123), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n482), .A2(G111), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n626), .B(new_n627), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(KEYINPUT83), .B(G2096), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n624), .A2(new_n625), .A3(new_n632), .ZN(G156));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n637), .A2(KEYINPUT14), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2451), .B(G2454), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT16), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n639), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2443), .B(G2446), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G1341), .B(G1348), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT84), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n644), .A2(new_n645), .ZN(new_n648));
  AND2_X1   g223(.A1(new_n648), .A2(G14), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n650), .A2(KEYINPUT85), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(KEYINPUT85), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT86), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2072), .B(G2078), .Z(new_n659));
  NOR3_X1   g234(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT18), .ZN(new_n661));
  XOR2_X1   g236(.A(KEYINPUT88), .B(KEYINPUT17), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n663), .A2(new_n657), .A3(new_n656), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n657), .B1(new_n656), .B2(new_n659), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT87), .ZN(new_n666));
  OAI22_X1  g241(.A1(new_n665), .A2(new_n666), .B1(new_n663), .B2(new_n656), .ZN(new_n667));
  INV_X1    g242(.A(new_n665), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n668), .A2(KEYINPUT87), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n661), .B(new_n664), .C1(new_n667), .C2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2096), .B(G2100), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT20), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n676), .B(new_n677), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n680), .B(new_n681), .C1(new_n675), .C2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT90), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n685), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n688), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(G229));
  XOR2_X1   g267(.A(KEYINPUT91), .B(G29), .Z(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n694), .A2(G35), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n695), .B1(G162), .B2(new_n694), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT29), .Z(new_n697));
  INV_X1    g272(.A(G2090), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G20), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT23), .Z(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(G299), .B2(G16), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1956), .ZN(new_n704));
  NAND2_X1  g279(.A1(G160), .A2(G29), .ZN(new_n705));
  INV_X1    g280(.A(KEYINPUT24), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n706), .A2(G34), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(G34), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n693), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n705), .A2(G2084), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n700), .A2(G5), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G171), .B2(new_n700), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(G1961), .ZN(new_n713));
  NOR2_X1   g288(.A1(G16), .A2(G19), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n550), .B2(G16), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n715), .A2(G1341), .ZN(new_n716));
  NAND4_X1  g291(.A1(new_n704), .A2(new_n710), .A3(new_n713), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n700), .A2(G21), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G168), .B2(new_n700), .ZN(new_n719));
  INV_X1    g294(.A(G1966), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n693), .A2(G26), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT28), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n477), .A2(G140), .ZN(new_n724));
  INV_X1    g299(.A(KEYINPUT94), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n727));
  INV_X1    g302(.A(G116), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(G2105), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(new_n483), .B2(G128), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n723), .B1(new_n731), .B2(G29), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(G2067), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n715), .A2(G1341), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n712), .A2(G1961), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n721), .A2(new_n733), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(G2084), .B1(new_n705), .B2(new_n709), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT98), .Z(new_n738));
  NOR4_X1   g313(.A1(new_n699), .A2(new_n717), .A3(new_n736), .A4(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n700), .A2(G4), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(new_n611), .B2(new_n700), .ZN(new_n741));
  INV_X1    g316(.A(G1348), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT30), .B(G28), .ZN(new_n744));
  INV_X1    g319(.A(G29), .ZN(new_n745));
  OR2_X1    g320(.A1(KEYINPUT31), .A2(G11), .ZN(new_n746));
  NAND2_X1  g321(.A1(KEYINPUT31), .A2(G11), .ZN(new_n747));
  AOI22_X1  g322(.A1(new_n744), .A2(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n630), .B2(new_n693), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT97), .B(KEYINPUT26), .Z(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n478), .A2(G105), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n483), .A2(G129), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n477), .A2(G141), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n758), .A2(new_n745), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n745), .B2(G32), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT27), .B(G1996), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n749), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n743), .B(new_n762), .C1(new_n760), .C2(new_n761), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n507), .A2(new_n694), .ZN(new_n764));
  INV_X1    g339(.A(G2078), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n693), .A2(G27), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT99), .ZN(new_n767));
  AND3_X1   g342(.A1(new_n764), .A2(new_n765), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n765), .B1(new_n764), .B2(new_n767), .ZN(new_n769));
  NOR3_X1   g344(.A1(new_n763), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n739), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n697), .A2(new_n698), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT100), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT96), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n619), .A2(G127), .ZN(new_n775));
  NAND2_X1  g350(.A1(G115), .A2(G2104), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n482), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT95), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT25), .ZN(new_n781));
  NAND2_X1  g356(.A1(G103), .A2(G2104), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(G2105), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n482), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n477), .A2(G139), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n777), .B2(new_n778), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n774), .B1(new_n780), .B2(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n777), .A2(new_n778), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n788), .A2(new_n779), .A3(KEYINPUT96), .A4(new_n785), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  MUX2_X1   g365(.A(G33), .B(new_n790), .S(G29), .Z(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(G2072), .Z(new_n792));
  NAND3_X1  g367(.A1(new_n771), .A2(new_n773), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n700), .A2(G6), .ZN(new_n794));
  INV_X1    g369(.A(G305), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n700), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT32), .B(G1981), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n572), .A2(new_n579), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(new_n700), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(new_n700), .B2(G23), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT33), .B(G1976), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n798), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n700), .A2(G22), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT93), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G166), .B2(new_n700), .ZN(new_n806));
  INV_X1    g381(.A(G1971), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n803), .B(new_n808), .C1(new_n801), .C2(new_n802), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT34), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n700), .A2(G24), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n592), .A2(new_n596), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(new_n700), .ZN(new_n813));
  INV_X1    g388(.A(G1986), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(KEYINPUT92), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(KEYINPUT92), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n477), .A2(G131), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n483), .A2(G119), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n482), .A2(G107), .ZN(new_n820));
  OAI21_X1  g395(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n818), .B(new_n819), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  MUX2_X1   g397(.A(G25), .B(new_n822), .S(new_n694), .Z(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT35), .B(G1991), .ZN(new_n824));
  XOR2_X1   g399(.A(new_n823), .B(new_n824), .Z(new_n825));
  NAND3_X1  g400(.A1(new_n816), .A2(new_n817), .A3(new_n825), .ZN(new_n826));
  OR3_X1    g401(.A1(new_n810), .A2(KEYINPUT36), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(KEYINPUT36), .B1(new_n810), .B2(new_n826), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n793), .B1(new_n827), .B2(new_n828), .ZN(G311));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n830), .A2(new_n771), .A3(new_n773), .A4(new_n792), .ZN(G150));
  NAND3_X1  g406(.A1(new_n523), .A2(G67), .A3(new_n525), .ZN(new_n832));
  NAND2_X1  g407(.A1(G80), .A2(G543), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n511), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(G55), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT101), .B(G93), .Z(new_n836));
  OAI22_X1  g411(.A1(new_n543), .A2(new_n835), .B1(new_n533), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(KEYINPUT102), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n834), .A2(KEYINPUT102), .A3(new_n837), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(G860), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT104), .Z(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT37), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n604), .A2(new_n612), .ZN(new_n846));
  XOR2_X1   g421(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  AND2_X1   g423(.A1(new_n549), .A2(G651), .ZN(new_n849));
  OAI22_X1  g424(.A1(new_n839), .A2(new_n840), .B1(new_n849), .B2(new_n546), .ZN(new_n850));
  NOR2_X1   g425(.A1(new_n834), .A2(new_n837), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n550), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n848), .B(new_n853), .Z(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n855), .A2(KEYINPUT39), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n842), .B1(new_n855), .B2(KEYINPUT39), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n845), .B1(new_n856), .B2(new_n857), .ZN(G145));
  NAND2_X1  g433(.A1(new_n477), .A2(G142), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n483), .A2(G130), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n482), .A2(G118), .ZN(new_n861));
  OAI21_X1  g436(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n859), .B(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT106), .Z(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(new_n621), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n621), .ZN(new_n866));
  AND3_X1   g441(.A1(new_n865), .A2(new_n866), .A3(new_n822), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n822), .B1(new_n865), .B2(new_n866), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n790), .A2(KEYINPUT105), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT105), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n787), .A2(new_n789), .A3(new_n871), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n758), .A2(new_n731), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n501), .A2(new_n502), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n758), .A2(new_n731), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n873), .A2(new_n499), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n873), .A2(new_n876), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n499), .A2(new_n875), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n870), .A2(new_n872), .A3(new_n877), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n877), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n882), .A2(KEYINPUT105), .A3(new_n790), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n869), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n480), .B(new_n630), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n886), .B(G162), .Z(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n883), .A2(new_n881), .A3(new_n869), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n885), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n889), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n887), .B1(new_n891), .B2(new_n884), .ZN(new_n892));
  INV_X1    g467(.A(G37), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n890), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(KEYINPUT107), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT107), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n890), .A2(new_n892), .A3(new_n896), .A4(new_n893), .ZN(new_n897));
  AND3_X1   g472(.A1(new_n895), .A2(KEYINPUT40), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT40), .B1(new_n895), .B2(new_n897), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(G395));
  NAND2_X1  g475(.A1(new_n812), .A2(G288), .ZN(new_n901));
  NAND2_X1  g476(.A1(G166), .A2(KEYINPUT108), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT108), .ZN(new_n903));
  NAND2_X1  g478(.A1(G303), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(new_n795), .ZN(new_n906));
  NAND2_X1  g481(.A1(G290), .A2(new_n799), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n902), .A2(G305), .A3(new_n904), .ZN(new_n908));
  AND4_X1   g483(.A1(new_n901), .A2(new_n906), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  AOI22_X1  g484(.A1(new_n901), .A2(new_n907), .B1(new_n906), .B2(new_n908), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT42), .ZN(new_n912));
  XNOR2_X1  g487(.A(new_n853), .B(new_n614), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n604), .A2(G299), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n599), .A2(new_n558), .A3(new_n563), .A4(new_n603), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n915), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n599), .A2(new_n603), .B1(new_n558), .B2(new_n563), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT41), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT41), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n914), .A2(new_n921), .A3(new_n915), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n917), .B1(new_n923), .B2(new_n913), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n912), .B(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(G868), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n926), .B1(G868), .B2(new_n841), .ZN(G295));
  OAI21_X1  g502(.A(new_n926), .B1(G868), .B2(new_n841), .ZN(G331));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT113), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT78), .ZN(new_n931));
  NAND2_X1  g506(.A1(G171), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(G286), .B1(new_n932), .B2(new_n565), .ZN(new_n933));
  NOR2_X1   g508(.A1(G171), .A2(G168), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n850), .B(new_n852), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(G168), .B1(new_n566), .B2(new_n567), .ZN(new_n936));
  INV_X1    g511(.A(new_n934), .ZN(new_n937));
  OR3_X1    g512(.A1(new_n834), .A2(KEYINPUT102), .A3(new_n837), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n550), .B1(new_n938), .B2(new_n838), .ZN(new_n939));
  INV_X1    g514(.A(new_n852), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n936), .B(new_n937), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n935), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n916), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n935), .A2(new_n941), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n920), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n922), .A2(KEYINPUT110), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n914), .A2(new_n949), .A3(new_n921), .A4(new_n915), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n916), .A2(KEYINPUT111), .A3(KEYINPUT41), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n947), .A2(new_n948), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n944), .A2(KEYINPUT112), .B1(new_n945), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n916), .B1(new_n935), .B2(new_n941), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n911), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n935), .A2(new_n923), .A3(new_n941), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n944), .A2(new_n911), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n893), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n930), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n911), .ZN(new_n962));
  INV_X1    g537(.A(new_n952), .ZN(new_n963));
  OAI22_X1  g538(.A1(new_n963), .A2(new_n942), .B1(new_n955), .B2(new_n954), .ZN(new_n964));
  INV_X1    g539(.A(new_n956), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n960), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(new_n967), .A3(KEYINPUT113), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n929), .B1(new_n961), .B2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n958), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n962), .B1(new_n970), .B2(new_n954), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT43), .B1(new_n967), .B2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT44), .B1(new_n969), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n971), .A2(new_n893), .A3(new_n959), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(KEYINPUT43), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT109), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n974), .A2(new_n977), .A3(KEYINPUT43), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n966), .A2(new_n967), .A3(new_n929), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n976), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n973), .A2(new_n982), .ZN(G397));
  XNOR2_X1  g558(.A(KEYINPUT114), .B(G1384), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n497), .B1(new_n493), .B2(new_n495), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n984), .B1(new_n985), .B2(new_n874), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n476), .A2(G40), .A3(new_n479), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n986), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1996), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(new_n991), .A3(new_n758), .ZN(new_n992));
  XOR2_X1   g567(.A(new_n992), .B(KEYINPUT115), .Z(new_n993));
  INV_X1    g568(.A(G2067), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n731), .B(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n991), .B2(new_n758), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n993), .B1(new_n990), .B2(new_n996), .ZN(new_n997));
  XOR2_X1   g572(.A(new_n822), .B(new_n824), .Z(new_n998));
  OAI21_X1  g573(.A(new_n997), .B1(new_n989), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n812), .A2(new_n814), .ZN(new_n1000));
  NAND2_X1  g575(.A1(G290), .A2(G1986), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n989), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT118), .ZN(new_n1004));
  NAND2_X1  g579(.A1(G303), .A2(G8), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT55), .ZN(new_n1006));
  OAI211_X1 g581(.A(KEYINPUT45), .B(new_n984), .C1(new_n985), .C2(new_n874), .ZN(new_n1007));
  AND2_X1   g582(.A1(new_n1007), .A2(new_n987), .ZN(new_n1008));
  INV_X1    g583(.A(G1384), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(new_n985), .B2(new_n505), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(new_n988), .ZN(new_n1011));
  AOI21_X1  g586(.A(G1971), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1009), .B1(new_n985), .B2(new_n874), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT50), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT117), .B1(new_n1014), .B2(new_n987), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT117), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n476), .A2(G40), .A3(new_n479), .ZN(new_n1017));
  AOI211_X1 g592(.A(new_n1016), .B(new_n1017), .C1(new_n1013), .C2(KEYINPUT50), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n1019));
  OAI211_X1 g594(.A(new_n1019), .B(new_n1009), .C1(new_n985), .C2(new_n505), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n1015), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1012), .B1(new_n1022), .B2(new_n698), .ZN(new_n1023));
  INV_X1    g598(.A(G8), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1004), .B(new_n1006), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1014), .A2(new_n987), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n1016), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1017), .B1(new_n1013), .B2(KEYINPUT50), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1021), .B1(new_n1028), .B2(KEYINPUT117), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n1029), .A3(new_n698), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1012), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1024), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1006), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT118), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1035));
  INV_X1    g610(.A(G48), .ZN(new_n1036));
  OAI22_X1  g611(.A1(new_n511), .A2(new_n1035), .B1(new_n543), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n533), .A2(new_n581), .ZN(new_n1038));
  OAI21_X1  g613(.A(G1981), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1039), .B1(G305), .B2(G1981), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT49), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n879), .A2(new_n987), .A3(new_n1009), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1039), .B(KEYINPUT49), .C1(G305), .C2(G1981), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1042), .A2(G8), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1046), .B(new_n1047), .C1(new_n799), .C2(G1976), .ZN(new_n1048));
  AOI21_X1  g623(.A(G1976), .B1(new_n572), .B2(new_n579), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT116), .B1(new_n1049), .B2(KEYINPUT52), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G1976), .ZN(new_n1052));
  OAI221_X1 g627(.A(G8), .B1(G288), .B2(new_n1052), .C1(new_n1017), .C2(new_n1013), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1045), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  AND2_X1   g629(.A1(new_n1053), .A2(KEYINPUT52), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n879), .A2(new_n1019), .A3(new_n1009), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1010), .A2(KEYINPUT50), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n987), .A3(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1059), .A2(G2090), .ZN(new_n1060));
  OAI211_X1 g635(.A(G8), .B(new_n1033), .C1(new_n1060), .C2(new_n1012), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1056), .A2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n987), .B1(new_n1013), .B2(KEYINPUT50), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1019), .B1(new_n507), .B2(new_n1009), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G2084), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1017), .B1(new_n1013), .B2(new_n988), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n1009), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1065), .A2(new_n1066), .B1(new_n1069), .B2(new_n720), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1070), .A2(new_n1024), .A3(G286), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1025), .A2(new_n1034), .A3(new_n1062), .A4(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(KEYINPUT119), .B(KEYINPUT63), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1071), .A2(KEYINPUT63), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1060), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1024), .B1(new_n1076), .B2(new_n1031), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n1078));
  AND2_X1   g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1006), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1075), .B(new_n1062), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1074), .A2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1011), .A2(new_n765), .A3(new_n987), .A4(new_n1007), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G1961), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1086), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1067), .A2(new_n1068), .A3(KEYINPUT53), .A4(new_n765), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n606), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1069), .A2(new_n720), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1057), .A2(new_n1058), .A3(new_n1066), .A4(new_n987), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(G168), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT51), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1094), .A2(KEYINPUT125), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(KEYINPUT125), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1093), .A2(G8), .A3(new_n1096), .A4(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(G8), .A3(G286), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1024), .B1(new_n1070), .B2(G168), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1098), .B(new_n1100), .C1(new_n1101), .C2(new_n1096), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1090), .B1(new_n1102), .B2(KEYINPUT62), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1056), .A2(new_n1061), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1006), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1104), .B1(new_n1105), .B2(KEYINPUT118), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1093), .A2(G8), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n1095), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1108), .A2(new_n1109), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1103), .A2(new_n1025), .A3(new_n1106), .A4(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1043), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1045), .A2(new_n1052), .A3(new_n799), .ZN(new_n1113));
  OR2_X1    g688(.A1(G305), .A2(G1981), .ZN(new_n1114));
  AOI211_X1 g689(.A(new_n1024), .B(new_n1112), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1061), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1115), .B1(new_n1116), .B2(new_n1056), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1082), .A2(new_n1111), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n986), .A2(new_n988), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1008), .A2(KEYINPUT53), .A3(new_n765), .A4(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1085), .A2(new_n1120), .A3(new_n1087), .A4(G301), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1090), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1085), .A2(new_n1120), .A3(new_n1087), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1123), .B1(new_n1124), .B2(G171), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .A4(G301), .ZN(new_n1126));
  AOI22_X1  g701(.A1(new_n1122), .A2(new_n1123), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1106), .A2(new_n1025), .A3(new_n1102), .A4(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(G1956), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1014), .A2(KEYINPUT117), .A3(new_n987), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n1020), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1129), .B1(new_n1131), .B2(new_n1015), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT57), .B1(new_n563), .B2(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g709(.A(G299), .B(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT56), .B(G2072), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1008), .A2(new_n1011), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1132), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1132), .A2(new_n1137), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1135), .B1(new_n1139), .B2(KEYINPUT122), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1132), .A2(new_n1141), .A3(new_n1137), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT123), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(G1956), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1137), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT122), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1135), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1146), .A2(new_n1142), .A3(KEYINPUT123), .A4(new_n1147), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1059), .A2(new_n742), .B1(new_n1112), .B2(new_n994), .ZN(new_n1149));
  INV_X1    g724(.A(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n611), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1148), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1138), .B1(new_n1143), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1154), .B1(new_n1149), .B2(KEYINPUT60), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1149), .A2(new_n1154), .A3(KEYINPUT60), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(new_n611), .A3(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1149), .A2(KEYINPUT60), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1159), .B1(new_n1155), .B2(new_n604), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1135), .B1(new_n1132), .B2(new_n1137), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1163));
  XNOR2_X1  g738(.A(KEYINPUT58), .B(G1341), .ZN(new_n1164));
  OAI22_X1  g739(.A1(new_n1163), .A2(G1996), .B1(new_n1112), .B2(new_n1164), .ZN(new_n1165));
  AND3_X1   g740(.A1(new_n1165), .A2(KEYINPUT59), .A3(new_n550), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT59), .B1(new_n1165), .B2(new_n550), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1162), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n1138), .A2(KEYINPUT61), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1138), .A2(KEYINPUT61), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1161), .A2(new_n1168), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1128), .B1(new_n1153), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1003), .B1(new_n1118), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n989), .B1(new_n995), .B2(new_n758), .ZN(new_n1174));
  XOR2_X1   g749(.A(new_n1174), .B(KEYINPUT126), .Z(new_n1175));
  NAND2_X1  g750(.A1(new_n990), .A2(new_n991), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1176), .B(KEYINPUT46), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  XOR2_X1   g753(.A(new_n1178), .B(KEYINPUT47), .Z(new_n1179));
  NOR2_X1   g754(.A1(new_n1000), .A2(new_n989), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1180), .B(KEYINPUT127), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(KEYINPUT48), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n999), .A2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n822), .A2(new_n824), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n997), .A2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n726), .A2(new_n994), .A3(new_n730), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n989), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1179), .A2(new_n1183), .A3(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1173), .A2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g764(.A1(G227), .A2(new_n459), .A3(new_n461), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n691), .A2(new_n1191), .ZN(new_n1192));
  AOI21_X1  g766(.A(new_n1192), .B1(new_n651), .B2(new_n652), .ZN(new_n1193));
  NAND2_X1  g767(.A1(new_n895), .A2(new_n897), .ZN(new_n1194));
  AND3_X1   g768(.A1(new_n1193), .A2(new_n980), .A3(new_n1194), .ZN(G308));
  NAND3_X1  g769(.A1(new_n1193), .A2(new_n980), .A3(new_n1194), .ZN(G225));
endmodule


