//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 1 0 0 1 0 0 0 0 0 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n805, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(G190gat), .ZN(new_n203));
  NAND3_X1  g002(.A1(new_n202), .A2(KEYINPUT28), .A3(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G183gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT27), .B1(new_n205), .B2(KEYINPUT66), .ZN(new_n206));
  OR3_X1    g005(.A1(new_n205), .A2(KEYINPUT66), .A3(KEYINPUT27), .ZN(new_n207));
  AND3_X1   g006(.A1(new_n206), .A2(new_n207), .A3(new_n203), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n204), .B1(new_n208), .B2(KEYINPUT28), .ZN(new_n209));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210));
  INV_X1    g009(.A(G169gat), .ZN(new_n211));
  INV_X1    g010(.A(G176gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT26), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n210), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT26), .B1(new_n211), .B2(new_n212), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n209), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n210), .A2(KEYINPUT24), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n205), .A2(G190gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n203), .A2(G183gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n220), .B1(new_n223), .B2(KEYINPUT24), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n211), .A2(new_n212), .A3(KEYINPUT23), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(new_n216), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(KEYINPUT65), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(G169gat), .B2(G176gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(KEYINPUT25), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n225), .A2(new_n232), .A3(new_n216), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n224), .A2(new_n227), .A3(new_n231), .A4(new_n233), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n225), .A2(new_n229), .A3(new_n216), .ZN(new_n235));
  AOI21_X1  g034(.A(KEYINPUT25), .B1(new_n224), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT64), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n234), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT25), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT24), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(G183gat), .A3(G190gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(G183gat), .B(G190gat), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n241), .B1(new_n242), .B2(new_n240), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n225), .A2(new_n229), .A3(new_n216), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n239), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(KEYINPUT64), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n219), .B1(new_n238), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G226gat), .ZN(new_n248));
  INV_X1    g047(.A(G233gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G197gat), .B(G204gat), .ZN(new_n252));
  INV_X1    g051(.A(G211gat), .ZN(new_n253));
  INV_X1    g052(.A(G218gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n252), .B1(KEYINPUT22), .B2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G211gat), .B(G218gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n236), .A2(new_n237), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT64), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(new_n261), .A3(new_n234), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT29), .B1(new_n262), .B2(new_n219), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n251), .B(new_n259), .C1(new_n263), .C2(new_n250), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT75), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT74), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT29), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n250), .B1(new_n247), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n250), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n269), .B1(new_n262), .B2(new_n219), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n266), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(KEYINPUT74), .B1(new_n263), .B2(new_n250), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n265), .B1(new_n273), .B2(new_n258), .ZN(new_n274));
  AOI211_X1 g073(.A(KEYINPUT75), .B(new_n259), .C1(new_n271), .C2(new_n272), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT76), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G8gat), .B(G36gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(G64gat), .B(G92gat), .ZN(new_n278));
  XOR2_X1   g077(.A(new_n277), .B(new_n278), .Z(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT75), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n243), .A2(new_n230), .ZN(new_n282));
  INV_X1    g081(.A(new_n233), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n232), .B1(new_n225), .B2(new_n216), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n245), .A2(KEYINPUT64), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  AOI22_X1  g085(.A1(new_n286), .A2(new_n260), .B1(new_n209), .B2(new_n218), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n269), .B1(new_n287), .B2(KEYINPUT29), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT74), .B1(new_n288), .B2(new_n251), .ZN(new_n289));
  INV_X1    g088(.A(new_n272), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n281), .B(new_n258), .C1(new_n289), .C2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT76), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n259), .B1(new_n271), .B2(new_n272), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n291), .B(new_n292), .C1(new_n293), .C2(new_n265), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n276), .A2(new_n280), .A3(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n291), .B1(new_n293), .B2(new_n265), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n296), .A2(KEYINPUT30), .A3(new_n279), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n279), .B1(new_n274), .B2(new_n275), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT30), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n295), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G225gat), .A2(G233gat), .ZN(new_n302));
  XOR2_X1   g101(.A(G141gat), .B(G148gat), .Z(new_n303));
  INV_X1    g102(.A(KEYINPUT2), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G155gat), .B(G162gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT77), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT77), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(G155gat), .B2(G162gat), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n305), .A2(new_n307), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT78), .B(G162gat), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n304), .B1(new_n311), .B2(G155gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n303), .A2(new_n306), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n310), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(G134gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G127gat), .ZN(new_n316));
  INV_X1    g115(.A(G127gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G134gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n316), .A2(new_n318), .A3(KEYINPUT67), .ZN(new_n319));
  XNOR2_X1  g118(.A(G113gat), .B(G120gat), .ZN(new_n320));
  OAI221_X1 g119(.A(new_n319), .B1(KEYINPUT67), .B2(new_n316), .C1(KEYINPUT1), .C2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT69), .ZN(new_n322));
  INV_X1    g121(.A(G120gat), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n322), .B1(new_n323), .B2(G113gat), .ZN(new_n324));
  OR2_X1    g123(.A1(KEYINPUT68), .A2(G120gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(KEYINPUT68), .A2(G120gat), .ZN(new_n326));
  AND2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n324), .B1(new_n327), .B2(G113gat), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n325), .A2(KEYINPUT69), .A3(G113gat), .A4(new_n326), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT1), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n329), .A2(new_n330), .A3(new_n316), .A4(new_n318), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n321), .B1(new_n328), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT4), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n314), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT70), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n314), .ZN(new_n337));
  OAI211_X1 g136(.A(new_n321), .B(KEYINPUT70), .C1(new_n328), .C2(new_n331), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n334), .B1(new_n339), .B2(new_n333), .ZN(new_n340));
  OR2_X1    g139(.A1(new_n313), .A2(new_n312), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n341), .A2(new_n342), .A3(new_n310), .ZN(new_n343));
  AOI211_X1 g142(.A(KEYINPUT79), .B(new_n342), .C1(new_n341), .C2(new_n310), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT79), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n345), .B1(new_n314), .B2(KEYINPUT3), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n332), .B(new_n343), .C1(new_n344), .C2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n302), .B1(new_n340), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n314), .B(new_n332), .ZN(new_n349));
  INV_X1    g148(.A(new_n302), .ZN(new_n350));
  OAI21_X1  g149(.A(KEYINPUT39), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OR2_X1    g150(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  XOR2_X1   g151(.A(G1gat), .B(G29gat), .Z(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT81), .ZN(new_n354));
  XOR2_X1   g153(.A(G57gat), .B(G85gat), .Z(new_n355));
  XNOR2_X1  g154(.A(new_n354), .B(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT39), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(new_n348), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT86), .B1(new_n352), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT40), .ZN(new_n362));
  AND2_X1   g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n358), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n333), .B1(new_n314), .B2(new_n332), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT4), .A4(new_n338), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n347), .A2(new_n302), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT5), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n368), .B1(new_n349), .B2(new_n350), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n340), .A2(new_n347), .A3(new_n368), .A4(new_n302), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n364), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n373), .B1(new_n361), .B2(new_n362), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n363), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n301), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n343), .A2(new_n267), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n258), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n342), .B1(new_n258), .B2(KEYINPUT29), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n314), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n378), .A2(KEYINPUT84), .ZN(new_n382));
  INV_X1    g181(.A(G228gat), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n382), .B1(new_n383), .B2(new_n249), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(G22gat), .ZN(new_n385));
  INV_X1    g184(.A(G22gat), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n382), .B(new_n386), .C1(new_n383), .C2(new_n249), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n381), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT85), .ZN(new_n390));
  XNOR2_X1  g189(.A(G78gat), .B(G106gat), .ZN(new_n391));
  INV_X1    g190(.A(G50gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  XOR2_X1   g192(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n394));
  XNOR2_X1  g193(.A(new_n393), .B(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n385), .A2(new_n381), .A3(new_n387), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n389), .A2(new_n390), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n395), .B(KEYINPUT85), .ZN(new_n398));
  INV_X1    g197(.A(new_n396), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n398), .B1(new_n399), .B2(new_n388), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT38), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n276), .A2(KEYINPUT37), .A3(new_n294), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT37), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n279), .B1(new_n296), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n402), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n370), .A2(new_n371), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(KEYINPUT6), .A3(new_n358), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT82), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT82), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n372), .A2(new_n410), .A3(KEYINPUT6), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n372), .A2(KEYINPUT6), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n370), .A2(new_n364), .A3(new_n371), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n409), .A2(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n296), .A2(new_n404), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n273), .A2(new_n259), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n268), .A2(new_n270), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n404), .B1(new_n417), .B2(new_n258), .ZN(new_n418));
  AOI21_X1  g217(.A(KEYINPUT38), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n415), .A2(new_n280), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n414), .A2(new_n420), .A3(new_n298), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n376), .B(new_n401), .C1(new_n406), .C2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT36), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n336), .A2(new_n338), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n247), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(G227gat), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n426), .A2(new_n249), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n262), .A2(new_n336), .A3(new_n338), .A4(new_n219), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n425), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n430), .A2(KEYINPUT73), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT72), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT32), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n425), .A2(new_n429), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n433), .B1(new_n434), .B2(new_n427), .ZN(new_n435));
  XNOR2_X1  g234(.A(G15gat), .B(G43gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(G71gat), .B(G99gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n436), .B(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT33), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n432), .B1(new_n435), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n428), .B1(new_n425), .B2(new_n429), .ZN(new_n443));
  NOR4_X1   g242(.A1(new_n443), .A2(KEYINPUT72), .A3(new_n433), .A4(new_n440), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n442), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n438), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n443), .B2(new_n433), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT71), .B1(new_n443), .B2(KEYINPUT33), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n247), .A2(new_n424), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n262), .A2(new_n219), .B1(new_n336), .B2(new_n338), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n427), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT71), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n452), .A3(new_n439), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n447), .B1(new_n448), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n431), .B1(new_n445), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n453), .A2(new_n448), .ZN(new_n456));
  INV_X1    g255(.A(new_n447), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n451), .A2(KEYINPUT32), .A3(new_n441), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT72), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n435), .A2(new_n432), .A3(new_n441), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n431), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n458), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n430), .A2(KEYINPUT73), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n465), .A2(KEYINPUT34), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n455), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n467), .B1(new_n455), .B2(new_n464), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n423), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n445), .A2(new_n454), .A3(new_n431), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n463), .B1(new_n458), .B2(new_n462), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n466), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n464), .A3(new_n467), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n473), .A2(KEYINPUT36), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT6), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n373), .A2(new_n476), .A3(new_n413), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n408), .A2(KEYINPUT82), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n410), .B1(new_n372), .B2(KEYINPUT6), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n480), .A2(new_n295), .A3(new_n297), .A4(new_n300), .ZN(new_n481));
  INV_X1    g280(.A(new_n401), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n470), .A2(new_n475), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n301), .A2(new_n414), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT35), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .A4(new_n401), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n473), .A2(new_n401), .A3(new_n474), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT35), .B1(new_n488), .B2(new_n481), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n422), .A2(new_n483), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G43gat), .B(G50gat), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT87), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT15), .ZN(new_n495));
  INV_X1    g294(.A(G43gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n496), .A2(KEYINPUT87), .A3(G50gat), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(G29gat), .A2(G36gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT14), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n492), .A2(KEYINPUT15), .ZN(new_n502));
  NAND2_X1  g301(.A1(G29gat), .A2(G36gat), .ZN(new_n503));
  XOR2_X1   g302(.A(new_n503), .B(KEYINPUT88), .Z(new_n504));
  NAND4_X1  g303(.A1(new_n498), .A2(new_n501), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n501), .A2(new_n503), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n505), .B1(new_n506), .B2(new_n502), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(KEYINPUT17), .ZN(new_n508));
  NAND2_X1  g307(.A1(G85gat), .A2(G92gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n510));
  XOR2_X1   g309(.A(new_n509), .B(new_n510), .Z(new_n511));
  NAND2_X1  g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512));
  INV_X1    g311(.A(G85gat), .ZN(new_n513));
  INV_X1    g312(.A(G92gat), .ZN(new_n514));
  AOI22_X1  g313(.A1(KEYINPUT8), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G99gat), .B(G106gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n508), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT95), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n508), .A2(KEYINPUT95), .A3(new_n519), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(G232gat), .A2(G233gat), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n518), .A2(new_n507), .B1(KEYINPUT41), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G190gat), .B(G218gat), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n529), .B(KEYINPUT96), .Z(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n526), .A2(KEYINPUT41), .ZN(new_n532));
  XNOR2_X1  g331(.A(G134gat), .B(G162gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(KEYINPUT97), .ZN(new_n535));
  INV_X1    g334(.A(new_n530), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n524), .A2(new_n536), .A3(new_n527), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n531), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n534), .B(KEYINPUT97), .Z(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n541), .B1(new_n531), .B2(new_n537), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G15gat), .B(G22gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT16), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n545), .B1(new_n546), .B2(G1gat), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(G1gat), .B2(new_n545), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(G8gat), .ZN(new_n549));
  XOR2_X1   g348(.A(G57gat), .B(G64gat), .Z(new_n550));
  NAND2_X1  g349(.A1(G71gat), .A2(G78gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT9), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n550), .B1(KEYINPUT90), .B2(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n553), .A2(KEYINPUT90), .ZN(new_n555));
  INV_X1    g354(.A(new_n551), .ZN(new_n556));
  OAI22_X1  g355(.A1(new_n554), .A2(new_n555), .B1(KEYINPUT89), .B2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(G71gat), .B(G78gat), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n557), .B(new_n558), .Z(new_n559));
  AOI21_X1  g358(.A(new_n549), .B1(new_n559), .B2(KEYINPUT21), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT93), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n559), .A2(KEYINPUT21), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n561), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G127gat), .B(G155gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT92), .ZN(new_n567));
  NAND2_X1  g366(.A1(G231gat), .A2(G233gat), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n568), .B(KEYINPUT91), .Z(new_n569));
  XNOR2_X1  g368(.A(new_n567), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G183gat), .B(G211gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n570), .B(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n565), .B(new_n572), .Z(new_n573));
  INV_X1    g372(.A(KEYINPUT98), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n518), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT10), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n557), .B(new_n558), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(new_n519), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n559), .A2(KEYINPUT10), .A3(new_n518), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G230gat), .A2(G233gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n575), .A2(new_n578), .ZN(new_n584));
  INV_X1    g383(.A(new_n582), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G120gat), .B(G148gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(G176gat), .B(G204gat), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n588), .B(new_n589), .Z(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n574), .B1(new_n587), .B2(new_n591), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n583), .A2(KEYINPUT98), .A3(new_n586), .A4(new_n590), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n587), .A2(new_n591), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n544), .A2(new_n573), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n549), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n508), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n549), .A2(new_n507), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G229gat), .A2(G233gat), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(KEYINPUT18), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n549), .B(new_n507), .ZN(new_n605));
  XOR2_X1   g404(.A(new_n603), .B(KEYINPUT13), .Z(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n600), .A2(new_n603), .A3(new_n601), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT18), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n604), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G113gat), .B(G141gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(G197gat), .ZN(new_n613));
  XOR2_X1   g412(.A(KEYINPUT11), .B(G169gat), .Z(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n615), .B(KEYINPUT12), .Z(new_n616));
  NAND2_X1  g415(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n616), .ZN(new_n618));
  NAND4_X1  g417(.A1(new_n604), .A2(new_n618), .A3(new_n607), .A4(new_n610), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n598), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n491), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(new_n414), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g425(.A(KEYINPUT16), .B(G8gat), .Z(new_n627));
  INV_X1    g426(.A(KEYINPUT42), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT100), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n627), .B(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n301), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n623), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n630), .B1(new_n632), .B2(new_n628), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT99), .ZN(new_n634));
  OAI22_X1  g433(.A1(new_n632), .A2(new_n634), .B1(new_n628), .B2(G8gat), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n623), .A2(KEYINPUT99), .A3(new_n631), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n637), .B(KEYINPUT101), .Z(G1325gat));
  AOI21_X1  g437(.A(G15gat), .B1(new_n624), .B2(new_n485), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(KEYINPUT102), .Z(new_n640));
  NAND2_X1  g439(.A1(new_n470), .A2(new_n475), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n642), .A2(G15gat), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n640), .B1(new_n624), .B2(new_n643), .ZN(G1326gat));
  NOR2_X1   g443(.A1(new_n623), .A2(new_n401), .ZN(new_n645));
  XOR2_X1   g444(.A(KEYINPUT43), .B(G22gat), .Z(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(G1327gat));
  INV_X1    g446(.A(KEYINPUT106), .ZN(new_n648));
  INV_X1    g447(.A(G29gat), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n544), .A2(KEYINPUT44), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT104), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n481), .A2(new_n482), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n422), .A2(new_n641), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n487), .A2(new_n489), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n651), .B1(new_n483), .B2(new_n422), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n650), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT44), .B1(new_n490), .B2(new_n544), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n573), .A2(new_n621), .A3(new_n596), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT105), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT105), .ZN(new_n662));
  INV_X1    g461(.A(new_n660), .ZN(new_n663));
  AOI211_X1 g462(.A(new_n662), .B(new_n663), .C1(new_n657), .C2(new_n658), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n649), .B1(new_n665), .B2(new_n414), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n490), .A2(new_n544), .A3(new_n663), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n667), .A2(new_n649), .A3(new_n414), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n648), .B1(new_n666), .B2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n670), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n661), .A2(new_n664), .A3(new_n480), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n672), .B(KEYINPUT106), .C1(new_n673), .C2(new_n649), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n671), .A2(new_n674), .ZN(G1328gat));
  INV_X1    g474(.A(G36gat), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n667), .A2(new_n676), .A3(new_n301), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT107), .B(KEYINPUT46), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n661), .A2(new_n664), .A3(new_n631), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n679), .B1(new_n680), .B2(new_n676), .ZN(G1329gat));
  NAND2_X1  g480(.A1(new_n659), .A2(new_n660), .ZN(new_n682));
  OAI21_X1  g481(.A(G43gat), .B1(new_n682), .B2(new_n641), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n667), .A2(new_n496), .A3(new_n485), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(KEYINPUT47), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n684), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n665), .A2(new_n642), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n686), .B1(new_n687), .B2(G43gat), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n685), .B1(new_n688), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g488(.A(G50gat), .B1(new_n682), .B2(new_n401), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n667), .A2(new_n392), .A3(new_n482), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n690), .A2(KEYINPUT48), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n691), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n665), .A2(new_n482), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n693), .B1(new_n694), .B2(G50gat), .ZN(new_n695));
  XOR2_X1   g494(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n696));
  OAI21_X1  g495(.A(new_n692), .B1(new_n695), .B2(new_n696), .ZN(G1331gat));
  OR2_X1    g496(.A1(new_n655), .A2(new_n656), .ZN(new_n698));
  INV_X1    g497(.A(new_n573), .ZN(new_n699));
  NOR4_X1   g498(.A1(new_n597), .A2(new_n699), .A3(new_n543), .A4(new_n620), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n414), .B(KEYINPUT109), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g503(.A(new_n301), .B(KEYINPUT110), .Z(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n701), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n707), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n708));
  XOR2_X1   g507(.A(KEYINPUT49), .B(G64gat), .Z(new_n709));
  OAI21_X1  g508(.A(new_n708), .B1(new_n707), .B2(new_n709), .ZN(G1333gat));
  NAND4_X1  g509(.A1(new_n698), .A2(G71gat), .A3(new_n642), .A4(new_n700), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT111), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n701), .A2(new_n485), .ZN(new_n713));
  INV_X1    g512(.A(G71gat), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT50), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT50), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n712), .A2(new_n718), .A3(new_n715), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n717), .A2(new_n719), .ZN(G1334gat));
  NAND2_X1  g519(.A1(new_n701), .A2(new_n482), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g521(.A1(new_n544), .A2(new_n573), .A3(new_n620), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n698), .A2(KEYINPUT51), .A3(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT51), .B1(new_n698), .B2(new_n723), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n596), .A2(new_n513), .A3(new_n414), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT112), .ZN(new_n729));
  INV_X1    g528(.A(new_n659), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n699), .A2(new_n621), .A3(new_n596), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n730), .A2(new_n480), .A3(new_n731), .ZN(new_n732));
  OAI22_X1  g531(.A1(new_n727), .A2(new_n729), .B1(new_n732), .B2(new_n513), .ZN(G1336gat));
  INV_X1    g532(.A(KEYINPUT52), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n730), .A2(new_n705), .A3(new_n731), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n705), .A2(G92gat), .A3(new_n597), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  OAI221_X1 g536(.A(new_n734), .B1(new_n735), .B2(new_n514), .C1(new_n727), .C2(new_n737), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n736), .B(KEYINPUT113), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n727), .A2(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n730), .A2(new_n731), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n514), .B1(new_n741), .B2(new_n301), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT52), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n738), .A2(new_n743), .ZN(G1337gat));
  NOR2_X1   g543(.A1(new_n727), .A2(new_n597), .ZN(new_n745));
  XOR2_X1   g544(.A(KEYINPUT114), .B(G99gat), .Z(new_n746));
  NAND3_X1  g545(.A1(new_n745), .A2(new_n485), .A3(new_n746), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n730), .A2(new_n641), .A3(new_n731), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(new_n746), .ZN(G1338gat));
  NOR3_X1   g548(.A1(new_n730), .A2(new_n401), .A3(new_n731), .ZN(new_n750));
  INV_X1    g549(.A(G106gat), .ZN(new_n751));
  OR2_X1    g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n401), .A2(G106gat), .ZN(new_n754));
  OAI211_X1 g553(.A(new_n596), .B(new_n754), .C1(new_n725), .C2(new_n726), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n752), .A2(KEYINPUT115), .A3(new_n753), .A4(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(KEYINPUT115), .B1(new_n750), .B2(new_n751), .ZN(new_n757));
  INV_X1    g556(.A(new_n755), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT53), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n756), .A2(new_n759), .ZN(G1339gat));
  INV_X1    g559(.A(new_n542), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n602), .A2(new_n603), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n605), .A2(new_n606), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n615), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n619), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n761), .A2(new_n766), .A3(new_n538), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n585), .B1(new_n579), .B2(new_n580), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT54), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n590), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n583), .A2(KEYINPUT54), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n581), .A2(new_n582), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT55), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  OAI211_X1 g574(.A(KEYINPUT55), .B(new_n770), .C1(new_n771), .C2(new_n772), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n775), .A2(new_n594), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(KEYINPUT116), .B1(new_n767), .B2(new_n777), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n539), .A2(new_n542), .A3(new_n765), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n775), .A2(new_n594), .A3(new_n776), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n778), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n596), .A2(new_n766), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n620), .A2(new_n594), .A3(new_n775), .A4(new_n776), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n543), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n699), .B1(new_n783), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n598), .A2(new_n620), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n790), .A2(new_n482), .ZN(new_n791));
  INV_X1    g590(.A(new_n485), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n706), .A2(new_n480), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(G113gat), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n794), .A2(new_n795), .A3(new_n621), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n787), .A2(new_n789), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n797), .A2(new_n401), .A3(new_n485), .A4(new_n702), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n798), .A2(new_n706), .ZN(new_n799));
  AOI21_X1  g598(.A(G113gat), .B1(new_n799), .B2(new_n620), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n796), .A2(new_n800), .ZN(G1340gat));
  OAI21_X1  g600(.A(G120gat), .B1(new_n794), .B2(new_n597), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n799), .A2(new_n327), .A3(new_n596), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(G1341gat));
  OAI21_X1  g603(.A(G127gat), .B1(new_n794), .B2(new_n699), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n799), .A2(new_n317), .A3(new_n573), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(G1342gat));
  OAI21_X1  g606(.A(G134gat), .B1(new_n794), .B2(new_n544), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT56), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n631), .A2(new_n543), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n798), .A2(G134gat), .A3(new_n810), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n811), .A2(KEYINPUT117), .A3(new_n809), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT117), .B1(new_n811), .B2(new_n809), .ZN(new_n813));
  OAI221_X1 g612(.A(new_n808), .B1(new_n809), .B2(new_n811), .C1(new_n812), .C2(new_n813), .ZN(G1343gat));
  INV_X1    g613(.A(KEYINPUT58), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n797), .A2(KEYINPUT121), .A3(new_n702), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n641), .A2(new_n482), .ZN(new_n817));
  INV_X1    g616(.A(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT121), .ZN(new_n820));
  INV_X1    g619(.A(new_n702), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n820), .B1(new_n790), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n621), .A2(G141gat), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n819), .A2(new_n705), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n815), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(G141gat), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n706), .A2(new_n480), .A3(new_n642), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n482), .A2(KEYINPUT57), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n777), .A2(KEYINPUT118), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n775), .A2(new_n594), .A3(new_n832), .A4(new_n776), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n831), .A2(new_n620), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n543), .B1(new_n834), .B2(new_n784), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n699), .B1(new_n835), .B2(new_n783), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n830), .B1(new_n836), .B2(new_n789), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(KEYINPUT119), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n797), .A2(new_n482), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841));
  AOI22_X1  g640(.A1(new_n837), .A2(KEYINPUT119), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n829), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n827), .B1(new_n843), .B2(new_n620), .ZN(new_n844));
  INV_X1    g643(.A(new_n824), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n826), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n837), .A2(KEYINPUT119), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n840), .A2(new_n841), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n828), .B1(new_n849), .B2(new_n838), .ZN(new_n850));
  OAI21_X1  g649(.A(G141gat), .B1(new_n850), .B2(new_n621), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n822), .A2(new_n705), .A3(new_n818), .A4(new_n816), .ZN(new_n852));
  INV_X1    g651(.A(new_n823), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n825), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT58), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n851), .A2(new_n855), .A3(new_n824), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n846), .A2(new_n856), .ZN(G1344gat));
  INV_X1    g656(.A(G148gat), .ZN(new_n858));
  AOI211_X1 g657(.A(KEYINPUT59), .B(new_n858), .C1(new_n843), .C2(new_n596), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860));
  INV_X1    g659(.A(new_n835), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n779), .A2(new_n780), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n573), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n841), .B(new_n482), .C1(new_n863), .C2(new_n788), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n840), .A2(KEYINPUT57), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n596), .A3(new_n828), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n860), .B1(new_n867), .B2(G148gat), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n596), .A2(new_n858), .ZN(new_n869));
  OAI22_X1  g668(.A1(new_n859), .A2(new_n868), .B1(new_n852), .B2(new_n869), .ZN(G1345gat));
  INV_X1    g669(.A(G155gat), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n871), .B1(new_n852), .B2(new_n699), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n573), .A2(G155gat), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT122), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n872), .B1(new_n850), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n872), .B(KEYINPUT123), .C1(new_n850), .C2(new_n874), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(G1346gat));
  OAI21_X1  g678(.A(new_n311), .B1(new_n850), .B2(new_n544), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n810), .A2(new_n311), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n819), .A2(new_n822), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(G1347gat));
  NOR4_X1   g682(.A1(new_n790), .A2(new_n414), .A3(new_n488), .A4(new_n705), .ZN(new_n884));
  AOI21_X1  g683(.A(G169gat), .B1(new_n884), .B2(new_n620), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n821), .A2(new_n301), .ZN(new_n886));
  NOR4_X1   g685(.A1(new_n790), .A2(new_n482), .A3(new_n792), .A4(new_n886), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n621), .A2(new_n211), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n885), .B1(new_n887), .B2(new_n888), .ZN(G1348gat));
  NAND3_X1  g688(.A1(new_n884), .A2(new_n212), .A3(new_n596), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n887), .A2(new_n596), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n890), .B1(new_n891), .B2(new_n212), .ZN(G1349gat));
  NAND3_X1  g691(.A1(new_n884), .A2(new_n202), .A3(new_n573), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n887), .A2(new_n573), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n894), .B2(new_n205), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g695(.A1(new_n884), .A2(new_n203), .A3(new_n543), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n887), .A2(new_n543), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(G190gat), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n899), .A2(KEYINPUT61), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(KEYINPUT61), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n897), .B1(new_n900), .B2(new_n901), .ZN(G1351gat));
  XNOR2_X1  g701(.A(KEYINPUT124), .B(G197gat), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n886), .A2(new_n642), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n866), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n903), .B1(new_n905), .B2(new_n621), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n797), .A2(new_n480), .A3(new_n706), .A4(new_n818), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n621), .A2(new_n903), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n906), .B1(new_n907), .B2(new_n908), .ZN(G1352gat));
  OAI21_X1  g708(.A(G204gat), .B1(new_n905), .B2(new_n597), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n907), .A2(G204gat), .A3(new_n597), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n912));
  OR2_X1    g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n912), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n910), .A2(new_n913), .A3(new_n914), .ZN(G1353gat));
  NAND3_X1  g714(.A1(new_n866), .A2(new_n573), .A3(new_n904), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n916), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT63), .B1(new_n916), .B2(G211gat), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n573), .A2(new_n253), .ZN(new_n919));
  OAI22_X1  g718(.A1(new_n917), .A2(new_n918), .B1(new_n907), .B2(new_n919), .ZN(G1354gat));
  AND2_X1   g719(.A1(new_n866), .A2(new_n904), .ZN(new_n921));
  OR2_X1    g720(.A1(new_n921), .A2(KEYINPUT126), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n543), .A2(G218gat), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n923), .B1(new_n921), .B2(KEYINPUT126), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n254), .B1(new_n907), .B2(new_n544), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT125), .ZN(new_n926));
  OR2_X1    g725(.A1(new_n925), .A2(KEYINPUT125), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n922), .A2(new_n924), .B1(new_n926), .B2(new_n927), .ZN(G1355gat));
endmodule


