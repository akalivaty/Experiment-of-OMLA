//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1 0 1 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n446, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n553, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n605, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT64), .B(G108), .Z(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT66), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G2104), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n467), .A2(G137), .A3(new_n468), .A4(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n464), .A2(new_n466), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(G101), .A3(new_n468), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n470), .A2(new_n475), .A3(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n478), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n474), .B1(new_n481), .B2(new_n482), .ZN(G160));
  NAND2_X1  g058(.A1(new_n467), .A2(new_n470), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G136), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n468), .A2(G112), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n467), .A2(new_n470), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n489), .A2(KEYINPUT69), .A3(G2105), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n491), .B1(new_n484), .B2(new_n468), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G124), .ZN(new_n494));
  OAI221_X1 g069(.A(new_n486), .B1(new_n487), .B2(new_n488), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  XNOR2_X1  g070(.A(new_n495), .B(KEYINPUT70), .ZN(G162));
  NAND2_X1  g071(.A1(new_n470), .A2(new_n475), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(new_n468), .A3(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n468), .A2(G138), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n467), .A2(new_n470), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n500), .B1(new_n502), .B2(KEYINPUT4), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n467), .A2(G126), .A3(G2105), .A4(new_n470), .ZN(new_n504));
  OR2_X1    g079(.A1(G102), .A2(G2105), .ZN(new_n505));
  OAI211_X1 g080(.A(new_n505), .B(G2104), .C1(G114), .C2(new_n468), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n503), .A2(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n515), .A2(new_n518), .ZN(G166));
  NAND2_X1  g094(.A1(new_n513), .A2(KEYINPUT71), .ZN(new_n520));
  INV_X1    g095(.A(G543), .ZN(new_n521));
  OR2_X1    g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT71), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n527), .A2(G51), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  XNOR2_X1  g105(.A(KEYINPUT72), .B(G89), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n510), .A2(new_n531), .B1(G63), .B2(G651), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT5), .B(G543), .Z(new_n533));
  OAI21_X1  g108(.A(new_n530), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n528), .A2(new_n534), .ZN(G168));
  AND2_X1   g110(.A1(new_n527), .A2(G52), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n537), .A2(new_n517), .B1(new_n511), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G171));
  XNOR2_X1  g115(.A(KEYINPUT73), .B(G43), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n527), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(G68), .A2(G543), .ZN(new_n543));
  INV_X1    g118(.A(G56), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n543), .B1(new_n533), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n511), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n545), .A2(G651), .B1(new_n546), .B2(G81), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g125(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n551));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  INV_X1    g129(.A(G53), .ZN(new_n555));
  OR3_X1    g130(.A1(new_n513), .A2(KEYINPUT75), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT75), .B1(new_n513), .B2(new_n555), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n556), .A2(KEYINPUT9), .A3(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  OAI211_X1 g134(.A(KEYINPUT75), .B(new_n559), .C1(new_n513), .C2(new_n555), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n533), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n563), .A2(G651), .B1(new_n546), .B2(G91), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n558), .A2(new_n560), .A3(new_n564), .ZN(G299));
  INV_X1    g140(.A(G171), .ZN(G301));
  INV_X1    g141(.A(G168), .ZN(G286));
  INV_X1    g142(.A(G166), .ZN(G303));
  NAND2_X1  g143(.A1(new_n546), .A2(G87), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n524), .A2(G49), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n533), .B2(new_n574), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n575), .A2(G651), .B1(G48), .B2(new_n524), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n577));
  INV_X1    g152(.A(G86), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n511), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n511), .A2(new_n578), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT76), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n576), .A2(new_n579), .A3(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  NOR3_X1   g158(.A1(new_n583), .A2(KEYINPUT77), .A3(new_n517), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(G85), .B2(new_n546), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT77), .B1(new_n583), .B2(new_n517), .ZN(new_n586));
  XOR2_X1   g161(.A(KEYINPUT78), .B(G47), .Z(new_n587));
  NAND2_X1  g162(.A1(new_n527), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(G290));
  AND3_X1   g164(.A1(new_n509), .A2(new_n510), .A3(G92), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n527), .A2(G54), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n593), .A2(new_n517), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(new_n596), .B2(G171), .ZN(G284));
  OAI21_X1  g173(.A(new_n597), .B1(new_n596), .B2(G171), .ZN(G321));
  NOR2_X1   g174(.A1(G286), .A2(new_n596), .ZN(new_n600));
  XNOR2_X1  g175(.A(G299), .B(KEYINPUT79), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(new_n596), .ZN(G297));
  AOI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(new_n596), .ZN(G280));
  AND3_X1   g178(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n604));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n605), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g184(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g185(.A(new_n497), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n611), .A2(new_n468), .A3(new_n472), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT12), .Z(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT13), .ZN(new_n614));
  XOR2_X1   g189(.A(new_n614), .B(G2100), .Z(new_n615));
  AND2_X1   g190(.A1(new_n490), .A2(new_n492), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G123), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT80), .ZN(new_n618));
  OR2_X1    g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n619), .B(G2104), .C1(G111), .C2(new_n468), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n485), .A2(G135), .ZN(new_n621));
  AND3_X1   g196(.A1(new_n618), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT81), .B(G2096), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n615), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(new_n623), .B2(new_n622), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT82), .Z(G156));
  INV_X1    g201(.A(KEYINPUT14), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2427), .B(G2430), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT83), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n629), .B2(new_n630), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n635), .B(new_n637), .Z(new_n638));
  XNOR2_X1  g213(.A(G1341), .B(G1348), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT84), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(G14), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n644), .B1(new_n638), .B2(new_n640), .ZN(new_n645));
  AND2_X1   g220(.A1(new_n643), .A2(new_n645), .ZN(G401));
  XOR2_X1   g221(.A(G2067), .B(G2678), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT85), .ZN(new_n648));
  NOR2_X1   g223(.A1(G2072), .A2(G2078), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n444), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2084), .B(G2090), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  NOR3_X1   g227(.A1(new_n648), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT18), .ZN(new_n654));
  INV_X1    g229(.A(new_n650), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n655), .A2(KEYINPUT86), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(KEYINPUT86), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n656), .A2(new_n648), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n650), .B(KEYINPUT17), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n658), .B(new_n652), .C1(new_n648), .C2(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n659), .A2(new_n648), .A3(new_n651), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n654), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2096), .B(G2100), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(G1971), .B(G1976), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT20), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n668), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n666), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n666), .B2(new_n672), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT87), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1991), .B(G1996), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(G229));
  NOR2_X1   g258(.A1(G29), .A2(G35), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(G162), .B2(G29), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT29), .ZN(new_n686));
  INV_X1    g261(.A(G2090), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G16), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n689), .A2(KEYINPUT90), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n689), .A2(KEYINPUT90), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G20), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT23), .ZN(new_n694));
  AND3_X1   g269(.A1(new_n558), .A2(new_n560), .A3(new_n564), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n694), .B1(new_n695), .B2(new_n689), .ZN(new_n696));
  INV_X1    g271(.A(G1956), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT93), .B(G2067), .ZN(new_n699));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G26), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT28), .Z(new_n702));
  NAND2_X1  g277(.A1(new_n616), .A2(G128), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n468), .A2(G116), .ZN(new_n704));
  OAI21_X1  g279(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  AOI22_X1  g281(.A1(new_n485), .A2(G140), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n702), .B1(new_n708), .B2(G29), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n698), .B1(new_n699), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n689), .A2(G21), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G168), .B2(new_n689), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT102), .B(G1966), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n692), .A2(G19), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(new_n548), .B2(new_n692), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n714), .B1(G1341), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n689), .A2(G5), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G171), .B2(new_n689), .ZN(new_n719));
  INV_X1    g294(.A(G1961), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n716), .A2(G1341), .ZN(new_n722));
  INV_X1    g297(.A(G28), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n723), .A2(KEYINPUT30), .ZN(new_n724));
  AOI21_X1  g299(.A(G29), .B1(new_n723), .B2(KEYINPUT30), .ZN(new_n725));
  OR2_X1    g300(.A1(KEYINPUT31), .A2(G11), .ZN(new_n726));
  NAND2_X1  g301(.A1(KEYINPUT31), .A2(G11), .ZN(new_n727));
  AOI22_X1  g302(.A1(new_n724), .A2(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n721), .A2(new_n722), .A3(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n700), .B1(KEYINPUT24), .B2(G34), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(KEYINPUT24), .B2(G34), .ZN(new_n731));
  INV_X1    g306(.A(G160), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(G29), .ZN(new_n733));
  INV_X1    g308(.A(G2084), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(G27), .A2(G29), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G164), .B2(G29), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G2078), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(G2078), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n735), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NOR4_X1   g315(.A1(new_n710), .A2(new_n717), .A3(new_n729), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n700), .A2(G32), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT100), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT99), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT26), .Z(new_n746));
  NAND3_X1  g321(.A1(new_n472), .A2(G105), .A3(new_n468), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n485), .A2(G141), .ZN(new_n748));
  AND3_X1   g323(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n616), .A2(G129), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT98), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n742), .B1(new_n753), .B2(new_n700), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT27), .B(G1996), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  AND2_X1   g332(.A1(new_n709), .A2(new_n699), .ZN(new_n758));
  NOR2_X1   g333(.A1(G4), .A2(G16), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT92), .Z(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n595), .B2(new_n689), .ZN(new_n761));
  INV_X1    g336(.A(G1348), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  AOI211_X1 g338(.A(new_n758), .B(new_n763), .C1(new_n622), .C2(G29), .ZN(new_n764));
  AND4_X1   g339(.A1(new_n688), .A2(new_n741), .A3(new_n757), .A4(new_n764), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n689), .A2(G6), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G305), .B2(G16), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT91), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT32), .B(G1981), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n689), .A2(G23), .ZN(new_n772));
  INV_X1    g347(.A(G288), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n689), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT33), .B(G1976), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n692), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(G22), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(G166), .B2(new_n777), .ZN(new_n779));
  XOR2_X1   g354(.A(new_n779), .B(G1971), .Z(new_n780));
  NAND4_X1  g355(.A1(new_n770), .A2(new_n771), .A3(new_n776), .A4(new_n780), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT34), .Z(new_n782));
  INV_X1    g357(.A(KEYINPUT36), .ZN(new_n783));
  MUX2_X1   g358(.A(G24), .B(G290), .S(new_n777), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(G1986), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n700), .A2(G25), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT88), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n616), .A2(G119), .ZN(new_n788));
  NOR2_X1   g363(.A1(G95), .A2(G2105), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT89), .Z(new_n790));
  INV_X1    g365(.A(G107), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n463), .B1(new_n791), .B2(G2105), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n485), .A2(G131), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n788), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n787), .B1(new_n794), .B2(G29), .ZN(new_n795));
  XOR2_X1   g370(.A(KEYINPUT35), .B(G1991), .Z(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n785), .A2(new_n797), .ZN(new_n798));
  AND3_X1   g373(.A1(new_n782), .A2(new_n783), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n783), .B1(new_n782), .B2(new_n798), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n765), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT97), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n485), .A2(G139), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT25), .Z(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT94), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n611), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n809), .A2(new_n468), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(KEYINPUT95), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT95), .ZN(new_n813));
  NAND3_X1  g388(.A1(new_n808), .A2(new_n813), .A3(new_n810), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(G29), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n700), .A2(G33), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT96), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n802), .B1(new_n819), .B2(G2072), .ZN(new_n820));
  OAI22_X1  g395(.A1(new_n754), .A2(new_n756), .B1(new_n734), .B2(new_n733), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(new_n819), .B2(G2072), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT96), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n818), .B(new_n823), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n824), .A2(KEYINPUT97), .A3(new_n442), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n820), .A2(new_n822), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(KEYINPUT101), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT101), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n820), .A2(new_n822), .A3(new_n828), .A4(new_n825), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n801), .B1(new_n827), .B2(new_n829), .ZN(G311));
  NAND2_X1  g405(.A1(new_n827), .A2(new_n829), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n799), .A2(new_n800), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n831), .A2(new_n832), .A3(new_n765), .ZN(G150));
  NAND2_X1  g408(.A1(new_n604), .A2(G559), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT38), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n527), .A2(G55), .ZN(new_n836));
  AOI22_X1  g411(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n837), .A2(new_n517), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT103), .B(G93), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n546), .A2(new_n839), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n548), .A2(new_n836), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n836), .A2(new_n838), .A3(new_n840), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n542), .A2(new_n547), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n835), .B(new_n846), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n847), .A2(KEYINPUT39), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(KEYINPUT39), .ZN(new_n849));
  NOR3_X1   g424(.A1(new_n848), .A2(new_n849), .A3(G860), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n843), .A2(G860), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT37), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n850), .A2(new_n852), .ZN(G145));
  AND2_X1   g428(.A1(new_n504), .A2(new_n506), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT104), .ZN(new_n855));
  AND2_X1   g430(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n854), .B(new_n855), .C1(new_n856), .C2(new_n500), .ZN(new_n857));
  OAI21_X1  g432(.A(KEYINPUT104), .B1(new_n503), .B2(new_n507), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n708), .B(new_n859), .Z(new_n860));
  NAND4_X1  g435(.A1(new_n812), .A2(new_n749), .A3(new_n814), .A4(new_n751), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  AOI22_X1  g437(.A1(new_n812), .A2(new_n814), .B1(new_n749), .B2(new_n751), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n860), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n863), .ZN(new_n865));
  INV_X1    g440(.A(new_n860), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n865), .A2(new_n861), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT106), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n788), .A2(new_n793), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(KEYINPUT105), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT105), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n794), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n613), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n616), .A2(G130), .ZN(new_n876));
  OR2_X1    g451(.A1(new_n468), .A2(G118), .ZN(new_n877));
  OAI21_X1  g452(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  AOI22_X1  g454(.A1(new_n485), .A2(G142), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n613), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n871), .A2(new_n883), .A3(new_n873), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n875), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n882), .B1(new_n875), .B2(new_n884), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n869), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n868), .A2(new_n888), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n886), .A2(new_n887), .A3(new_n869), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n875), .A2(new_n884), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n881), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT106), .B1(new_n892), .B2(new_n885), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n889), .B1(new_n894), .B2(new_n868), .ZN(new_n895));
  XNOR2_X1  g470(.A(G162), .B(G160), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n622), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(G37), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n897), .B(new_n889), .C1(new_n894), .C2(new_n868), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT40), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n892), .A2(KEYINPUT106), .A3(new_n885), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n868), .B1(new_n902), .B2(new_n888), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n868), .A2(new_n888), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n898), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  AND4_X1   g481(.A1(KEYINPUT40), .A2(new_n905), .A3(new_n900), .A4(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n901), .A2(new_n907), .ZN(G395));
  NAND2_X1  g483(.A1(new_n842), .A2(new_n845), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(new_n607), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT107), .B1(new_n604), .B2(G299), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n604), .A2(G299), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n695), .A2(new_n595), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n912), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n910), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT41), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n911), .A2(KEYINPUT41), .A3(new_n914), .A4(new_n912), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n916), .B1(new_n920), .B2(new_n910), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n921), .A2(KEYINPUT42), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(KEYINPUT42), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(G166), .B(KEYINPUT108), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(G305), .ZN(new_n926));
  XNOR2_X1  g501(.A(G290), .B(new_n773), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n926), .B(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n596), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n928), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n922), .A2(new_n930), .A3(new_n923), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n929), .A2(KEYINPUT109), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n929), .A2(new_n931), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT109), .B1(new_n843), .B2(new_n596), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(G295));
  AOI21_X1  g510(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(G331));
  NAND2_X1  g511(.A1(new_n846), .A2(G301), .ZN(new_n937));
  AOI21_X1  g512(.A(G301), .B1(new_n842), .B2(new_n845), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n937), .A2(G168), .A3(new_n939), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n909), .A2(G171), .ZN(new_n941));
  OAI21_X1  g516(.A(G286), .B1(new_n941), .B2(new_n938), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(new_n915), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n918), .A2(new_n919), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(new_n940), .A3(new_n942), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n928), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n906), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n928), .B1(new_n944), .B2(new_n946), .ZN(new_n949));
  OR3_X1    g524(.A1(new_n948), .A2(KEYINPUT43), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n940), .B(new_n942), .C1(KEYINPUT110), .C2(new_n919), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n918), .A2(KEYINPUT110), .A3(new_n919), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n944), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n948), .B1(new_n930), .B2(new_n954), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n950), .B(KEYINPUT44), .C1(new_n951), .C2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT111), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n954), .A2(new_n930), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n958), .A2(new_n951), .A3(new_n906), .A4(new_n947), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT43), .B1(new_n948), .B2(new_n949), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n957), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI211_X1 g538(.A(KEYINPUT111), .B(KEYINPUT44), .C1(new_n959), .C2(new_n960), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n956), .B1(new_n963), .B2(new_n964), .ZN(G397));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n857), .A2(new_n966), .A3(new_n858), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n471), .A2(new_n473), .ZN(new_n970));
  AOI21_X1  g545(.A(KEYINPUT67), .B1(new_n478), .B2(G2105), .ZN(new_n971));
  AOI211_X1 g546(.A(new_n480), .B(new_n468), .C1(new_n476), .C2(new_n477), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n970), .B(G40), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n969), .A2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n708), .A2(G2067), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT112), .ZN(new_n977));
  INV_X1    g552(.A(G2067), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n703), .B2(new_n707), .ZN(new_n979));
  OR3_X1    g554(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n977), .B1(new_n976), .B2(new_n979), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n975), .B1(new_n982), .B2(new_n753), .ZN(new_n983));
  INV_X1    g558(.A(G1996), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n975), .ZN(new_n987));
  NOR2_X1   g562(.A1(G290), .A2(G1986), .ZN(new_n988));
  AND2_X1   g563(.A1(G290), .A2(G1986), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n984), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(new_n752), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n794), .B(new_n796), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT113), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n987), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n986), .A2(new_n990), .A3(new_n993), .A4(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(KEYINPUT115), .B(G8), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n966), .B1(new_n503), .B2(new_n507), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n973), .B1(new_n968), .B2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n857), .A2(KEYINPUT45), .A3(new_n966), .A4(new_n858), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1971), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1004), .B(new_n966), .C1(new_n503), .C2(new_n507), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1000), .A2(KEYINPUT50), .ZN(new_n1006));
  AND4_X1   g581(.A1(new_n687), .A2(new_n974), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n999), .B1(new_n1003), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n1009));
  INV_X1    g584(.A(G8), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1009), .B1(G166), .B2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g586(.A(KEYINPUT55), .B(G8), .C1(new_n515), .C2(new_n518), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1008), .A2(new_n1013), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1011), .A2(KEYINPUT114), .A3(new_n1012), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT114), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n1017), .B(G8), .C1(new_n1003), .C2(new_n1007), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n999), .B1(new_n973), .B2(new_n1000), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n773), .A2(G1976), .ZN(new_n1021));
  INV_X1    g596(.A(G1976), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(G288), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1981), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n576), .A2(new_n581), .A3(new_n1025), .A4(new_n579), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n524), .A2(G48), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1027), .B1(new_n1028), .B2(new_n517), .ZN(new_n1029));
  OAI21_X1  g604(.A(G1981), .B1(new_n1029), .B2(new_n580), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT49), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1026), .A2(KEYINPUT49), .A3(new_n1030), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1020), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(G288), .A2(new_n1022), .ZN(new_n1036));
  OAI21_X1  g611(.A(KEYINPUT52), .B1(new_n1019), .B2(new_n1036), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1024), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1000), .A2(new_n968), .ZN(new_n1039));
  OAI211_X1 g614(.A(KEYINPUT45), .B(new_n966), .C1(new_n503), .C2(new_n507), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n974), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(G1966), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT117), .B(G2084), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n974), .A2(new_n1006), .A3(new_n1005), .A4(new_n1044), .ZN(new_n1045));
  AOI211_X1 g620(.A(G286), .B(new_n998), .C1(new_n1043), .C2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1014), .A2(new_n1018), .A3(new_n1038), .A4(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT63), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n974), .A2(new_n1006), .A3(new_n1005), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  AOI22_X1  g626(.A1(new_n1051), .A2(new_n1044), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1052));
  NOR4_X1   g627(.A1(new_n1052), .A2(new_n1048), .A3(G286), .A4(new_n998), .ZN(new_n1053));
  OAI21_X1  g628(.A(G8), .B1(new_n1003), .B2(new_n1007), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(new_n1013), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1053), .A2(new_n1018), .A3(new_n1038), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1049), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1026), .ZN(new_n1058));
  NOR2_X1   g633(.A1(G288), .A2(G1976), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1058), .B1(new_n1035), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1020), .B1(new_n1060), .B2(KEYINPUT116), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1060), .A2(KEYINPUT116), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1018), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1062), .A2(new_n1063), .B1(new_n1064), .B2(new_n1038), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1057), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1067), .B1(new_n1052), .B2(new_n998), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1069), .A2(KEYINPUT122), .A3(new_n999), .ZN(new_n1070));
  NOR2_X1   g645(.A1(G168), .A2(new_n998), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1071), .A2(KEYINPUT51), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1068), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(KEYINPUT121), .B(KEYINPUT51), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1010), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1074), .B1(new_n1075), .B2(new_n1071), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1073), .A2(new_n1076), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT62), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n443), .A2(KEYINPUT53), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1001), .A2(new_n1081), .A3(new_n1040), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1050), .A2(new_n720), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1001), .A2(new_n443), .A3(new_n1002), .ZN(new_n1085));
  XOR2_X1   g660(.A(KEYINPUT123), .B(KEYINPUT53), .Z(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(G301), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1088), .A2(new_n1014), .A3(new_n1018), .A4(new_n1038), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT122), .B1(new_n1069), .B2(new_n999), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1076), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1089), .B1(new_n1094), .B2(KEYINPUT62), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1066), .B1(new_n1079), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT57), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n695), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1050), .A2(new_n697), .ZN(new_n1101));
  XNOR2_X1  g676(.A(KEYINPUT56), .B(G2072), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1001), .A2(new_n1002), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1100), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  NOR3_X1   g679(.A1(new_n973), .A2(new_n1000), .A3(G2067), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1105), .B1(new_n1050), .B2(new_n762), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1106), .A2(new_n595), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1104), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1103), .A2(new_n1101), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1111), .A2(new_n1104), .A3(KEYINPUT61), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1113), .A2(KEYINPUT119), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1001), .A2(new_n984), .A3(new_n1002), .ZN(new_n1115));
  XOR2_X1   g690(.A(KEYINPUT58), .B(G1341), .Z(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(new_n973), .B2(new_n1000), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT118), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT118), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1119), .B(new_n1116), .C1(new_n973), .C2(new_n1000), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1115), .A2(new_n1118), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(new_n548), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(KEYINPUT59), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1121), .A2(new_n1124), .A3(new_n548), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1123), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1111), .A2(new_n1104), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1114), .A2(new_n1126), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1111), .A2(new_n1104), .A3(new_n1131), .A4(KEYINPUT61), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1050), .A2(new_n762), .ZN(new_n1133));
  INV_X1    g708(.A(new_n1105), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n595), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1133), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT120), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n595), .A2(new_n1135), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1106), .A2(KEYINPUT120), .A3(new_n1136), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1139), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1141), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1132), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1112), .B1(new_n1130), .B2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n970), .A2(G40), .A3(new_n479), .A4(new_n1081), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1147), .B1(new_n967), .B2(new_n968), .ZN(new_n1148));
  AOI22_X1  g723(.A1(new_n1148), .A2(new_n1002), .B1(new_n720), .B2(new_n1050), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(new_n1087), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT124), .B1(new_n1150), .B2(G171), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1084), .A2(new_n1087), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(G171), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1149), .A2(new_n1154), .A3(G301), .A4(new_n1087), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1151), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT54), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1087), .A2(new_n1082), .A3(G301), .A4(new_n1083), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT54), .ZN(new_n1160));
  AOI21_X1  g735(.A(G301), .B1(new_n1149), .B2(new_n1087), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT125), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1150), .A2(G171), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1163), .A2(new_n1164), .A3(KEYINPUT54), .A4(new_n1159), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1014), .A2(new_n1018), .A3(new_n1038), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1167), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1146), .A2(new_n1158), .A3(new_n1166), .A4(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n997), .B1(new_n1096), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n870), .A2(new_n796), .ZN(new_n1171));
  AOI211_X1 g746(.A(new_n1171), .B(new_n992), .C1(new_n983), .C2(new_n985), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n987), .B1(new_n1172), .B2(new_n976), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n987), .A2(new_n988), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT48), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n986), .A2(new_n993), .A3(new_n996), .A4(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT47), .ZN(new_n1177));
  AOI21_X1  g752(.A(KEYINPUT46), .B1(new_n987), .B2(new_n984), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n983), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n987), .A2(KEYINPUT46), .A3(new_n984), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1180), .B(KEYINPUT126), .ZN(new_n1181));
  AOI21_X1  g756(.A(new_n1177), .B1(new_n1179), .B2(new_n1181), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1179), .A2(new_n1177), .A3(new_n1181), .ZN(new_n1183));
  OAI211_X1 g758(.A(new_n1173), .B(new_n1176), .C1(new_n1182), .C2(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(KEYINPUT127), .B1(new_n1170), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n997), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1112), .ZN(new_n1187));
  AND3_X1   g762(.A1(new_n1114), .A2(new_n1126), .A3(new_n1129), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1113), .ZN(new_n1189));
  INV_X1    g764(.A(new_n1142), .ZN(new_n1190));
  AOI21_X1  g765(.A(KEYINPUT120), .B1(new_n1106), .B2(new_n1136), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1140), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1139), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1193));
  AOI22_X1  g768(.A1(new_n1189), .A2(new_n1131), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1187), .B1(new_n1188), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1168), .A2(new_n1158), .A3(new_n1166), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1064), .A2(new_n1038), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1063), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1198), .B1(new_n1199), .B2(new_n1061), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1200), .B1(new_n1049), .B2(new_n1056), .ZN(new_n1201));
  INV_X1    g776(.A(new_n1089), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1202), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1094), .A2(KEYINPUT62), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1201), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1186), .B1(new_n1197), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1176), .B1(new_n1183), .B2(new_n1182), .ZN(new_n1207));
  NAND4_X1  g782(.A1(new_n986), .A2(new_n796), .A3(new_n870), .A4(new_n993), .ZN(new_n1208));
  INV_X1    g783(.A(new_n976), .ZN(new_n1209));
  AOI21_X1  g784(.A(new_n975), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g785(.A1(new_n1207), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n1212));
  NAND3_X1  g787(.A1(new_n1206), .A2(new_n1211), .A3(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1185), .A2(new_n1213), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g789(.A1(new_n899), .A2(new_n900), .ZN(new_n1216));
  INV_X1    g790(.A(G319), .ZN(new_n1217));
  NOR2_X1   g791(.A1(G227), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g792(.A1(new_n682), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g793(.A(new_n1219), .B1(new_n643), .B2(new_n645), .ZN(new_n1220));
  AND3_X1   g794(.A1(new_n1216), .A2(new_n1220), .A3(new_n961), .ZN(G308));
  NAND3_X1  g795(.A1(new_n1216), .A2(new_n1220), .A3(new_n961), .ZN(G225));
endmodule


