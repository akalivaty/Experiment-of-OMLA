

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U550 ( .A1(n546), .A2(n545), .ZN(G160) );
  NOR2_X2 U551 ( .A1(n710), .A2(n709), .ZN(n716) );
  NOR2_X2 U552 ( .A1(G168), .A2(n689), .ZN(n690) );
  XNOR2_X1 U553 ( .A(n533), .B(KEYINPUT23), .ZN(n534) );
  INV_X1 U554 ( .A(KEYINPUT64), .ZN(n533) );
  AND2_X1 U555 ( .A1(n687), .A2(n738), .ZN(n688) );
  XNOR2_X1 U556 ( .A(n542), .B(n541), .ZN(n556) );
  XNOR2_X1 U557 ( .A(n540), .B(KEYINPUT17), .ZN(n542) );
  INV_X1 U558 ( .A(KEYINPUT66), .ZN(n540) );
  XNOR2_X1 U559 ( .A(n593), .B(KEYINPUT73), .ZN(n703) );
  OR2_X1 U560 ( .A1(n897), .A2(n712), .ZN(n516) );
  XOR2_X1 U561 ( .A(KEYINPUT32), .B(n734), .Z(n517) );
  NOR2_X2 U562 ( .A1(n769), .A2(n770), .ZN(n708) );
  NOR2_X1 U563 ( .A1(G2084), .A2(n727), .ZN(n736) );
  XNOR2_X1 U564 ( .A(KEYINPUT13), .B(KEYINPUT72), .ZN(n587) );
  XNOR2_X1 U565 ( .A(n588), .B(n587), .ZN(n590) );
  INV_X1 U566 ( .A(KEYINPUT87), .ZN(n557) );
  XNOR2_X1 U567 ( .A(n558), .B(n557), .ZN(n560) );
  NOR2_X1 U568 ( .A1(n627), .A2(n525), .ZN(n642) );
  BUF_X1 U569 ( .A(n556), .Z(n875) );
  XOR2_X1 U570 ( .A(KEYINPUT1), .B(n519), .Z(n646) );
  XNOR2_X1 U571 ( .A(n535), .B(n534), .ZN(n538) );
  INV_X1 U572 ( .A(n703), .ZN(n995) );
  XOR2_X1 U573 ( .A(G543), .B(KEYINPUT0), .Z(n627) );
  NOR2_X1 U574 ( .A1(G651), .A2(n627), .ZN(n647) );
  NAND2_X1 U575 ( .A1(n647), .A2(G51), .ZN(n518) );
  XNOR2_X1 U576 ( .A(n518), .B(KEYINPUT76), .ZN(n521) );
  XNOR2_X1 U577 ( .A(KEYINPUT67), .B(G651), .ZN(n525) );
  NOR2_X1 U578 ( .A1(G543), .A2(n525), .ZN(n519) );
  NAND2_X1 U579 ( .A1(G63), .A2(n646), .ZN(n520) );
  NAND2_X1 U580 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U581 ( .A(KEYINPUT6), .B(n522), .ZN(n530) );
  NOR2_X1 U582 ( .A1(G651), .A2(G543), .ZN(n641) );
  NAND2_X1 U583 ( .A1(G89), .A2(n641), .ZN(n523) );
  XOR2_X1 U584 ( .A(KEYINPUT4), .B(n523), .Z(n524) );
  XNOR2_X1 U585 ( .A(n524), .B(KEYINPUT75), .ZN(n527) );
  NAND2_X1 U586 ( .A1(G76), .A2(n642), .ZN(n526) );
  NAND2_X1 U587 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U588 ( .A(KEYINPUT5), .B(n528), .Z(n529) );
  NOR2_X1 U589 ( .A1(n530), .A2(n529), .ZN(n532) );
  XNOR2_X1 U590 ( .A(KEYINPUT7), .B(KEYINPUT77), .ZN(n531) );
  XNOR2_X1 U591 ( .A(n532), .B(n531), .ZN(G168) );
  XOR2_X1 U592 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U593 ( .A(G2105), .ZN(n539) );
  AND2_X2 U594 ( .A1(n539), .A2(G2104), .ZN(n877) );
  NAND2_X1 U595 ( .A1(G101), .A2(n877), .ZN(n535) );
  NAND2_X1 U596 ( .A1(G2105), .A2(G2104), .ZN(n536) );
  XNOR2_X1 U597 ( .A(n536), .B(KEYINPUT65), .ZN(n871) );
  NAND2_X1 U598 ( .A1(G113), .A2(n871), .ZN(n537) );
  NAND2_X1 U599 ( .A1(n538), .A2(n537), .ZN(n546) );
  NOR2_X1 U600 ( .A1(G2104), .A2(n539), .ZN(n872) );
  NAND2_X1 U601 ( .A1(n872), .A2(G125), .ZN(n544) );
  NOR2_X1 U602 ( .A1(G2104), .A2(G2105), .ZN(n541) );
  NAND2_X1 U603 ( .A1(G137), .A2(n875), .ZN(n543) );
  NAND2_X1 U604 ( .A1(n544), .A2(n543), .ZN(n545) );
  AND2_X1 U605 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U606 ( .A1(G111), .A2(n871), .ZN(n547) );
  XNOR2_X1 U607 ( .A(n547), .B(KEYINPUT78), .ZN(n554) );
  NAND2_X1 U608 ( .A1(n877), .A2(G99), .ZN(n549) );
  NAND2_X1 U609 ( .A1(G135), .A2(n875), .ZN(n548) );
  NAND2_X1 U610 ( .A1(n549), .A2(n548), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n872), .A2(G123), .ZN(n550) );
  XOR2_X1 U612 ( .A(KEYINPUT18), .B(n550), .Z(n551) );
  NOR2_X1 U613 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U614 ( .A1(n554), .A2(n553), .ZN(n927) );
  XNOR2_X1 U615 ( .A(G2096), .B(n927), .ZN(n555) );
  OR2_X1 U616 ( .A1(G2100), .A2(n555), .ZN(G156) );
  NAND2_X1 U617 ( .A1(G138), .A2(n556), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n877), .A2(G102), .ZN(n559) );
  NAND2_X1 U619 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U620 ( .A(n561), .B(KEYINPUT88), .ZN(n565) );
  NAND2_X1 U621 ( .A1(G114), .A2(n871), .ZN(n563) );
  NAND2_X1 U622 ( .A1(G126), .A2(n872), .ZN(n562) );
  NAND2_X1 U623 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U624 ( .A1(n565), .A2(n564), .ZN(n681) );
  BUF_X1 U625 ( .A(n681), .Z(G164) );
  INV_X1 U626 ( .A(G132), .ZN(G219) );
  INV_X1 U627 ( .A(G82), .ZN(G220) );
  INV_X1 U628 ( .A(G57), .ZN(G237) );
  INV_X1 U629 ( .A(G108), .ZN(G238) );
  INV_X1 U630 ( .A(G120), .ZN(G236) );
  NAND2_X1 U631 ( .A1(n641), .A2(G88), .ZN(n567) );
  NAND2_X1 U632 ( .A1(G75), .A2(n642), .ZN(n566) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n647), .A2(G50), .ZN(n569) );
  NAND2_X1 U635 ( .A1(G62), .A2(n646), .ZN(n568) );
  NAND2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(G166) );
  NAND2_X1 U638 ( .A1(n647), .A2(G52), .ZN(n573) );
  NAND2_X1 U639 ( .A1(G64), .A2(n646), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n578) );
  NAND2_X1 U641 ( .A1(n641), .A2(G90), .ZN(n575) );
  NAND2_X1 U642 ( .A1(G77), .A2(n642), .ZN(n574) );
  NAND2_X1 U643 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U644 ( .A(KEYINPUT9), .B(n576), .Z(n577) );
  NOR2_X1 U645 ( .A1(n578), .A2(n577), .ZN(G171) );
  INV_X1 U646 ( .A(G171), .ZN(G301) );
  NAND2_X1 U647 ( .A1(G7), .A2(G661), .ZN(n579) );
  XOR2_X1 U648 ( .A(n579), .B(KEYINPUT10), .Z(n918) );
  NAND2_X1 U649 ( .A1(n918), .A2(G567), .ZN(n580) );
  XOR2_X1 U650 ( .A(KEYINPUT11), .B(n580), .Z(G234) );
  XOR2_X1 U651 ( .A(KEYINPUT70), .B(KEYINPUT14), .Z(n582) );
  NAND2_X1 U652 ( .A1(G56), .A2(n646), .ZN(n581) );
  XNOR2_X1 U653 ( .A(n582), .B(n581), .ZN(n592) );
  NAND2_X1 U654 ( .A1(n642), .A2(G68), .ZN(n586) );
  XOR2_X1 U655 ( .A(KEYINPUT71), .B(KEYINPUT12), .Z(n584) );
  NAND2_X1 U656 ( .A1(G81), .A2(n641), .ZN(n583) );
  XNOR2_X1 U657 ( .A(n584), .B(n583), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U659 ( .A1(G43), .A2(n647), .ZN(n589) );
  NAND2_X1 U660 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U661 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U662 ( .A1(n995), .A2(G860), .ZN(G153) );
  NAND2_X1 U663 ( .A1(G92), .A2(n641), .ZN(n595) );
  NAND2_X1 U664 ( .A1(G54), .A2(n647), .ZN(n594) );
  NAND2_X1 U665 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U666 ( .A1(G79), .A2(n642), .ZN(n597) );
  NAND2_X1 U667 ( .A1(G66), .A2(n646), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U669 ( .A1(n599), .A2(n598), .ZN(n601) );
  XNOR2_X1 U670 ( .A(KEYINPUT74), .B(KEYINPUT15), .ZN(n600) );
  XOR2_X1 U671 ( .A(n601), .B(n600), .Z(n997) );
  INV_X1 U672 ( .A(n997), .ZN(n897) );
  NOR2_X1 U673 ( .A1(n897), .A2(G868), .ZN(n603) );
  INV_X1 U674 ( .A(G868), .ZN(n660) );
  NOR2_X1 U675 ( .A1(n660), .A2(G301), .ZN(n602) );
  NOR2_X1 U676 ( .A1(n603), .A2(n602), .ZN(G284) );
  NAND2_X1 U677 ( .A1(n647), .A2(G53), .ZN(n605) );
  NAND2_X1 U678 ( .A1(G65), .A2(n646), .ZN(n604) );
  NAND2_X1 U679 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U680 ( .A1(n641), .A2(G91), .ZN(n607) );
  NAND2_X1 U681 ( .A1(G78), .A2(n642), .ZN(n606) );
  NAND2_X1 U682 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U683 ( .A1(n609), .A2(n608), .ZN(n1002) );
  XNOR2_X1 U684 ( .A(n1002), .B(KEYINPUT69), .ZN(G299) );
  NAND2_X1 U685 ( .A1(G286), .A2(G868), .ZN(n611) );
  NAND2_X1 U686 ( .A1(n660), .A2(G299), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n611), .A2(n610), .ZN(G297) );
  INV_X1 U688 ( .A(G860), .ZN(n618) );
  NAND2_X1 U689 ( .A1(n618), .A2(G559), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n612), .A2(n997), .ZN(n613) );
  XNOR2_X1 U691 ( .A(n613), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U692 ( .A1(n897), .A2(G559), .ZN(n614) );
  NOR2_X1 U693 ( .A1(n660), .A2(n614), .ZN(n616) );
  NOR2_X1 U694 ( .A1(n995), .A2(G868), .ZN(n615) );
  OR2_X1 U695 ( .A1(n616), .A2(n615), .ZN(G282) );
  NAND2_X1 U696 ( .A1(n997), .A2(G559), .ZN(n617) );
  XNOR2_X1 U697 ( .A(n617), .B(n995), .ZN(n657) );
  NAND2_X1 U698 ( .A1(n618), .A2(n657), .ZN(n626) );
  NAND2_X1 U699 ( .A1(G93), .A2(n641), .ZN(n620) );
  NAND2_X1 U700 ( .A1(G55), .A2(n647), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n620), .A2(n619), .ZN(n623) );
  NAND2_X1 U702 ( .A1(G67), .A2(n646), .ZN(n621) );
  XNOR2_X1 U703 ( .A(KEYINPUT79), .B(n621), .ZN(n622) );
  NOR2_X1 U704 ( .A1(n623), .A2(n622), .ZN(n625) );
  NAND2_X1 U705 ( .A1(G80), .A2(n642), .ZN(n624) );
  NAND2_X1 U706 ( .A1(n625), .A2(n624), .ZN(n661) );
  XNOR2_X1 U707 ( .A(n626), .B(n661), .ZN(G145) );
  NAND2_X1 U708 ( .A1(G87), .A2(n627), .ZN(n629) );
  NAND2_X1 U709 ( .A1(G74), .A2(G651), .ZN(n628) );
  NAND2_X1 U710 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U711 ( .A1(n646), .A2(n630), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n647), .A2(G49), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n632), .A2(n631), .ZN(G288) );
  XOR2_X1 U714 ( .A(KEYINPUT80), .B(KEYINPUT2), .Z(n634) );
  NAND2_X1 U715 ( .A1(G73), .A2(n642), .ZN(n633) );
  XNOR2_X1 U716 ( .A(n634), .B(n633), .ZN(n638) );
  NAND2_X1 U717 ( .A1(G86), .A2(n641), .ZN(n636) );
  NAND2_X1 U718 ( .A1(G48), .A2(n647), .ZN(n635) );
  NAND2_X1 U719 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U720 ( .A1(n638), .A2(n637), .ZN(n640) );
  NAND2_X1 U721 ( .A1(G61), .A2(n646), .ZN(n639) );
  NAND2_X1 U722 ( .A1(n640), .A2(n639), .ZN(G305) );
  NAND2_X1 U723 ( .A1(n641), .A2(G85), .ZN(n644) );
  NAND2_X1 U724 ( .A1(G72), .A2(n642), .ZN(n643) );
  NAND2_X1 U725 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U726 ( .A(KEYINPUT68), .B(n645), .Z(n651) );
  NAND2_X1 U727 ( .A1(n646), .A2(G60), .ZN(n649) );
  NAND2_X1 U728 ( .A1(n647), .A2(G47), .ZN(n648) );
  AND2_X1 U729 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(G290) );
  XOR2_X1 U731 ( .A(KEYINPUT19), .B(G166), .Z(n652) );
  XNOR2_X1 U732 ( .A(n652), .B(G288), .ZN(n653) );
  XNOR2_X1 U733 ( .A(n653), .B(G305), .ZN(n654) );
  XNOR2_X1 U734 ( .A(n654), .B(n661), .ZN(n655) );
  XNOR2_X1 U735 ( .A(n655), .B(G290), .ZN(n656) );
  XNOR2_X1 U736 ( .A(n656), .B(G299), .ZN(n896) );
  XNOR2_X1 U737 ( .A(n896), .B(n657), .ZN(n658) );
  NAND2_X1 U738 ( .A1(n658), .A2(G868), .ZN(n659) );
  XOR2_X1 U739 ( .A(KEYINPUT81), .B(n659), .Z(n663) );
  NAND2_X1 U740 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U741 ( .A1(n663), .A2(n662), .ZN(G295) );
  NAND2_X1 U742 ( .A1(G2078), .A2(G2084), .ZN(n664) );
  XOR2_X1 U743 ( .A(KEYINPUT20), .B(n664), .Z(n665) );
  NAND2_X1 U744 ( .A1(n665), .A2(G2090), .ZN(n666) );
  XNOR2_X1 U745 ( .A(n666), .B(KEYINPUT82), .ZN(n667) );
  XNOR2_X1 U746 ( .A(KEYINPUT21), .B(n667), .ZN(n668) );
  NAND2_X1 U747 ( .A1(n668), .A2(G2072), .ZN(n669) );
  XOR2_X1 U748 ( .A(KEYINPUT83), .B(n669), .Z(G158) );
  XNOR2_X1 U749 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U750 ( .A1(G236), .A2(G238), .ZN(n670) );
  NAND2_X1 U751 ( .A1(G69), .A2(n670), .ZN(n671) );
  NOR2_X1 U752 ( .A1(n671), .A2(G237), .ZN(n672) );
  XNOR2_X1 U753 ( .A(n672), .B(KEYINPUT85), .ZN(n827) );
  NAND2_X1 U754 ( .A1(n827), .A2(G567), .ZN(n678) );
  NOR2_X1 U755 ( .A1(G220), .A2(G219), .ZN(n673) );
  XNOR2_X1 U756 ( .A(KEYINPUT22), .B(n673), .ZN(n674) );
  NAND2_X1 U757 ( .A1(n674), .A2(G96), .ZN(n675) );
  NOR2_X1 U758 ( .A1(G218), .A2(n675), .ZN(n676) );
  XOR2_X1 U759 ( .A(KEYINPUT84), .B(n676), .Z(n826) );
  NAND2_X1 U760 ( .A1(n826), .A2(G2106), .ZN(n677) );
  NAND2_X1 U761 ( .A1(n678), .A2(n677), .ZN(n829) );
  NAND2_X1 U762 ( .A1(G661), .A2(G483), .ZN(n679) );
  XNOR2_X1 U763 ( .A(KEYINPUT86), .B(n679), .ZN(n680) );
  NOR2_X1 U764 ( .A1(n829), .A2(n680), .ZN(n825) );
  NAND2_X1 U765 ( .A1(n825), .A2(G36), .ZN(G176) );
  INV_X1 U766 ( .A(G166), .ZN(G303) );
  INV_X1 U767 ( .A(G8), .ZN(n682) );
  OR2_X2 U768 ( .A1(n681), .A2(G1384), .ZN(n769) );
  NAND2_X1 U769 ( .A1(G160), .A2(G40), .ZN(n770) );
  OR2_X4 U770 ( .A1(n769), .A2(n770), .ZN(n727) );
  NOR2_X1 U771 ( .A1(n682), .A2(n736), .ZN(n687) );
  INV_X1 U772 ( .A(G1966), .ZN(n683) );
  AND2_X1 U773 ( .A1(n683), .A2(G8), .ZN(n684) );
  NAND2_X1 U774 ( .A1(n727), .A2(n684), .ZN(n686) );
  INV_X1 U775 ( .A(KEYINPUT97), .ZN(n685) );
  XNOR2_X1 U776 ( .A(n686), .B(n685), .ZN(n738) );
  XOR2_X1 U777 ( .A(n688), .B(KEYINPUT30), .Z(n689) );
  XNOR2_X1 U778 ( .A(n690), .B(KEYINPUT101), .ZN(n694) );
  XOR2_X1 U779 ( .A(G2078), .B(KEYINPUT25), .Z(n973) );
  NOR2_X1 U780 ( .A1(n973), .A2(n727), .ZN(n692) );
  NOR2_X1 U781 ( .A1(n708), .A2(G1961), .ZN(n691) );
  NOR2_X1 U782 ( .A1(n692), .A2(n691), .ZN(n721) );
  NAND2_X1 U783 ( .A1(n721), .A2(G301), .ZN(n693) );
  NAND2_X1 U784 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U785 ( .A(n695), .B(KEYINPUT31), .ZN(n725) );
  NAND2_X1 U786 ( .A1(n727), .A2(G1341), .ZN(n696) );
  XNOR2_X1 U787 ( .A(n696), .B(KEYINPUT98), .ZN(n701) );
  NAND2_X1 U788 ( .A1(G1348), .A2(n727), .ZN(n697) );
  XOR2_X1 U789 ( .A(KEYINPUT99), .B(n697), .Z(n699) );
  NAND2_X1 U790 ( .A1(G2067), .A2(n708), .ZN(n698) );
  NAND2_X1 U791 ( .A1(n699), .A2(n698), .ZN(n712) );
  NAND2_X1 U792 ( .A1(n712), .A2(n897), .ZN(n700) );
  AND2_X1 U793 ( .A1(n701), .A2(n700), .ZN(n706) );
  NAND2_X1 U794 ( .A1(G1996), .A2(n708), .ZN(n702) );
  XOR2_X1 U795 ( .A(KEYINPUT26), .B(n702), .Z(n704) );
  NOR2_X1 U796 ( .A1(n704), .A2(n703), .ZN(n705) );
  AND2_X1 U797 ( .A1(n706), .A2(n705), .ZN(n715) );
  NAND2_X1 U798 ( .A1(n708), .A2(G2072), .ZN(n707) );
  XNOR2_X1 U799 ( .A(n707), .B(KEYINPUT27), .ZN(n710) );
  INV_X1 U800 ( .A(G1956), .ZN(n1003) );
  NOR2_X1 U801 ( .A1(n1003), .A2(n708), .ZN(n709) );
  NAND2_X1 U802 ( .A1(n716), .A2(n1002), .ZN(n711) );
  XNOR2_X1 U803 ( .A(n711), .B(KEYINPUT100), .ZN(n713) );
  NAND2_X1 U804 ( .A1(n713), .A2(n516), .ZN(n714) );
  NOR2_X1 U805 ( .A1(n715), .A2(n714), .ZN(n719) );
  NOR2_X1 U806 ( .A1(n1002), .A2(n716), .ZN(n717) );
  XNOR2_X1 U807 ( .A(n717), .B(KEYINPUT28), .ZN(n718) );
  NOR2_X1 U808 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U809 ( .A(n720), .B(KEYINPUT29), .ZN(n723) );
  OR2_X1 U810 ( .A1(G301), .A2(n721), .ZN(n722) );
  NAND2_X1 U811 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U812 ( .A1(n725), .A2(n724), .ZN(n735) );
  NAND2_X1 U813 ( .A1(n735), .A2(G286), .ZN(n726) );
  XNOR2_X1 U814 ( .A(n726), .B(KEYINPUT102), .ZN(n732) );
  NAND2_X1 U815 ( .A1(G8), .A2(n727), .ZN(n766) );
  NOR2_X1 U816 ( .A1(G1971), .A2(n766), .ZN(n729) );
  NOR2_X1 U817 ( .A1(G2090), .A2(n727), .ZN(n728) );
  NOR2_X1 U818 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U819 ( .A1(n730), .A2(G303), .ZN(n731) );
  NAND2_X1 U820 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U821 ( .A1(n733), .A2(G8), .ZN(n734) );
  INV_X1 U822 ( .A(n735), .ZN(n741) );
  NAND2_X1 U823 ( .A1(G8), .A2(n736), .ZN(n737) );
  XNOR2_X1 U824 ( .A(n737), .B(KEYINPUT96), .ZN(n739) );
  NAND2_X1 U825 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U826 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U827 ( .A1(n517), .A2(n742), .ZN(n747) );
  NAND2_X1 U828 ( .A1(G8), .A2(G166), .ZN(n743) );
  NOR2_X1 U829 ( .A1(G2090), .A2(n743), .ZN(n744) );
  NOR2_X1 U830 ( .A1(n747), .A2(n744), .ZN(n745) );
  XNOR2_X1 U831 ( .A(n745), .B(KEYINPUT103), .ZN(n746) );
  NAND2_X1 U832 ( .A1(n746), .A2(n766), .ZN(n762) );
  INV_X1 U833 ( .A(n747), .ZN(n751) );
  NOR2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n754) );
  NOR2_X1 U835 ( .A1(G1971), .A2(G303), .ZN(n748) );
  NOR2_X1 U836 ( .A1(n754), .A2(n748), .ZN(n1007) );
  INV_X1 U837 ( .A(KEYINPUT33), .ZN(n749) );
  AND2_X1 U838 ( .A1(n1007), .A2(n749), .ZN(n750) );
  NAND2_X1 U839 ( .A1(n751), .A2(n750), .ZN(n760) );
  XOR2_X1 U840 ( .A(G1981), .B(G305), .Z(n989) );
  INV_X1 U841 ( .A(n766), .ZN(n752) );
  NAND2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n1006) );
  AND2_X1 U843 ( .A1(n752), .A2(n1006), .ZN(n753) );
  NOR2_X1 U844 ( .A1(KEYINPUT33), .A2(n753), .ZN(n757) );
  NAND2_X1 U845 ( .A1(n754), .A2(KEYINPUT33), .ZN(n755) );
  NOR2_X1 U846 ( .A1(n755), .A2(n766), .ZN(n756) );
  NOR2_X1 U847 ( .A1(n757), .A2(n756), .ZN(n758) );
  AND2_X1 U848 ( .A1(n989), .A2(n758), .ZN(n759) );
  NAND2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U850 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U851 ( .A(n763), .B(KEYINPUT104), .ZN(n768) );
  NOR2_X1 U852 ( .A1(G1981), .A2(G305), .ZN(n764) );
  XOR2_X1 U853 ( .A(n764), .B(KEYINPUT24), .Z(n765) );
  NOR2_X1 U854 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n803) );
  INV_X1 U856 ( .A(n769), .ZN(n771) );
  NOR2_X1 U857 ( .A1(n771), .A2(n770), .ZN(n818) );
  XNOR2_X1 U858 ( .A(KEYINPUT37), .B(G2067), .ZN(n816) );
  NAND2_X1 U859 ( .A1(n877), .A2(G104), .ZN(n773) );
  NAND2_X1 U860 ( .A1(G140), .A2(n875), .ZN(n772) );
  NAND2_X1 U861 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U862 ( .A(KEYINPUT34), .B(n774), .ZN(n781) );
  NAND2_X1 U863 ( .A1(n871), .A2(G116), .ZN(n775) );
  XNOR2_X1 U864 ( .A(KEYINPUT91), .B(n775), .ZN(n778) );
  NAND2_X1 U865 ( .A1(n872), .A2(G128), .ZN(n776) );
  XOR2_X1 U866 ( .A(KEYINPUT90), .B(n776), .Z(n777) );
  NOR2_X1 U867 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U868 ( .A(n779), .B(KEYINPUT35), .ZN(n780) );
  NOR2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U870 ( .A(KEYINPUT36), .B(n782), .ZN(n892) );
  NOR2_X1 U871 ( .A1(n816), .A2(n892), .ZN(n938) );
  NAND2_X1 U872 ( .A1(n818), .A2(n938), .ZN(n814) );
  NAND2_X1 U873 ( .A1(n871), .A2(G107), .ZN(n784) );
  NAND2_X1 U874 ( .A1(G131), .A2(n875), .ZN(n783) );
  NAND2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n877), .A2(G95), .ZN(n785) );
  XOR2_X1 U877 ( .A(KEYINPUT92), .B(n785), .Z(n786) );
  NOR2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n789) );
  NAND2_X1 U879 ( .A1(n872), .A2(G119), .ZN(n788) );
  NAND2_X1 U880 ( .A1(n789), .A2(n788), .ZN(n889) );
  NAND2_X1 U881 ( .A1(G1991), .A2(n889), .ZN(n800) );
  NAND2_X1 U882 ( .A1(n877), .A2(G105), .ZN(n790) );
  XNOR2_X1 U883 ( .A(n790), .B(KEYINPUT38), .ZN(n792) );
  NAND2_X1 U884 ( .A1(G117), .A2(n871), .ZN(n791) );
  NAND2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n795) );
  NAND2_X1 U886 ( .A1(G129), .A2(n872), .ZN(n793) );
  XNOR2_X1 U887 ( .A(KEYINPUT93), .B(n793), .ZN(n794) );
  NOR2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U889 ( .A(n796), .B(KEYINPUT94), .ZN(n798) );
  NAND2_X1 U890 ( .A1(G141), .A2(n875), .ZN(n797) );
  NAND2_X1 U891 ( .A1(n798), .A2(n797), .ZN(n866) );
  NAND2_X1 U892 ( .A1(G1996), .A2(n866), .ZN(n799) );
  NAND2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n934) );
  NAND2_X1 U894 ( .A1(n818), .A2(n934), .ZN(n801) );
  XOR2_X1 U895 ( .A(KEYINPUT95), .B(n801), .Z(n807) );
  NAND2_X1 U896 ( .A1(n814), .A2(n807), .ZN(n802) );
  NOR2_X1 U897 ( .A1(n803), .A2(n802), .ZN(n806) );
  XOR2_X1 U898 ( .A(G1986), .B(KEYINPUT89), .Z(n804) );
  XNOR2_X1 U899 ( .A(G290), .B(n804), .ZN(n994) );
  NAND2_X1 U900 ( .A1(n994), .A2(n818), .ZN(n805) );
  NAND2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n821) );
  NOR2_X1 U902 ( .A1(G1996), .A2(n866), .ZN(n924) );
  INV_X1 U903 ( .A(n807), .ZN(n811) );
  NOR2_X1 U904 ( .A1(G1991), .A2(n889), .ZN(n808) );
  XOR2_X1 U905 ( .A(KEYINPUT105), .B(n808), .Z(n930) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n809) );
  NOR2_X1 U907 ( .A1(n930), .A2(n809), .ZN(n810) );
  NOR2_X1 U908 ( .A1(n811), .A2(n810), .ZN(n812) );
  NOR2_X1 U909 ( .A1(n924), .A2(n812), .ZN(n813) );
  XNOR2_X1 U910 ( .A(n813), .B(KEYINPUT39), .ZN(n815) );
  NAND2_X1 U911 ( .A1(n815), .A2(n814), .ZN(n817) );
  NAND2_X1 U912 ( .A1(n816), .A2(n892), .ZN(n939) );
  NAND2_X1 U913 ( .A1(n817), .A2(n939), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U915 ( .A1(n821), .A2(n820), .ZN(n822) );
  XNOR2_X1 U916 ( .A(KEYINPUT40), .B(n822), .ZN(G329) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n918), .ZN(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n823) );
  NAND2_X1 U919 ( .A1(G661), .A2(n823), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U921 ( .A1(n825), .A2(n824), .ZN(G188) );
  INV_X1 U923 ( .A(G96), .ZN(G221) );
  NOR2_X1 U924 ( .A1(n827), .A2(n826), .ZN(n828) );
  XOR2_X1 U925 ( .A(n828), .B(KEYINPUT106), .Z(G261) );
  INV_X1 U926 ( .A(G261), .ZN(G325) );
  INV_X1 U927 ( .A(n829), .ZN(G319) );
  XNOR2_X1 U928 ( .A(G2090), .B(G2084), .ZN(n830) );
  XNOR2_X1 U929 ( .A(n830), .B(KEYINPUT107), .ZN(n840) );
  XOR2_X1 U930 ( .A(KEYINPUT42), .B(G2678), .Z(n832) );
  XNOR2_X1 U931 ( .A(KEYINPUT108), .B(G2096), .ZN(n831) );
  XNOR2_X1 U932 ( .A(n832), .B(n831), .ZN(n836) );
  XOR2_X1 U933 ( .A(G2100), .B(G2072), .Z(n834) );
  XNOR2_X1 U934 ( .A(G2067), .B(G2078), .ZN(n833) );
  XNOR2_X1 U935 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U936 ( .A(n836), .B(n835), .Z(n838) );
  XNOR2_X1 U937 ( .A(KEYINPUT43), .B(KEYINPUT109), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(G227) );
  XOR2_X1 U940 ( .A(G1971), .B(G1961), .Z(n842) );
  XNOR2_X1 U941 ( .A(G1986), .B(G1966), .ZN(n841) );
  XNOR2_X1 U942 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U943 ( .A(n843), .B(G2474), .Z(n845) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1991), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U946 ( .A(KEYINPUT41), .B(G1976), .Z(n847) );
  XOR2_X1 U947 ( .A(G1981), .B(n1003), .Z(n846) );
  XNOR2_X1 U948 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(G229) );
  NAND2_X1 U950 ( .A1(G124), .A2(n872), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n850), .B(KEYINPUT44), .ZN(n852) );
  NAND2_X1 U952 ( .A1(n871), .A2(G112), .ZN(n851) );
  NAND2_X1 U953 ( .A1(n852), .A2(n851), .ZN(n856) );
  NAND2_X1 U954 ( .A1(n877), .A2(G100), .ZN(n854) );
  NAND2_X1 U955 ( .A1(G136), .A2(n875), .ZN(n853) );
  NAND2_X1 U956 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U957 ( .A1(n856), .A2(n855), .ZN(G162) );
  NAND2_X1 U958 ( .A1(n877), .A2(G103), .ZN(n858) );
  NAND2_X1 U959 ( .A1(G139), .A2(n875), .ZN(n857) );
  NAND2_X1 U960 ( .A1(n858), .A2(n857), .ZN(n865) );
  XNOR2_X1 U961 ( .A(KEYINPUT114), .B(KEYINPUT47), .ZN(n863) );
  NAND2_X1 U962 ( .A1(n871), .A2(G115), .ZN(n861) );
  NAND2_X1 U963 ( .A1(n872), .A2(G127), .ZN(n859) );
  XOR2_X1 U964 ( .A(KEYINPUT113), .B(n859), .Z(n860) );
  NAND2_X1 U965 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U966 ( .A(n863), .B(n862), .Z(n864) );
  NOR2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n919) );
  XNOR2_X1 U968 ( .A(n919), .B(n866), .ZN(n867) );
  XNOR2_X1 U969 ( .A(n867), .B(n927), .ZN(n888) );
  XOR2_X1 U970 ( .A(KEYINPUT115), .B(KEYINPUT48), .Z(n869) );
  XNOR2_X1 U971 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n868) );
  XNOR2_X1 U972 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U973 ( .A(n870), .B(KEYINPUT116), .Z(n886) );
  NAND2_X1 U974 ( .A1(G118), .A2(n871), .ZN(n874) );
  NAND2_X1 U975 ( .A1(G130), .A2(n872), .ZN(n873) );
  NAND2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n883) );
  NAND2_X1 U977 ( .A1(G142), .A2(n875), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n876), .B(KEYINPUT110), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G106), .A2(n877), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U981 ( .A(KEYINPUT111), .B(n880), .ZN(n881) );
  XNOR2_X1 U982 ( .A(KEYINPUT45), .B(n881), .ZN(n882) );
  NOR2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U984 ( .A(G160), .B(n884), .ZN(n885) );
  XNOR2_X1 U985 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U986 ( .A(n888), .B(n887), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n889), .B(G162), .ZN(n890) );
  XNOR2_X1 U988 ( .A(n891), .B(n890), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n892), .B(G164), .ZN(n893) );
  XNOR2_X1 U990 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U991 ( .A1(G37), .A2(n895), .ZN(G395) );
  XOR2_X1 U992 ( .A(n896), .B(G286), .Z(n899) );
  XOR2_X1 U993 ( .A(G301), .B(n897), .Z(n898) );
  XNOR2_X1 U994 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U995 ( .A(n995), .B(n900), .Z(n901) );
  NOR2_X1 U996 ( .A1(G37), .A2(n901), .ZN(G397) );
  XOR2_X1 U997 ( .A(G2451), .B(G2430), .Z(n903) );
  XNOR2_X1 U998 ( .A(G2438), .B(G2443), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n909) );
  XOR2_X1 U1000 ( .A(G2435), .B(G2454), .Z(n905) );
  XNOR2_X1 U1001 ( .A(G1348), .B(G1341), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(n907) );
  XOR2_X1 U1003 ( .A(G2446), .B(G2427), .Z(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1005 ( .A(n909), .B(n908), .Z(n910) );
  NAND2_X1 U1006 ( .A1(G14), .A2(n910), .ZN(n917) );
  NAND2_X1 U1007 ( .A1(G319), .A2(n917), .ZN(n914) );
  NOR2_X1 U1008 ( .A1(G227), .A2(G229), .ZN(n911) );
  XOR2_X1 U1009 ( .A(KEYINPUT49), .B(n911), .Z(n912) );
  XNOR2_X1 U1010 ( .A(n912), .B(KEYINPUT117), .ZN(n913) );
  NOR2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(n916) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G69), .ZN(G235) );
  INV_X1 U1016 ( .A(n917), .ZN(G401) );
  INV_X1 U1017 ( .A(n918), .ZN(G223) );
  XOR2_X1 U1018 ( .A(G2072), .B(n919), .Z(n921) );
  XOR2_X1 U1019 ( .A(G164), .B(G2078), .Z(n920) );
  NOR2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1021 ( .A(KEYINPUT50), .B(n922), .ZN(n936) );
  XOR2_X1 U1022 ( .A(G2090), .B(G162), .Z(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1024 ( .A(KEYINPUT51), .B(n925), .Z(n932) );
  XNOR2_X1 U1025 ( .A(G160), .B(G2084), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(n926), .B(KEYINPUT118), .ZN(n928) );
  NAND2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  NOR2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1031 ( .A1(n936), .A2(n935), .ZN(n937) );
  NOR2_X1 U1032 ( .A1(n938), .A2(n937), .ZN(n940) );
  NAND2_X1 U1033 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1034 ( .A(KEYINPUT52), .B(n941), .ZN(n942) );
  NAND2_X1 U1035 ( .A1(n942), .A2(G29), .ZN(n1022) );
  XOR2_X1 U1036 ( .A(G16), .B(KEYINPUT123), .Z(n967) );
  XNOR2_X1 U1037 ( .A(G1966), .B(G21), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(G5), .B(G1961), .ZN(n943) );
  NOR2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n963) );
  XOR2_X1 U1040 ( .A(G20), .B(G1956), .Z(n948) );
  XNOR2_X1 U1041 ( .A(G1981), .B(G6), .ZN(n946) );
  XNOR2_X1 U1042 ( .A(G1341), .B(G19), .ZN(n945) );
  NOR2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n951) );
  XOR2_X1 U1045 ( .A(KEYINPUT59), .B(G1348), .Z(n949) );
  XNOR2_X1 U1046 ( .A(G4), .B(n949), .ZN(n950) );
  NOR2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1048 ( .A(KEYINPUT60), .B(n952), .Z(n961) );
  XOR2_X1 U1049 ( .A(G1976), .B(G23), .Z(n955) );
  XOR2_X1 U1050 ( .A(G22), .B(KEYINPUT124), .Z(n953) );
  XNOR2_X1 U1051 ( .A(n953), .B(G1971), .ZN(n954) );
  NAND2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n958) );
  XOR2_X1 U1053 ( .A(KEYINPUT125), .B(G1986), .Z(n956) );
  XNOR2_X1 U1054 ( .A(G24), .B(n956), .ZN(n957) );
  NOR2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1056 ( .A(KEYINPUT58), .B(n959), .Z(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(n964), .B(KEYINPUT61), .ZN(n965) );
  XNOR2_X1 U1060 ( .A(n965), .B(KEYINPUT126), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1062 ( .A(KEYINPUT127), .B(n968), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n969), .A2(G11), .ZN(n1020) );
  XOR2_X1 U1064 ( .A(G1991), .B(G25), .Z(n970) );
  NAND2_X1 U1065 ( .A1(n970), .A2(G28), .ZN(n979) );
  XNOR2_X1 U1066 ( .A(G1996), .B(G32), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(G33), .B(G2072), .ZN(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(G2067), .B(G26), .ZN(n975) );
  XNOR2_X1 U1070 ( .A(G27), .B(n973), .ZN(n974) );
  NOR2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1074 ( .A(KEYINPUT53), .B(n980), .Z(n983) );
  XOR2_X1 U1075 ( .A(G34), .B(KEYINPUT54), .Z(n981) );
  XNOR2_X1 U1076 ( .A(G2084), .B(n981), .ZN(n982) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(G35), .B(G2090), .ZN(n984) );
  NOR2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1080 ( .A(KEYINPUT119), .B(n986), .Z(n987) );
  NOR2_X1 U1081 ( .A1(G29), .A2(n987), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(n988), .B(KEYINPUT55), .ZN(n1018) );
  XNOR2_X1 U1083 ( .A(KEYINPUT56), .B(G16), .ZN(n1016) );
  XNOR2_X1 U1084 ( .A(G1966), .B(G168), .ZN(n990) );
  NAND2_X1 U1085 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1086 ( .A(n991), .B(KEYINPUT57), .ZN(n992) );
  XOR2_X1 U1087 ( .A(KEYINPUT120), .B(n992), .Z(n993) );
  NOR2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n1014) );
  XNOR2_X1 U1089 ( .A(n995), .B(G1341), .ZN(n996) );
  XNOR2_X1 U1090 ( .A(n996), .B(KEYINPUT122), .ZN(n1001) );
  XOR2_X1 U1091 ( .A(G171), .B(G1961), .Z(n999) );
  XOR2_X1 U1092 ( .A(n997), .B(G1348), .Z(n998) );
  NOR2_X1 U1093 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1012) );
  XOR2_X1 U1095 ( .A(n1003), .B(n1002), .Z(n1005) );
  NAND2_X1 U1096 ( .A1(G1971), .A2(G303), .ZN(n1004) );
  NAND2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(KEYINPUT121), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(KEYINPUT62), .B(n1023), .ZN(G150) );
  INV_X1 U1108 ( .A(G150), .ZN(G311) );
endmodule

