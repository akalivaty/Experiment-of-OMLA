//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1264, new_n1265, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT65), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G87), .A2(G250), .ZN(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT66), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT64), .B(G77), .ZN(new_n215));
  AOI22_X1  g0015(.A1(new_n213), .A2(new_n214), .B1(G244), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(KEYINPUT66), .B1(new_n208), .B2(new_n212), .ZN(new_n217));
  AND2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  INV_X1    g0019(.A(G116), .ZN(new_n220));
  INV_X1    g0020(.A(G270), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G68), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n206), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT1), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n206), .A2(G13), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT0), .Z(new_n230));
  OAI21_X1  g0030(.A(G50), .B1(G58), .B2(G68), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR3_X1   g0033(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NOR3_X1   g0034(.A1(new_n227), .A2(new_n230), .A3(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XOR2_X1   g0044(.A(G50), .B(G58), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT67), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  AND2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G1698), .ZN(new_n255));
  OAI21_X1  g0055(.A(KEYINPUT69), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT3), .B(G33), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT69), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(new_n258), .A3(G1698), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n256), .A2(new_n259), .A3(G223), .ZN(new_n260));
  OR2_X1    g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  AOI21_X1  g0062(.A(G1698), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G222), .ZN(new_n264));
  INV_X1    g0064(.A(new_n215), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n260), .B(new_n264), .C1(new_n265), .C2(new_n257), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  OAI211_X1 g0068(.A(G1), .B(G13), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AND2_X1   g0070(.A1(new_n266), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G1), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n272), .B1(G41), .B2(G45), .ZN(new_n273));
  INV_X1    g0073(.A(G274), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AND2_X1   g0075(.A1(new_n269), .A2(new_n273), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n275), .B1(new_n276), .B2(G226), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n277), .B(KEYINPUT68), .ZN(new_n278));
  OR2_X1    g0078(.A1(new_n271), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G169), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n203), .A2(G20), .ZN(new_n282));
  INV_X1    g0082(.A(G150), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n232), .A2(new_n267), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n232), .A2(G33), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  OAI221_X1 g0086(.A(new_n282), .B1(new_n283), .B2(new_n284), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(new_n233), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n272), .A2(G13), .A3(G20), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n202), .ZN(new_n293));
  INV_X1    g0093(.A(new_n289), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n272), .A2(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n290), .B(new_n293), .C1(new_n202), .C2(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n271), .A2(new_n278), .ZN(new_n298));
  INV_X1    g0098(.A(G179), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n281), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT70), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT70), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g0106(.A(KEYINPUT7), .B1(new_n254), .B2(new_n232), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n232), .A4(new_n262), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(G68), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT75), .ZN(new_n311));
  NOR2_X1   g0111(.A1(G20), .A2(G33), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n311), .B1(new_n312), .B2(G159), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n312), .A2(new_n311), .A3(G159), .ZN(new_n315));
  XNOR2_X1  g0115(.A(G58), .B(G68), .ZN(new_n316));
  AOI22_X1  g0116(.A1(new_n314), .A2(new_n315), .B1(new_n316), .B2(G20), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n310), .A2(KEYINPUT16), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(G20), .ZN(new_n319));
  INV_X1    g0119(.A(new_n315), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(new_n313), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT76), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n308), .A2(new_n322), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n254), .A2(KEYINPUT76), .A3(KEYINPUT7), .A4(new_n232), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT7), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n325), .B1(new_n257), .B2(G20), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n323), .A2(new_n324), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n321), .B1(new_n327), .B2(G68), .ZN(new_n328));
  OAI211_X1 g0128(.A(new_n289), .B(new_n318), .C1(new_n328), .C2(KEYINPUT16), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n219), .A2(G1698), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n330), .B1(G223), .B2(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G87), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n270), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n275), .B1(new_n276), .B2(G232), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n334), .A2(new_n335), .A3(G190), .ZN(new_n336));
  INV_X1    g0136(.A(new_n286), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n296), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(new_n292), .B2(new_n337), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n269), .B1(new_n331), .B2(new_n332), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n273), .A2(new_n274), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n269), .A2(new_n273), .ZN(new_n342));
  INV_X1    g0142(.A(G232), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(G200), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n329), .A2(new_n336), .A3(new_n339), .A4(new_n345), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n346), .B(KEYINPUT17), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT18), .ZN(new_n348));
  AND2_X1   g0148(.A1(new_n329), .A2(new_n339), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n280), .B1(new_n334), .B2(new_n335), .ZN(new_n350));
  NOR3_X1   g0150(.A1(new_n340), .A2(new_n344), .A3(new_n299), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n348), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n329), .A2(new_n339), .ZN(new_n354));
  INV_X1    g0154(.A(new_n352), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(new_n355), .A3(KEYINPUT18), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n306), .A2(new_n347), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n298), .A2(G190), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n297), .B(KEYINPUT9), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT72), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n361), .B1(new_n279), .B2(G200), .ZN(new_n362));
  INV_X1    g0162(.A(G200), .ZN(new_n363));
  NOR3_X1   g0163(.A1(new_n298), .A2(KEYINPUT72), .A3(new_n363), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n359), .B(new_n360), .C1(new_n362), .C2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT10), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n365), .B(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT74), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G33), .A2(G97), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n257), .B1(G232), .B2(new_n255), .ZN(new_n370));
  NOR2_X1   g0170(.A1(G226), .A2(G1698), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n270), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n276), .A2(G238), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n341), .A3(new_n374), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n375), .A2(KEYINPUT13), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n375), .A2(KEYINPUT13), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n368), .B(KEYINPUT14), .C1(new_n378), .C2(new_n280), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(G179), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n368), .A2(KEYINPUT14), .ZN(new_n381));
  OAI211_X1 g0181(.A(G169), .B(new_n381), .C1(new_n376), .C2(new_n377), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n296), .A2(new_n223), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n384), .B(KEYINPUT73), .ZN(new_n385));
  OAI22_X1  g0185(.A1(new_n284), .A2(new_n202), .B1(new_n232), .B2(G68), .ZN(new_n386));
  INV_X1    g0186(.A(G77), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n285), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n289), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g0189(.A(new_n389), .B(KEYINPUT11), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n292), .A2(new_n223), .ZN(new_n391));
  XNOR2_X1  g0191(.A(new_n391), .B(KEYINPUT12), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n385), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n383), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G244), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n342), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n256), .A2(new_n259), .A3(G238), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n263), .A2(G232), .B1(new_n254), .B2(G107), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI211_X1 g0199(.A(new_n396), .B(new_n275), .C1(new_n399), .C2(new_n270), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n299), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n215), .A2(new_n291), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n337), .A2(new_n312), .B1(new_n215), .B2(G20), .ZN(new_n403));
  XOR2_X1   g0203(.A(KEYINPUT15), .B(G87), .Z(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n403), .B1(new_n285), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n402), .B1(new_n406), .B2(new_n289), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n387), .B2(new_n296), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n401), .B(new_n408), .C1(G169), .C2(new_n400), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n378), .A2(G190), .ZN(new_n410));
  INV_X1    g0210(.A(new_n393), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n410), .B(new_n411), .C1(new_n363), .C2(new_n378), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n394), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n275), .B1(new_n399), .B2(new_n270), .ZN(new_n414));
  INV_X1    g0214(.A(new_n396), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n363), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(KEYINPUT71), .B1(new_n416), .B2(new_n408), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n400), .A2(G190), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n296), .A2(new_n387), .ZN(new_n419));
  AOI211_X1 g0219(.A(new_n419), .B(new_n402), .C1(new_n406), .C2(new_n289), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT71), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n420), .B(new_n421), .C1(new_n400), .C2(new_n363), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n417), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NOR4_X1   g0224(.A1(new_n358), .A2(new_n367), .A3(new_n413), .A4(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT83), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n232), .B1(new_n210), .B2(G33), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G283), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT77), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(KEYINPUT77), .A2(G33), .A3(G283), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n427), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n289), .B1(new_n232), .B2(G116), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n426), .B(KEYINPUT20), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n430), .A2(new_n431), .ZN(new_n435));
  INV_X1    g0235(.A(new_n427), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n426), .A2(KEYINPUT20), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n426), .A2(KEYINPUT20), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n288), .A2(new_n233), .B1(G20), .B2(new_n220), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n437), .A2(new_n438), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n292), .A2(new_n220), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n272), .A2(G33), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n294), .A2(G116), .A3(new_n291), .A4(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n434), .A2(new_n441), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n445), .A2(G169), .ZN(new_n446));
  INV_X1    g0246(.A(G45), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(G1), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n268), .A2(KEYINPUT5), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT5), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G41), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n448), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n269), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT81), .B1(new_n453), .B2(new_n221), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT81), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n452), .A2(new_n455), .A3(G270), .A4(new_n269), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n452), .A2(new_n274), .ZN(new_n458));
  OAI211_X1 g0258(.A(G257), .B(new_n255), .C1(new_n252), .C2(new_n253), .ZN(new_n459));
  OAI211_X1 g0259(.A(G264), .B(G1698), .C1(new_n252), .C2(new_n253), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n261), .A2(G303), .A3(new_n262), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT82), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n462), .A2(new_n463), .A3(new_n270), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n463), .B1(new_n462), .B2(new_n270), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n457), .B(new_n458), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n446), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT21), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n466), .A2(G200), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n462), .A2(new_n270), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT82), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n462), .A2(new_n463), .A3(new_n270), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n474), .A2(G190), .A3(new_n458), .A4(new_n457), .ZN(new_n475));
  INV_X1    g0275(.A(new_n445), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n470), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n466), .A2(new_n299), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n445), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n446), .A2(KEYINPUT21), .A3(new_n466), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n469), .A2(new_n477), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT84), .ZN(new_n482));
  AND3_X1   g0282(.A1(new_n446), .A2(KEYINPUT21), .A3(new_n466), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT21), .B1(new_n446), .B2(new_n466), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT84), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n485), .A2(new_n486), .A3(new_n479), .A4(new_n477), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n294), .A2(new_n291), .A3(new_n443), .ZN(new_n489));
  INV_X1    g0289(.A(G107), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n292), .A2(new_n490), .ZN(new_n493));
  XNOR2_X1  g0293(.A(new_n493), .B(KEYINPUT25), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT23), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT85), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT85), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT23), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n497), .A2(new_n499), .B1(G20), .B2(new_n490), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n496), .A2(KEYINPUT85), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n490), .A2(G20), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n232), .B(G87), .C1(new_n252), .C2(new_n253), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT22), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n285), .A2(new_n220), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n257), .A2(KEYINPUT22), .A3(new_n232), .A4(G87), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n504), .A2(new_n507), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT24), .ZN(new_n512));
  INV_X1    g0312(.A(new_n505), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n508), .B1(new_n513), .B2(KEYINPUT22), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT24), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n514), .A2(new_n515), .A3(new_n507), .A4(new_n504), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n492), .B(new_n495), .C1(new_n517), .C2(new_n294), .ZN(new_n518));
  OAI211_X1 g0318(.A(G250), .B(new_n255), .C1(new_n252), .C2(new_n253), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT86), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT86), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n257), .A2(new_n521), .A3(G250), .A4(new_n255), .ZN(new_n522));
  NAND2_X1  g0322(.A1(G33), .A2(G294), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n257), .A2(G257), .A3(G1698), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n520), .A2(new_n522), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n270), .ZN(new_n526));
  INV_X1    g0326(.A(new_n453), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(G264), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n458), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n280), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n525), .A2(new_n270), .B1(G264), .B2(new_n527), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(new_n299), .A3(new_n458), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n518), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(G190), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n526), .A2(new_n534), .A3(new_n458), .A4(new_n528), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT87), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n529), .A2(new_n363), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT87), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n531), .A2(new_n538), .A3(new_n534), .A4(new_n458), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n294), .B1(new_n512), .B2(new_n516), .ZN(new_n541));
  NOR3_X1   g0341(.A1(new_n541), .A2(new_n491), .A3(new_n494), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n533), .A2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(G244), .B(new_n255), .C1(new_n252), .C2(new_n253), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT4), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n257), .A2(KEYINPUT4), .A3(G244), .A4(new_n255), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n257), .A2(G250), .A3(G1698), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n435), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n270), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n453), .A2(new_n211), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n552), .A2(new_n458), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT78), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n547), .A2(new_n548), .A3(new_n435), .A4(new_n550), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n553), .B1(new_n558), .B2(new_n270), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n559), .A2(KEYINPUT78), .A3(new_n458), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n557), .A2(G200), .A3(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n291), .A2(G97), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n489), .A2(new_n210), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n327), .A2(G107), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n490), .A2(KEYINPUT6), .A3(G97), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n210), .A2(new_n490), .ZN(new_n566));
  NOR2_X1   g0366(.A1(G97), .A2(G107), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n565), .B1(new_n568), .B2(KEYINPUT6), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n569), .A2(G20), .B1(G77), .B2(new_n312), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n564), .A2(new_n570), .ZN(new_n571));
  AOI211_X1 g0371(.A(new_n562), .B(new_n563), .C1(new_n571), .C2(new_n289), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n559), .A2(G190), .A3(new_n458), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n561), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n571), .A2(new_n289), .ZN(new_n575));
  INV_X1    g0375(.A(new_n563), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n555), .A2(new_n299), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n280), .B1(new_n559), .B2(new_n458), .ZN(new_n579));
  OAI22_X1  g0379(.A1(new_n577), .A2(new_n562), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT19), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n582), .A2(new_n232), .A3(G33), .A4(G97), .ZN(new_n583));
  INV_X1    g0383(.A(G87), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n567), .A2(new_n584), .B1(new_n369), .B2(new_n232), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n583), .B1(new_n585), .B2(new_n582), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n232), .B(G68), .C1(new_n252), .C2(new_n253), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(KEYINPUT79), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT79), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n257), .A2(new_n589), .A3(new_n232), .A4(G68), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n586), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n289), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n405), .A2(new_n292), .ZN(new_n593));
  INV_X1    g0393(.A(new_n489), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n404), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT80), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n269), .B(G250), .C1(G1), .C2(new_n447), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n448), .A2(G274), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n224), .A2(new_n255), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n395), .A2(G1698), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n601), .B(new_n602), .C1(new_n252), .C2(new_n253), .ZN(new_n603));
  NAND2_X1  g0403(.A1(G33), .A2(G116), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n600), .B1(new_n270), .B2(new_n605), .ZN(new_n606));
  OR2_X1    g0406(.A1(new_n606), .A2(G169), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n299), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT80), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n592), .A2(new_n609), .A3(new_n593), .A4(new_n595), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n597), .A2(new_n607), .A3(new_n608), .A4(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n594), .A2(G87), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n592), .A2(new_n593), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n606), .A2(G190), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n613), .B(new_n614), .C1(new_n363), .C2(new_n606), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n544), .A2(new_n581), .A3(new_n616), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n425), .A2(new_n488), .A3(new_n617), .ZN(G372));
  AND2_X1   g0418(.A1(new_n574), .A2(new_n580), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT89), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT88), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n605), .B2(new_n270), .ZN(new_n622));
  AOI211_X1 g0422(.A(KEYINPUT88), .B(new_n269), .C1(new_n603), .C2(new_n604), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n599), .B(new_n598), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n280), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n597), .A2(new_n625), .A3(new_n608), .A4(new_n610), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n624), .A2(G200), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n627), .A2(new_n613), .A3(new_n614), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n619), .A2(new_n620), .A3(new_n543), .A4(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n574), .A2(new_n543), .A3(new_n580), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n626), .A2(new_n628), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT89), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n466), .A2(new_n476), .A3(new_n299), .ZN(new_n634));
  NOR3_X1   g0434(.A1(new_n483), .A2(new_n484), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n533), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n630), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n578), .A2(new_n579), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(new_n572), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n629), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(KEYINPUT26), .B1(new_n616), .B2(new_n580), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n641), .A2(new_n626), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n637), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n425), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n306), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n367), .A2(KEYINPUT90), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n365), .B(KEYINPUT10), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT90), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n394), .A2(new_n409), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(new_n412), .A3(new_n347), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(new_n357), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n646), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n645), .A2(new_n655), .ZN(G369));
  AOI21_X1  g0456(.A(new_n486), .B1(new_n635), .B2(new_n477), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n481), .A2(KEYINPUT84), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT92), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(G13), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n660), .A2(G20), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n272), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT27), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n661), .A2(new_n664), .A3(new_n272), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n663), .A2(G213), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT91), .ZN(new_n667));
  INV_X1    g0467(.A(G343), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(new_n476), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT92), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n482), .A2(new_n487), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n659), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n469), .A2(new_n479), .A3(new_n480), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n671), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT93), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT93), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n675), .A2(new_n680), .A3(new_n677), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n544), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n542), .B2(new_n670), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n518), .A2(new_n530), .A3(new_n532), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(new_n669), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n682), .A2(G330), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n676), .A2(new_n670), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(new_n544), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n669), .B(KEYINPUT94), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n691), .B1(new_n685), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n689), .A2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n228), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n567), .A2(new_n584), .A3(new_n220), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n697), .A2(G1), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(new_n231), .B2(new_n697), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT28), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n466), .A2(new_n529), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n703), .A2(new_n299), .A3(new_n555), .A4(new_n624), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n531), .A2(new_n559), .A3(new_n458), .A4(new_n606), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n705), .B1(new_n707), .B2(new_n478), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n474), .A2(G179), .A3(new_n458), .A4(new_n457), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n709), .A2(new_n706), .A3(KEYINPUT30), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n704), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT95), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI211_X1 g0513(.A(new_n704), .B(KEYINPUT95), .C1(new_n708), .C2(new_n710), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n713), .A2(new_n669), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT31), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n617), .A2(new_n488), .A3(new_n692), .ZN(new_n718));
  INV_X1    g0518(.A(new_n692), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n711), .A2(KEYINPUT31), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G330), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n629), .A2(new_n543), .A3(new_n580), .A4(new_n574), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n685), .A2(new_n676), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT96), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n574), .A2(new_n543), .A3(new_n580), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT96), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n726), .A2(new_n636), .A3(new_n727), .A4(new_n629), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT26), .B1(new_n632), .B2(new_n580), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n640), .A2(new_n638), .A3(new_n611), .A4(new_n615), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n730), .A2(new_n626), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n725), .A2(new_n728), .A3(new_n729), .A4(new_n731), .ZN(new_n732));
  AND3_X1   g0532(.A1(new_n732), .A2(KEYINPUT29), .A3(new_n670), .ZN(new_n733));
  AOI21_X1  g0533(.A(KEYINPUT29), .B1(new_n644), .B2(new_n692), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n722), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n702), .B1(new_n736), .B2(G1), .ZN(G364));
  AND3_X1   g0537(.A1(new_n675), .A2(new_n680), .A3(new_n677), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n680), .B1(new_n675), .B2(new_n677), .ZN(new_n739));
  OAI21_X1  g0539(.A(G330), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(G330), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n679), .A2(new_n741), .A3(new_n681), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n661), .A2(G45), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n697), .A2(G1), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n740), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n745), .A2(KEYINPUT97), .ZN(new_n746));
  XNOR2_X1  g0546(.A(KEYINPUT98), .B(G169), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  INV_X1    g0548(.A(new_n233), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n232), .A2(G190), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n363), .A2(G179), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G107), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G179), .A2(G200), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n232), .B1(new_n756), .B2(G190), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n299), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(new_n751), .ZN(new_n759));
  OAI221_X1 g0559(.A(new_n755), .B1(new_n210), .B2(new_n757), .C1(new_n265), .C2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n299), .A2(new_n363), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n751), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n760), .B1(G68), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n232), .A2(new_n534), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(new_n752), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n584), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n765), .A2(new_n761), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n765), .A2(new_n758), .ZN(new_n770));
  INV_X1    g0570(.A(G58), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n769), .A2(new_n202), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT32), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n751), .A2(new_n756), .ZN(new_n774));
  INV_X1    g0574(.A(G159), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n774), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(KEYINPUT32), .A3(G159), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n772), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n764), .A2(new_n257), .A3(new_n768), .A4(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G303), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n254), .B1(new_n766), .B2(new_n781), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT100), .Z(new_n783));
  INV_X1    g0583(.A(G322), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n770), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(G283), .ZN(new_n786));
  INV_X1    g0586(.A(G329), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n753), .A2(new_n786), .B1(new_n774), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(KEYINPUT33), .B(G317), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n785), .B(new_n788), .C1(new_n763), .C2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n759), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G311), .ZN(new_n792));
  INV_X1    g0592(.A(new_n769), .ZN(new_n793));
  INV_X1    g0593(.A(new_n757), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n793), .A2(G326), .B1(new_n794), .B2(G294), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n783), .A2(new_n790), .A3(new_n792), .A4(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n750), .B1(new_n780), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n750), .ZN(new_n798));
  NOR2_X1   g0598(.A1(G13), .A2(G33), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(G20), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT99), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n695), .A2(new_n257), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(new_n246), .B2(G45), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(G45), .B2(new_n231), .ZN(new_n807));
  INV_X1    g0607(.A(G355), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n257), .A2(new_n228), .ZN(new_n809));
  OAI221_X1 g0609(.A(new_n807), .B1(G116), .B2(new_n228), .C1(new_n808), .C2(new_n809), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n744), .B(new_n797), .C1(new_n803), .C2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n801), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n682), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n745), .A2(KEYINPUT97), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n746), .A2(new_n813), .A3(new_n814), .ZN(G396));
  NAND2_X1  g0615(.A1(new_n408), .A2(new_n669), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n423), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(new_n409), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n409), .A2(new_n669), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(new_n644), .B2(new_n692), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n719), .B(new_n820), .C1(new_n637), .C2(new_n643), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n722), .ZN(new_n825));
  OAI211_X1 g0625(.A(G330), .B(new_n721), .C1(new_n822), .C2(new_n823), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n825), .A2(new_n744), .A3(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT103), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n753), .A2(new_n584), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n762), .A2(new_n786), .B1(new_n757), .B2(new_n210), .ZN(new_n830));
  INV_X1    g0630(.A(new_n770), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n829), .B(new_n830), .C1(G294), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n791), .A2(G116), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n793), .A2(G303), .B1(new_n777), .B2(G311), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n254), .B1(new_n766), .B2(new_n490), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT101), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n832), .A2(new_n833), .A3(new_n834), .A4(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(G143), .A2(new_n831), .B1(new_n791), .B2(G159), .ZN(new_n838));
  INV_X1    g0638(.A(G137), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n838), .B1(new_n839), .B2(new_n769), .C1(new_n283), .C2(new_n762), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT102), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT34), .ZN(new_n842));
  INV_X1    g0642(.A(G132), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n774), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n753), .A2(new_n223), .ZN(new_n845));
  INV_X1    g0645(.A(new_n766), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n844), .B(new_n845), .C1(G50), .C2(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n842), .A2(new_n257), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n757), .A2(new_n771), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n837), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n798), .A2(new_n799), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n850), .A2(new_n798), .B1(new_n387), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n800), .B2(new_n821), .ZN(new_n853));
  INV_X1    g0653(.A(new_n744), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  AND3_X1   g0655(.A1(new_n827), .A2(new_n828), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n828), .B1(new_n827), .B2(new_n855), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n856), .A2(new_n857), .ZN(G384));
  NAND4_X1  g0658(.A1(new_n349), .A2(KEYINPUT17), .A3(new_n336), .A4(new_n345), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT17), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n346), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(KEYINPUT18), .B1(new_n354), .B2(new_n355), .ZN(new_n862));
  AOI211_X1 g0662(.A(new_n348), .B(new_n352), .C1(new_n339), .C2(new_n329), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n859), .B(new_n861), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n349), .A2(new_n667), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n329), .A2(new_n339), .B1(new_n352), .B2(new_n667), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n867), .A2(new_n868), .A3(new_n346), .ZN(new_n869));
  INV_X1    g0669(.A(new_n346), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT37), .B1(new_n870), .B2(new_n866), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n864), .A2(new_n865), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT105), .B1(new_n872), .B2(KEYINPUT38), .ZN(new_n873));
  AOI21_X1  g0673(.A(KEYINPUT16), .B1(new_n310), .B2(new_n317), .ZN(new_n874));
  OAI21_X1  g0674(.A(KEYINPUT104), .B1(new_n874), .B2(new_n294), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT104), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n326), .A2(new_n308), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n321), .B1(new_n877), .B2(G68), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n876), .B(new_n289), .C1(new_n878), .C2(KEYINPUT16), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n875), .A2(new_n318), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n667), .B1(new_n880), .B2(new_n339), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n352), .B1(new_n880), .B2(new_n339), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n881), .A2(new_n882), .A3(new_n870), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n869), .B1(new_n883), .B2(new_n868), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n864), .A2(new_n881), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n884), .A2(KEYINPUT38), .A3(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT105), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT38), .ZN(new_n888));
  INV_X1    g0688(.A(new_n865), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n357), .B2(new_n347), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n869), .A2(new_n871), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n887), .B(new_n888), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n873), .A2(new_n886), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n669), .A4(new_n714), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n717), .A2(new_n718), .A3(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n394), .A2(new_n669), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n393), .A2(new_n669), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n383), .A2(new_n393), .B1(new_n412), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n896), .A2(new_n821), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(KEYINPUT40), .B1(new_n894), .B2(new_n901), .ZN(new_n902));
  AND3_X1   g0702(.A1(new_n896), .A2(new_n821), .A3(new_n900), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT38), .B1(new_n884), .B2(new_n885), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(KEYINPUT40), .B1(new_n905), .B2(new_n886), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n903), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n741), .B1(new_n902), .B2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n425), .A2(new_n896), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n908), .B1(G330), .B2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT106), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n911), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n903), .A2(new_n893), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n914), .A2(KEYINPUT40), .B1(new_n903), .B2(new_n906), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n425), .A2(new_n896), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n912), .B(new_n913), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n733), .A2(new_n734), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n425), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n655), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n917), .B(new_n920), .Z(new_n921));
  NAND2_X1  g0721(.A1(new_n905), .A2(new_n886), .ZN(new_n922));
  INV_X1    g0722(.A(new_n819), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n922), .B(new_n900), .C1(new_n823), .C2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n667), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n357), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n870), .A2(new_n866), .A3(KEYINPUT37), .ZN(new_n928));
  INV_X1    g0728(.A(new_n881), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n880), .A2(new_n339), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n355), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n929), .A2(new_n931), .A3(new_n346), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n928), .B1(new_n932), .B2(KEYINPUT37), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n929), .B1(new_n357), .B2(new_n347), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n933), .A2(new_n934), .A3(new_n888), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT39), .B1(new_n935), .B2(new_n904), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT39), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n873), .A2(new_n937), .A3(new_n892), .A4(new_n886), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n897), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n924), .B(new_n927), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n921), .B(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n272), .B2(new_n661), .ZN(new_n943));
  OAI211_X1 g0743(.A(G20), .B(new_n749), .C1(new_n569), .C2(KEYINPUT35), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n220), .B(new_n944), .C1(KEYINPUT35), .C2(new_n569), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n945), .B(KEYINPUT36), .Z(new_n946));
  INV_X1    g0746(.A(new_n231), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n771), .B2(new_n223), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n948), .A2(new_n265), .B1(G50), .B2(new_n223), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(G1), .A3(new_n660), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n943), .A2(new_n946), .A3(new_n950), .ZN(G367));
  AOI22_X1  g0751(.A1(G159), .A2(new_n763), .B1(new_n791), .B2(G50), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n794), .A2(G68), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n952), .B(new_n953), .C1(new_n283), .C2(new_n770), .ZN(new_n954));
  INV_X1    g0754(.A(G143), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n769), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n774), .A2(new_n839), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n257), .B1(new_n766), .B2(new_n771), .C1(new_n265), .C2(new_n753), .ZN(new_n958));
  NOR4_X1   g0758(.A1(new_n954), .A2(new_n956), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(G311), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n769), .A2(new_n960), .B1(new_n770), .B2(new_n781), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT111), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n962), .B1(G97), .B2(new_n754), .ZN(new_n963));
  INV_X1    g0763(.A(G317), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n963), .B1(new_n490), .B2(new_n757), .C1(new_n964), .C2(new_n774), .ZN(new_n965));
  INV_X1    g0765(.A(G294), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n762), .A2(new_n966), .B1(new_n759), .B2(new_n786), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n965), .A2(new_n257), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(KEYINPUT112), .B1(new_n766), .B2(new_n220), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT46), .Z(new_n970));
  AOI21_X1  g0770(.A(new_n959), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n971), .B(KEYINPUT47), .Z(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n798), .ZN(new_n973));
  OR2_X1    g0773(.A1(new_n670), .A2(new_n613), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n974), .A2(new_n626), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n629), .A2(new_n974), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n975), .A2(new_n976), .A3(new_n801), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n802), .B1(new_n228), .B2(new_n405), .C1(new_n242), .C2(new_n805), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n973), .A2(new_n977), .A3(new_n854), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n743), .A2(G1), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT109), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n691), .B1(new_n687), .B2(new_n690), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n740), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n982), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n984), .B(G330), .C1(new_n738), .C2(new_n739), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n981), .B1(new_n986), .B2(new_n736), .ZN(new_n987));
  AOI211_X1 g0787(.A(KEYINPUT109), .B(new_n735), .C1(new_n983), .C2(new_n985), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n692), .A2(new_n580), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT107), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n619), .B1(new_n572), .B2(new_n692), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n693), .ZN(new_n995));
  AOI21_X1  g0795(.A(KEYINPUT44), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT44), .ZN(new_n997));
  NOR3_X1   g0797(.A1(new_n993), .A2(new_n693), .A3(new_n997), .ZN(new_n998));
  AND3_X1   g0798(.A1(new_n993), .A2(KEYINPUT45), .A3(new_n693), .ZN(new_n999));
  AOI21_X1  g0799(.A(KEYINPUT45), .B1(new_n993), .B2(new_n693), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n996), .A2(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n689), .B(new_n1001), .ZN(new_n1002));
  AOI21_X1  g0802(.A(KEYINPUT110), .B1(new_n989), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n984), .B1(new_n682), .B2(G330), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n741), .B(new_n982), .C1(new_n679), .C2(new_n681), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n736), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(KEYINPUT109), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n735), .B1(new_n983), .B2(new_n985), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n981), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1007), .A2(new_n1002), .A3(new_n1009), .A4(KEYINPUT110), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n736), .B1(new_n1003), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n696), .B(KEYINPUT41), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n980), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n993), .A2(new_n691), .ZN(new_n1015));
  XOR2_X1   g0815(.A(KEYINPUT108), .B(KEYINPUT42), .Z(new_n1016));
  XNOR2_X1  g0816(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n580), .B1(new_n994), .B2(new_n533), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1018), .A2(new_n692), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n975), .A2(new_n976), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(new_n1017), .A2(new_n1019), .B1(KEYINPUT43), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1020), .A2(KEYINPUT43), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1021), .B(new_n1022), .Z(new_n1023));
  OR3_X1    g0823(.A1(new_n1023), .A2(new_n689), .A3(new_n994), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1023), .B1(new_n689), .B2(new_n994), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n979), .B1(new_n1014), .B2(new_n1026), .ZN(G387));
  XOR2_X1   g0827(.A(KEYINPUT113), .B(G150), .Z(new_n1028));
  NOR2_X1   g0828(.A1(new_n1028), .A2(new_n774), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G68), .A2(new_n791), .B1(new_n794), .B2(new_n404), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1030), .B1(new_n775), .B2(new_n769), .C1(new_n286), .C2(new_n762), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1029), .B(new_n1031), .C1(G50), .C2(new_n831), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n754), .A2(G97), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n846), .A2(new_n215), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1032), .A2(new_n257), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n770), .A2(new_n964), .B1(new_n759), .B2(new_n781), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT114), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1037), .B1(new_n960), .B2(new_n762), .C1(new_n784), .C2(new_n769), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT48), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n786), .B2(new_n757), .C1(new_n966), .C2(new_n766), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT49), .Z(new_n1041));
  AOI21_X1  g0841(.A(new_n257), .B1(new_n777), .B2(G326), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n220), .B2(new_n753), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1035), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT115), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g0846(.A(KEYINPUT115), .B(new_n1035), .C1(new_n1041), .C2(new_n1043), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1046), .A2(new_n798), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n687), .A2(new_n801), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n286), .A2(G50), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT50), .ZN(new_n1051));
  AOI21_X1  g0851(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1051), .A2(new_n699), .A3(new_n1052), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n804), .B(new_n1053), .C1(new_n239), .C2(new_n447), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1054), .B1(G107), .B2(new_n228), .C1(new_n699), .C2(new_n809), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n803), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1048), .A2(new_n854), .A3(new_n1049), .A4(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT116), .ZN(new_n1058));
  AND2_X1   g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g0859(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n980), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n983), .B2(new_n985), .ZN(new_n1062));
  NOR3_X1   g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n983), .A2(new_n735), .A3(new_n985), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1006), .A2(new_n696), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(KEYINPUT117), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT117), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1063), .A2(new_n1068), .A3(new_n1065), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1069), .ZN(G393));
  NAND2_X1  g0870(.A1(new_n1002), .A2(new_n980), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n994), .A2(new_n801), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n802), .B1(new_n210), .B2(new_n228), .C1(new_n250), .C2(new_n805), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n769), .A2(new_n283), .B1(new_n770), .B2(new_n775), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1074), .A2(KEYINPUT51), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(KEYINPUT51), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1075), .A2(new_n1076), .B1(G50), .B2(new_n763), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n766), .A2(new_n223), .B1(new_n774), .B2(new_n955), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1078), .A2(KEYINPUT118), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n759), .A2(new_n286), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n829), .B(new_n1080), .C1(new_n1078), .C2(KEYINPUT118), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n254), .B1(new_n794), .B2(G77), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1077), .A2(new_n1079), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT119), .Z(new_n1084));
  AOI22_X1  g0884(.A1(new_n763), .A2(G303), .B1(new_n794), .B2(G116), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n784), .B2(new_n774), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(G283), .B2(new_n846), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n257), .B1(new_n791), .B2(G294), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n769), .A2(new_n964), .B1(new_n770), .B2(new_n960), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT52), .ZN(new_n1090));
  AND4_X1   g0890(.A1(new_n755), .A2(new_n1087), .A3(new_n1088), .A4(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n798), .B1(new_n1084), .B2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1072), .A2(new_n854), .A3(new_n1073), .A4(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1071), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1007), .A2(new_n1002), .A3(new_n1009), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT110), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1095), .B1(new_n1098), .B2(new_n1010), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1094), .B1(new_n1099), .B2(new_n696), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(G390));
  NAND2_X1  g0901(.A1(new_n936), .A2(new_n938), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n900), .B1(new_n823), .B2(new_n923), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1102), .B1(new_n1103), .B2(new_n940), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n893), .A2(new_n940), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n899), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n732), .A2(new_n670), .A3(new_n818), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n819), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1105), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n721), .A2(new_n900), .A3(G330), .A4(new_n821), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NOR3_X1   g0911(.A1(new_n1104), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n901), .A2(new_n741), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n900), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n644), .A2(new_n692), .A3(new_n821), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n819), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n939), .B1(new_n1117), .B2(new_n897), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n893), .A2(new_n940), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1107), .A2(new_n819), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1119), .B1(new_n1120), .B2(new_n899), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1114), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1112), .A2(new_n1122), .ZN(new_n1123));
  XOR2_X1   g0923(.A(KEYINPUT54), .B(G143), .Z(new_n1124));
  AOI22_X1  g0924(.A1(G132), .A2(new_n831), .B1(new_n791), .B2(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n793), .A2(G128), .B1(new_n794), .B2(G159), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1125), .B(new_n1126), .C1(new_n202), .C2(new_n753), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1028), .A2(new_n766), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(new_n1128), .B(KEYINPUT53), .ZN(new_n1129));
  INV_X1    g0929(.A(G125), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1129), .B(new_n257), .C1(new_n1130), .C2(new_n774), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1127), .B(new_n1131), .C1(G137), .C2(new_n763), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(G294), .A2(new_n777), .B1(new_n794), .B2(G77), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n1133), .B1(new_n220), .B2(new_n770), .C1(new_n786), .C2(new_n769), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n254), .B1(new_n759), .B2(new_n210), .C1(new_n490), .C2(new_n762), .ZN(new_n1135));
  NOR4_X1   g0935(.A1(new_n1134), .A2(new_n767), .A3(new_n845), .A4(new_n1135), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1132), .A2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1137), .A2(new_n750), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1102), .A2(new_n800), .ZN(new_n1139));
  AOI211_X1 g0939(.A(new_n1138), .B(new_n1139), .C1(new_n286), .C2(new_n851), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1123), .A2(new_n980), .B1(new_n854), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n425), .A2(G330), .A3(new_n896), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n919), .A2(new_n1142), .A3(new_n655), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n823), .A2(new_n923), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT120), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n721), .A2(G330), .A3(new_n821), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1146), .B1(new_n1147), .B2(new_n1115), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1148), .A2(new_n1113), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1147), .A2(new_n1146), .A3(new_n1115), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1145), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n896), .A2(G330), .A3(new_n821), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n1115), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1120), .A2(new_n1153), .A3(new_n1110), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1144), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1113), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1118), .A2(new_n1121), .A3(new_n1110), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n696), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1154), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1147), .A2(new_n1146), .A3(new_n1115), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n1161), .A2(new_n1148), .A3(new_n1113), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1160), .B1(new_n1162), .B2(new_n1145), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1163), .A2(new_n1144), .B1(new_n1157), .B2(new_n1156), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1141), .B1(new_n1159), .B2(new_n1164), .ZN(G378));
  INV_X1    g0965(.A(KEYINPUT57), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n651), .A2(new_n301), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n925), .A2(new_n297), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT55), .Z(new_n1169));
  NAND2_X1  g0969(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1169), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n651), .A2(new_n301), .A3(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1171), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1172), .B1(new_n651), .B2(new_n301), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n302), .B(new_n1169), .C1(new_n650), .C2(new_n647), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1174), .A2(new_n1178), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n908), .A2(new_n941), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n908), .A2(new_n941), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1179), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n926), .B1(new_n1102), .B2(new_n897), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n924), .B(new_n1183), .C1(new_n915), .C2(new_n741), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n1174), .A2(new_n1178), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n908), .A2(new_n941), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1182), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1143), .B1(new_n1123), .B2(new_n1163), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1166), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1147), .A2(new_n1115), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(KEYINPUT120), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1192), .A2(new_n1114), .A3(new_n1150), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1145), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1154), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1144), .B1(new_n1158), .B2(new_n1195), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1196), .A2(KEYINPUT57), .A3(new_n1187), .A4(new_n1182), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1190), .A2(new_n696), .A3(new_n1197), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1182), .A2(new_n1187), .A3(new_n980), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n202), .B1(new_n252), .B2(G41), .ZN(new_n1200));
  AOI21_X1  g1000(.A(G41), .B1(new_n777), .B2(G124), .ZN(new_n1201));
  AOI21_X1  g1001(.A(G33), .B1(new_n754), .B2(G159), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n769), .A2(new_n1130), .B1(new_n757), .B2(new_n283), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n831), .A2(G128), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n759), .B2(new_n839), .C1(new_n843), .C2(new_n762), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n1203), .B(new_n1205), .C1(new_n846), .C2(new_n1124), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT59), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1201), .B(new_n1202), .C1(new_n1206), .C2(new_n1207), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1200), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n763), .A2(G97), .B1(new_n777), .B2(G283), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1211), .B(new_n1034), .C1(new_n490), .C2(new_n770), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n404), .A2(new_n791), .B1(new_n754), .B2(G58), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n257), .B1(new_n793), .B2(G116), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1213), .A2(new_n953), .A3(new_n1214), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n1212), .A2(new_n1215), .A3(G41), .ZN(new_n1216));
  XOR2_X1   g1016(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n1217));
  XNOR2_X1  g1017(.A(new_n1216), .B(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1210), .A2(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1219), .A2(new_n750), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n744), .B(new_n1220), .C1(new_n202), .C2(new_n851), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n1185), .B2(new_n800), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1199), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1198), .A2(new_n1224), .ZN(G375));
  NAND2_X1  g1025(.A1(new_n1115), .A2(new_n799), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n763), .A2(new_n1124), .B1(new_n777), .B2(G128), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1227), .B(new_n257), .C1(new_n283), .C2(new_n759), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G159), .A2(new_n846), .B1(new_n754), .B2(G58), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n843), .B2(new_n769), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n770), .A2(new_n839), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n757), .A2(new_n202), .ZN(new_n1232));
  NOR4_X1   g1032(.A1(new_n1228), .A2(new_n1230), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(G77), .A2(new_n754), .B1(new_n794), .B2(new_n404), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n490), .B2(new_n759), .ZN(new_n1235));
  OAI221_X1 g1035(.A(new_n254), .B1(new_n774), .B2(new_n781), .C1(new_n786), .C2(new_n770), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n762), .A2(new_n220), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n769), .A2(new_n966), .B1(new_n766), .B2(new_n210), .ZN(new_n1238));
  NOR4_X1   g1038(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n798), .B1(new_n1233), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n851), .A2(new_n223), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1226), .A2(new_n854), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n1195), .B2(new_n1061), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1195), .A2(new_n1143), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1160), .B(new_n1143), .C1(new_n1162), .C2(new_n1145), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT123), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1195), .A2(KEYINPUT123), .A3(new_n1143), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1244), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1243), .B1(new_n1249), .B2(new_n1013), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(G381));
  INV_X1    g1051(.A(G396), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1067), .A2(new_n1252), .A3(new_n1069), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n857), .B2(new_n856), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(new_n1254), .B(KEYINPUT124), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1196), .A2(new_n1187), .A3(new_n1182), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n697), .B1(new_n1256), .B2(new_n1166), .ZN(new_n1257));
  AOI211_X1 g1057(.A(G378), .B(new_n1223), .C1(new_n1257), .C2(new_n1197), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1255), .A2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n979), .B(new_n1100), .C1(new_n1014), .C2(new_n1026), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n1250), .ZN(new_n1262));
  OR2_X1    g1062(.A1(new_n1259), .A2(new_n1262), .ZN(G407));
  INV_X1    g1063(.A(G378), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1198), .A2(new_n1264), .A3(new_n1224), .ZN(new_n1265));
  OAI221_X1 g1065(.A(G213), .B1(G343), .B2(new_n1265), .C1(new_n1259), .C2(new_n1262), .ZN(G409));
  AOI21_X1  g1066(.A(new_n1264), .B1(new_n1198), .B2(new_n1224), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n668), .A2(G213), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1013), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1199), .B(new_n1222), .C1(new_n1256), .C2(new_n1269), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1268), .B1(new_n1270), .B2(G378), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1267), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1243), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT125), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(new_n856), .B2(new_n857), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1247), .A2(new_n1248), .B1(new_n1155), .B2(KEYINPUT60), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT60), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n696), .B1(new_n1245), .B2(new_n1277), .ZN(new_n1278));
  OAI211_X1 g1078(.A(new_n1273), .B(new_n1275), .C1(new_n1276), .C2(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT123), .B1(new_n1195), .B2(new_n1143), .ZN(new_n1281));
  OAI22_X1  g1081(.A1(new_n1280), .A2(new_n1281), .B1(new_n1244), .B2(new_n1277), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1278), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1243), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  XNOR2_X1  g1084(.A(G384), .B(new_n1274), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1279), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(KEYINPUT63), .B1(new_n1272), .B2(new_n1287), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT63), .ZN(new_n1289));
  NOR4_X1   g1089(.A1(new_n1267), .A2(new_n1286), .A3(new_n1271), .A4(new_n1289), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1288), .A2(new_n1290), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1252), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1292));
  OR2_X1    g1092(.A1(new_n1253), .A2(new_n1292), .ZN(new_n1293));
  AND2_X1   g1093(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1098), .A2(new_n1010), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1269), .B1(new_n1295), .B2(new_n736), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1294), .B1(new_n1296), .B2(new_n980), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1100), .B1(new_n1297), .B2(new_n979), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1293), .B1(new_n1261), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G387), .A2(G390), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1253), .A2(new_n1292), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1300), .A2(new_n1260), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT61), .ZN(new_n1304));
  OR2_X1    g1104(.A1(new_n1267), .A2(new_n1271), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n668), .A2(G213), .A3(G2897), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1287), .A2(new_n1307), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1307), .B(new_n1279), .C1(new_n1284), .C2(new_n1285), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1305), .B1(new_n1308), .B2(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1291), .A2(new_n1303), .A3(new_n1304), .A4(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(KEYINPUT62), .B1(new_n1305), .B2(new_n1286), .ZN(new_n1313));
  XOR2_X1   g1113(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1314));
  INV_X1    g1114(.A(KEYINPUT62), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1272), .A2(new_n1315), .A3(new_n1287), .ZN(new_n1316));
  AND4_X1   g1116(.A1(new_n1311), .A2(new_n1313), .A3(new_n1314), .A4(new_n1316), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1312), .B1(new_n1317), .B2(new_n1303), .ZN(G405));
  NAND2_X1  g1118(.A1(G375), .A2(G378), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1319), .A2(new_n1265), .A3(new_n1286), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1287), .B1(new_n1258), .B2(new_n1267), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1299), .A2(new_n1322), .A3(new_n1302), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(KEYINPUT127), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1322), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1303), .A2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT127), .ZN(new_n1327));
  NAND4_X1  g1127(.A1(new_n1299), .A2(new_n1322), .A3(new_n1302), .A4(new_n1327), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1324), .A2(new_n1326), .A3(new_n1328), .ZN(G402));
endmodule


