

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604;

  NOR2_X1 U325 ( .A1(n500), .A2(n602), .ZN(n481) );
  XNOR2_X1 U326 ( .A(n350), .B(KEYINPUT95), .ZN(n351) );
  XNOR2_X1 U327 ( .A(n385), .B(n293), .ZN(n386) );
  XNOR2_X1 U328 ( .A(n348), .B(n347), .ZN(n488) );
  XNOR2_X1 U329 ( .A(KEYINPUT103), .B(KEYINPUT38), .ZN(n463) );
  INV_X1 U330 ( .A(n504), .ZN(n461) );
  AND2_X1 U331 ( .A1(G232GAT), .A2(G233GAT), .ZN(n293) );
  XOR2_X1 U332 ( .A(n449), .B(n359), .Z(n294) );
  AND2_X1 U333 ( .A1(n417), .A2(n500), .ZN(n295) );
  INV_X1 U334 ( .A(KEYINPUT25), .ZN(n350) );
  NOR2_X1 U335 ( .A1(n473), .A2(n581), .ZN(n474) );
  INV_X1 U336 ( .A(KEYINPUT33), .ZN(n440) );
  XNOR2_X1 U337 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U338 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U339 ( .A(n433), .B(n386), .ZN(n387) );
  XNOR2_X1 U340 ( .A(n389), .B(n454), .ZN(n390) );
  XNOR2_X1 U341 ( .A(n388), .B(n334), .ZN(n335) );
  INV_X1 U342 ( .A(n452), .ZN(n456) );
  XNOR2_X1 U343 ( .A(n391), .B(n390), .ZN(n393) );
  XNOR2_X1 U344 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U345 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U346 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U347 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U348 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U349 ( .A(n464), .B(n463), .ZN(n518) );
  XNOR2_X1 U350 ( .A(n497), .B(G176GAT), .ZN(n498) );
  XNOR2_X1 U351 ( .A(n467), .B(G43GAT), .ZN(n468) );
  XNOR2_X1 U352 ( .A(n469), .B(n468), .ZN(G1330GAT) );
  XOR2_X1 U353 ( .A(KEYINPUT102), .B(KEYINPUT37), .Z(n419) );
  XOR2_X1 U354 ( .A(KEYINPUT17), .B(KEYINPUT86), .Z(n297) );
  XNOR2_X1 U355 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n296) );
  XNOR2_X1 U356 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U357 ( .A(KEYINPUT19), .B(n298), .Z(n336) );
  XOR2_X1 U358 ( .A(G120GAT), .B(G71GAT), .Z(n449) );
  XOR2_X1 U359 ( .A(G127GAT), .B(KEYINPUT81), .Z(n300) );
  XNOR2_X1 U360 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n299) );
  XNOR2_X1 U361 ( .A(n300), .B(n299), .ZN(n359) );
  NAND2_X1 U362 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U363 ( .A(n294), .B(n301), .ZN(n313) );
  XOR2_X1 U364 ( .A(G99GAT), .B(G190GAT), .Z(n303) );
  XNOR2_X1 U365 ( .A(G43GAT), .B(G113GAT), .ZN(n302) );
  XNOR2_X1 U366 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U367 ( .A(KEYINPUT82), .B(G176GAT), .Z(n305) );
  XNOR2_X1 U368 ( .A(G169GAT), .B(G15GAT), .ZN(n304) );
  XNOR2_X1 U369 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U370 ( .A(n307), .B(n306), .Z(n311) );
  XOR2_X1 U371 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n309) );
  XNOR2_X1 U372 ( .A(KEYINPUT85), .B(KEYINPUT83), .ZN(n308) );
  XNOR2_X1 U373 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U374 ( .A(n336), .B(n314), .Z(n539) );
  INV_X1 U375 ( .A(n539), .ZN(n547) );
  XOR2_X1 U376 ( .A(G211GAT), .B(KEYINPUT87), .Z(n316) );
  XNOR2_X1 U377 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n315) );
  XNOR2_X1 U378 ( .A(n316), .B(n315), .ZN(n344) );
  XOR2_X1 U379 ( .A(KEYINPUT69), .B(G78GAT), .Z(n318) );
  XNOR2_X1 U380 ( .A(G148GAT), .B(G106GAT), .ZN(n317) );
  XNOR2_X1 U381 ( .A(n318), .B(n317), .ZN(n452) );
  XNOR2_X1 U382 ( .A(n344), .B(n452), .ZN(n330) );
  XOR2_X1 U383 ( .A(KEYINPUT88), .B(KEYINPUT3), .Z(n320) );
  XNOR2_X1 U384 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n319) );
  XNOR2_X1 U385 ( .A(n320), .B(n319), .ZN(n355) );
  XOR2_X1 U386 ( .A(n355), .B(KEYINPUT23), .Z(n322) );
  NAND2_X1 U387 ( .A1(G228GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U388 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U389 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n324) );
  XNOR2_X1 U390 ( .A(G204GAT), .B(G218GAT), .ZN(n323) );
  XNOR2_X1 U391 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U392 ( .A(n326), .B(n325), .Z(n328) );
  XOR2_X1 U393 ( .A(G50GAT), .B(G162GAT), .Z(n385) );
  XOR2_X1 U394 ( .A(G22GAT), .B(G155GAT), .Z(n403) );
  XNOR2_X1 U395 ( .A(n385), .B(n403), .ZN(n327) );
  XNOR2_X1 U396 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U397 ( .A(n330), .B(n329), .ZN(n493) );
  NAND2_X1 U398 ( .A1(n547), .A2(n493), .ZN(n331) );
  XNOR2_X1 U399 ( .A(n331), .B(KEYINPUT26), .ZN(n332) );
  XOR2_X1 U400 ( .A(KEYINPUT94), .B(n332), .Z(n565) );
  XOR2_X1 U401 ( .A(G169GAT), .B(G8GAT), .Z(n424) );
  XNOR2_X1 U402 ( .A(G36GAT), .B(G190GAT), .ZN(n333) );
  XNOR2_X1 U403 ( .A(n333), .B(G218GAT), .ZN(n388) );
  XOR2_X1 U404 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n334) );
  XOR2_X1 U405 ( .A(n424), .B(n337), .Z(n348) );
  INV_X1 U406 ( .A(G204GAT), .ZN(n338) );
  NAND2_X1 U407 ( .A1(n338), .A2(G64GAT), .ZN(n341) );
  INV_X1 U408 ( .A(G64GAT), .ZN(n339) );
  NAND2_X1 U409 ( .A1(n339), .A2(G204GAT), .ZN(n340) );
  NAND2_X1 U410 ( .A1(n341), .A2(n340), .ZN(n343) );
  XNOR2_X1 U411 ( .A(G176GAT), .B(G92GAT), .ZN(n342) );
  XNOR2_X1 U412 ( .A(n343), .B(n342), .ZN(n443) );
  XNOR2_X1 U413 ( .A(n443), .B(n344), .ZN(n346) );
  NAND2_X1 U414 ( .A1(G226GAT), .A2(G233GAT), .ZN(n345) );
  INV_X1 U415 ( .A(n488), .ZN(n537) );
  XNOR2_X1 U416 ( .A(n537), .B(KEYINPUT27), .ZN(n376) );
  NAND2_X1 U417 ( .A1(n565), .A2(n376), .ZN(n354) );
  NOR2_X1 U418 ( .A1(n488), .A2(n547), .ZN(n349) );
  NOR2_X1 U419 ( .A1(n493), .A2(n349), .ZN(n352) );
  NAND2_X1 U420 ( .A1(n354), .A2(n353), .ZN(n374) );
  XOR2_X1 U421 ( .A(G113GAT), .B(G1GAT), .Z(n425) );
  XOR2_X1 U422 ( .A(n355), .B(n425), .Z(n357) );
  NAND2_X1 U423 ( .A1(G225GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U424 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U425 ( .A(n358), .B(G57GAT), .Z(n361) );
  XNOR2_X1 U426 ( .A(n359), .B(G120GAT), .ZN(n360) );
  XNOR2_X1 U427 ( .A(n361), .B(n360), .ZN(n365) );
  XOR2_X1 U428 ( .A(KEYINPUT6), .B(G85GAT), .Z(n363) );
  XNOR2_X1 U429 ( .A(G29GAT), .B(G162GAT), .ZN(n362) );
  XNOR2_X1 U430 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U431 ( .A(n365), .B(n364), .Z(n373) );
  XOR2_X1 U432 ( .A(G155GAT), .B(KEYINPUT89), .Z(n367) );
  XNOR2_X1 U433 ( .A(KEYINPUT90), .B(KEYINPUT5), .ZN(n366) );
  XNOR2_X1 U434 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U435 ( .A(KEYINPUT91), .B(G148GAT), .Z(n369) );
  XNOR2_X1 U436 ( .A(KEYINPUT4), .B(KEYINPUT1), .ZN(n368) );
  XNOR2_X1 U437 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U438 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U439 ( .A(n373), .B(n372), .Z(n491) );
  NAND2_X1 U440 ( .A1(n374), .A2(n491), .ZN(n375) );
  XNOR2_X1 U441 ( .A(n375), .B(KEYINPUT96), .ZN(n379) );
  XNOR2_X1 U442 ( .A(n493), .B(KEYINPUT28), .ZN(n550) );
  INV_X1 U443 ( .A(n491), .ZN(n534) );
  NAND2_X1 U444 ( .A1(n534), .A2(n376), .ZN(n545) );
  NOR2_X1 U445 ( .A1(n550), .A2(n545), .ZN(n377) );
  NAND2_X1 U446 ( .A1(n377), .A2(n547), .ZN(n378) );
  NAND2_X1 U447 ( .A1(n379), .A2(n378), .ZN(n380) );
  XOR2_X1 U448 ( .A(KEYINPUT97), .B(n380), .Z(n502) );
  XOR2_X1 U449 ( .A(KEYINPUT9), .B(G106GAT), .Z(n382) );
  XNOR2_X1 U450 ( .A(KEYINPUT11), .B(KEYINPUT10), .ZN(n381) );
  XNOR2_X1 U451 ( .A(n382), .B(n381), .ZN(n395) );
  XOR2_X1 U452 ( .A(G29GAT), .B(G43GAT), .Z(n384) );
  XNOR2_X1 U453 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n383) );
  XNOR2_X1 U454 ( .A(n384), .B(n383), .ZN(n433) );
  XNOR2_X1 U455 ( .A(n387), .B(KEYINPUT74), .ZN(n391) );
  XNOR2_X1 U456 ( .A(n388), .B(KEYINPUT75), .ZN(n389) );
  XOR2_X1 U457 ( .A(G99GAT), .B(G85GAT), .Z(n454) );
  XNOR2_X1 U458 ( .A(G134GAT), .B(G92GAT), .ZN(n392) );
  XNOR2_X1 U459 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U460 ( .A(n395), .B(n394), .ZN(n472) );
  INV_X1 U461 ( .A(KEYINPUT36), .ZN(n396) );
  XNOR2_X1 U462 ( .A(n472), .B(n396), .ZN(n602) );
  INV_X1 U463 ( .A(n602), .ZN(n417) );
  XOR2_X1 U464 ( .A(G64GAT), .B(G127GAT), .Z(n398) );
  XNOR2_X1 U465 ( .A(G1GAT), .B(G183GAT), .ZN(n397) );
  XNOR2_X1 U466 ( .A(n398), .B(n397), .ZN(n402) );
  XOR2_X1 U467 ( .A(G78GAT), .B(G211GAT), .Z(n400) );
  XNOR2_X1 U468 ( .A(G8GAT), .B(G71GAT), .ZN(n399) );
  XNOR2_X1 U469 ( .A(n400), .B(n399), .ZN(n401) );
  XOR2_X1 U470 ( .A(n402), .B(n401), .Z(n408) );
  XOR2_X1 U471 ( .A(G57GAT), .B(KEYINPUT13), .Z(n453) );
  XOR2_X1 U472 ( .A(n403), .B(KEYINPUT80), .Z(n405) );
  NAND2_X1 U473 ( .A1(G231GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U474 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U475 ( .A(n453), .B(n406), .ZN(n407) );
  XNOR2_X1 U476 ( .A(n408), .B(n407), .ZN(n416) );
  XOR2_X1 U477 ( .A(KEYINPUT14), .B(KEYINPUT15), .Z(n410) );
  XNOR2_X1 U478 ( .A(G15GAT), .B(KEYINPUT76), .ZN(n409) );
  XNOR2_X1 U479 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U480 ( .A(KEYINPUT79), .B(KEYINPUT77), .Z(n412) );
  XNOR2_X1 U481 ( .A(KEYINPUT78), .B(KEYINPUT12), .ZN(n411) );
  XNOR2_X1 U482 ( .A(n412), .B(n411), .ZN(n413) );
  XOR2_X1 U483 ( .A(n414), .B(n413), .Z(n415) );
  XOR2_X1 U484 ( .A(n416), .B(n415), .Z(n500) );
  NAND2_X1 U485 ( .A1(n502), .A2(n295), .ZN(n418) );
  XNOR2_X1 U486 ( .A(n419), .B(n418), .ZN(n533) );
  INV_X1 U487 ( .A(n533), .ZN(n462) );
  XOR2_X1 U488 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n421) );
  XNOR2_X1 U489 ( .A(G141GAT), .B(G197GAT), .ZN(n420) );
  XNOR2_X1 U490 ( .A(n421), .B(n420), .ZN(n437) );
  XOR2_X1 U491 ( .A(KEYINPUT67), .B(G22GAT), .Z(n423) );
  XNOR2_X1 U492 ( .A(G15GAT), .B(KEYINPUT68), .ZN(n422) );
  XNOR2_X1 U493 ( .A(n423), .B(n422), .ZN(n429) );
  XOR2_X1 U494 ( .A(G50GAT), .B(G36GAT), .Z(n427) );
  XNOR2_X1 U495 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U496 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U497 ( .A(n429), .B(n428), .Z(n431) );
  NAND2_X1 U498 ( .A1(G229GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U499 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U500 ( .A(n432), .B(KEYINPUT66), .Z(n435) );
  XNOR2_X1 U501 ( .A(n433), .B(KEYINPUT65), .ZN(n434) );
  XNOR2_X1 U502 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U503 ( .A(n437), .B(n436), .ZN(n520) );
  INV_X1 U504 ( .A(n520), .ZN(n589) );
  XOR2_X1 U505 ( .A(KEYINPUT71), .B(KEYINPUT72), .Z(n439) );
  XNOR2_X1 U506 ( .A(KEYINPUT32), .B(KEYINPUT73), .ZN(n438) );
  XNOR2_X1 U507 ( .A(n439), .B(n438), .ZN(n460) );
  NAND2_X1 U508 ( .A1(G230GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U509 ( .A(n443), .B(n442), .ZN(n446) );
  INV_X1 U510 ( .A(n446), .ZN(n444) );
  NAND2_X1 U511 ( .A1(n444), .A2(KEYINPUT70), .ZN(n448) );
  INV_X1 U512 ( .A(KEYINPUT70), .ZN(n445) );
  NAND2_X1 U513 ( .A1(n446), .A2(n445), .ZN(n447) );
  NAND2_X1 U514 ( .A1(n448), .A2(n447), .ZN(n451) );
  XNOR2_X1 U515 ( .A(n449), .B(KEYINPUT31), .ZN(n450) );
  XNOR2_X1 U516 ( .A(n451), .B(n450), .ZN(n458) );
  XNOR2_X1 U517 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U518 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X1 U519 ( .A(n460), .B(n459), .Z(n594) );
  NAND2_X1 U520 ( .A1(n589), .A2(n594), .ZN(n504) );
  NAND2_X1 U521 ( .A1(n462), .A2(n461), .ZN(n464) );
  NAND2_X1 U522 ( .A1(n518), .A2(n537), .ZN(n466) );
  XNOR2_X1 U523 ( .A(G36GAT), .B(KEYINPUT104), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n466), .B(n465), .ZN(G1329GAT) );
  NAND2_X1 U525 ( .A1(n539), .A2(n518), .ZN(n469) );
  XOR2_X1 U526 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n467) );
  INV_X1 U527 ( .A(KEYINPUT41), .ZN(n470) );
  XNOR2_X1 U528 ( .A(n594), .B(n470), .ZN(n571) );
  XOR2_X1 U529 ( .A(n571), .B(KEYINPUT106), .Z(n554) );
  NOR2_X1 U530 ( .A1(n571), .A2(n520), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n471), .B(KEYINPUT46), .ZN(n473) );
  BUF_X1 U532 ( .A(n472), .Z(n581) );
  INV_X1 U533 ( .A(n500), .ZN(n597) );
  NAND2_X1 U534 ( .A1(n474), .A2(n500), .ZN(n477) );
  INV_X1 U535 ( .A(n477), .ZN(n476) );
  XOR2_X1 U536 ( .A(KEYINPUT47), .B(KEYINPUT111), .Z(n478) );
  INV_X1 U537 ( .A(n478), .ZN(n475) );
  NAND2_X1 U538 ( .A1(n476), .A2(n475), .ZN(n480) );
  NAND2_X1 U539 ( .A1(n478), .A2(n477), .ZN(n479) );
  NAND2_X1 U540 ( .A1(n480), .A2(n479), .ZN(n486) );
  XNOR2_X1 U541 ( .A(n481), .B(KEYINPUT45), .ZN(n482) );
  NAND2_X1 U542 ( .A1(n482), .A2(n594), .ZN(n483) );
  NOR2_X1 U543 ( .A1(n589), .A2(n483), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n484), .B(KEYINPUT112), .ZN(n485) );
  NOR2_X1 U545 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U546 ( .A(KEYINPUT48), .B(n487), .ZN(n544) );
  NOR2_X1 U547 ( .A1(n544), .A2(n488), .ZN(n489) );
  XNOR2_X1 U548 ( .A(KEYINPUT54), .B(n489), .ZN(n490) );
  AND2_X1 U549 ( .A1(n491), .A2(n490), .ZN(n492) );
  XOR2_X1 U550 ( .A(KEYINPUT64), .B(n492), .Z(n588) );
  NOR2_X1 U551 ( .A1(n588), .A2(n493), .ZN(n494) );
  XNOR2_X1 U552 ( .A(n494), .B(KEYINPUT55), .ZN(n495) );
  NOR2_X2 U553 ( .A1(n547), .A2(n495), .ZN(n496) );
  XOR2_X2 U554 ( .A(KEYINPUT123), .B(n496), .Z(n582) );
  NAND2_X1 U555 ( .A1(n554), .A2(n582), .ZN(n499) );
  XOR2_X1 U556 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n497) );
  XNOR2_X1 U557 ( .A(n499), .B(n498), .ZN(G1349GAT) );
  NOR2_X1 U558 ( .A1(n500), .A2(n581), .ZN(n501) );
  XNOR2_X1 U559 ( .A(n501), .B(KEYINPUT16), .ZN(n503) );
  NAND2_X1 U560 ( .A1(n503), .A2(n502), .ZN(n522) );
  NOR2_X1 U561 ( .A1(n504), .A2(n522), .ZN(n513) );
  NAND2_X1 U562 ( .A1(n513), .A2(n534), .ZN(n505) );
  XNOR2_X1 U563 ( .A(n505), .B(KEYINPUT34), .ZN(n506) );
  XNOR2_X1 U564 ( .A(G1GAT), .B(n506), .ZN(G1324GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n508) );
  NAND2_X1 U566 ( .A1(n513), .A2(n537), .ZN(n507) );
  XNOR2_X1 U567 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U568 ( .A(G8GAT), .B(n509), .ZN(G1325GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT35), .B(KEYINPUT100), .Z(n511) );
  NAND2_X1 U570 ( .A1(n513), .A2(n539), .ZN(n510) );
  XNOR2_X1 U571 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U572 ( .A(G15GAT), .B(n512), .ZN(G1326GAT) );
  XOR2_X1 U573 ( .A(G22GAT), .B(KEYINPUT101), .Z(n515) );
  NAND2_X1 U574 ( .A1(n513), .A2(n550), .ZN(n514) );
  XNOR2_X1 U575 ( .A(n515), .B(n514), .ZN(G1327GAT) );
  XOR2_X1 U576 ( .A(G29GAT), .B(KEYINPUT39), .Z(n517) );
  NAND2_X1 U577 ( .A1(n534), .A2(n518), .ZN(n516) );
  XNOR2_X1 U578 ( .A(n517), .B(n516), .ZN(G1328GAT) );
  NAND2_X1 U579 ( .A1(n518), .A2(n550), .ZN(n519) );
  XNOR2_X1 U580 ( .A(n519), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U581 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n524) );
  NAND2_X1 U582 ( .A1(n520), .A2(n554), .ZN(n521) );
  XOR2_X1 U583 ( .A(KEYINPUT107), .B(n521), .Z(n532) );
  NOR2_X1 U584 ( .A1(n532), .A2(n522), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n534), .A2(n528), .ZN(n523) );
  XNOR2_X1 U586 ( .A(n524), .B(n523), .ZN(G1332GAT) );
  NAND2_X1 U587 ( .A1(n537), .A2(n528), .ZN(n525) );
  XNOR2_X1 U588 ( .A(n525), .B(KEYINPUT108), .ZN(n526) );
  XNOR2_X1 U589 ( .A(G64GAT), .B(n526), .ZN(G1333GAT) );
  NAND2_X1 U590 ( .A1(n528), .A2(n539), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n527), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n530) );
  NAND2_X1 U593 ( .A1(n528), .A2(n550), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U595 ( .A(G78GAT), .B(n531), .Z(G1335GAT) );
  NOR2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n534), .A2(n541), .ZN(n535) );
  XNOR2_X1 U598 ( .A(KEYINPUT110), .B(n535), .ZN(n536) );
  XNOR2_X1 U599 ( .A(G85GAT), .B(n536), .ZN(G1336GAT) );
  NAND2_X1 U600 ( .A1(n537), .A2(n541), .ZN(n538) );
  XNOR2_X1 U601 ( .A(n538), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U602 ( .A1(n541), .A2(n539), .ZN(n540) );
  XNOR2_X1 U603 ( .A(n540), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U604 ( .A1(n550), .A2(n541), .ZN(n542) );
  XNOR2_X1 U605 ( .A(n542), .B(KEYINPUT44), .ZN(n543) );
  XNOR2_X1 U606 ( .A(G106GAT), .B(n543), .ZN(G1339GAT) );
  XOR2_X1 U607 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n552) );
  NOR2_X1 U608 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U609 ( .A(n546), .B(KEYINPUT113), .ZN(n566) );
  NOR2_X1 U610 ( .A1(n547), .A2(n566), .ZN(n548) );
  XOR2_X1 U611 ( .A(KEYINPUT114), .B(n548), .Z(n549) );
  NOR2_X1 U612 ( .A1(n550), .A2(n549), .ZN(n561) );
  NAND2_X1 U613 ( .A1(n561), .A2(n589), .ZN(n551) );
  XNOR2_X1 U614 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U615 ( .A(G113GAT), .B(n553), .ZN(G1340GAT) );
  XOR2_X1 U616 ( .A(G120GAT), .B(KEYINPUT49), .Z(n556) );
  NAND2_X1 U617 ( .A1(n561), .A2(n554), .ZN(n555) );
  XNOR2_X1 U618 ( .A(n556), .B(n555), .ZN(G1341GAT) );
  XNOR2_X1 U619 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n560) );
  XOR2_X1 U620 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n558) );
  NAND2_X1 U621 ( .A1(n561), .A2(n597), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U623 ( .A(n560), .B(n559), .ZN(G1342GAT) );
  XOR2_X1 U624 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n563) );
  NAND2_X1 U625 ( .A1(n561), .A2(n581), .ZN(n562) );
  XNOR2_X1 U626 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U627 ( .A(G134GAT), .B(n564), .Z(G1343GAT) );
  INV_X1 U628 ( .A(n565), .ZN(n587) );
  NOR2_X1 U629 ( .A1(n566), .A2(n587), .ZN(n577) );
  NAND2_X1 U630 ( .A1(n589), .A2(n577), .ZN(n567) );
  XNOR2_X1 U631 ( .A(G141GAT), .B(n567), .ZN(G1344GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT122), .B(KEYINPUT53), .Z(n569) );
  XNOR2_X1 U633 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n575) );
  INV_X1 U635 ( .A(n577), .ZN(n570) );
  NOR2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n573) );
  XNOR2_X1 U637 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n575), .B(n574), .ZN(G1345GAT) );
  NAND2_X1 U640 ( .A1(n597), .A2(n577), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U642 ( .A1(n581), .A2(n577), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U644 ( .A1(n589), .A2(n582), .ZN(n579) );
  XNOR2_X1 U645 ( .A(G169GAT), .B(n579), .ZN(G1348GAT) );
  NAND2_X1 U646 ( .A1(n597), .A2(n582), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n580), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U648 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n584) );
  NAND2_X1 U649 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(G1351GAT) );
  XOR2_X1 U651 ( .A(KEYINPUT126), .B(KEYINPUT60), .Z(n586) );
  XNOR2_X1 U652 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n585) );
  XNOR2_X1 U653 ( .A(n586), .B(n585), .ZN(n593) );
  XOR2_X1 U654 ( .A(G197GAT), .B(KEYINPUT59), .Z(n591) );
  NOR2_X1 U655 ( .A1(n588), .A2(n587), .ZN(n598) );
  NAND2_X1 U656 ( .A1(n598), .A2(n589), .ZN(n590) );
  XNOR2_X1 U657 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U658 ( .A(n593), .B(n592), .ZN(G1352GAT) );
  XOR2_X1 U659 ( .A(G204GAT), .B(KEYINPUT61), .Z(n596) );
  INV_X1 U660 ( .A(n598), .ZN(n601) );
  OR2_X1 U661 ( .A1(n601), .A2(n594), .ZN(n595) );
  XNOR2_X1 U662 ( .A(n596), .B(n595), .ZN(G1353GAT) );
  XOR2_X1 U663 ( .A(G211GAT), .B(KEYINPUT127), .Z(n600) );
  NAND2_X1 U664 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U665 ( .A(n600), .B(n599), .ZN(G1354GAT) );
  NOR2_X1 U666 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U667 ( .A(KEYINPUT62), .B(n603), .Z(n604) );
  XNOR2_X1 U668 ( .A(G218GAT), .B(n604), .ZN(G1355GAT) );
endmodule

