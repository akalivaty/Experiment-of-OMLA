//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n602, new_n603,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n820, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n849, new_n850, new_n851;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n202));
  NAND2_X1  g001(.A1(G227gat), .A2(G233gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT72), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT24), .ZN(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G183gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT65), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT65), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G183gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G190gat), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n208), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n206), .A2(new_n207), .A3(new_n205), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n218), .A2(KEYINPUT23), .ZN(new_n219));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(KEYINPUT23), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  AND3_X1   g021(.A1(new_n217), .A2(KEYINPUT25), .A3(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n224), .B1(new_n205), .B2(new_n206), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(new_n205), .B2(new_n206), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT25), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n229));
  NOR2_X1   g028(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n230));
  XNOR2_X1  g029(.A(KEYINPUT65), .B(G183gat), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n230), .B1(new_n231), .B2(KEYINPUT27), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n229), .B1(new_n232), .B2(G190gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT28), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n210), .A2(new_n212), .A3(KEYINPUT27), .ZN(new_n235));
  INV_X1    g034(.A(new_n230), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n237), .A2(KEYINPUT66), .A3(new_n214), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n233), .A2(new_n234), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n233), .A2(KEYINPUT67), .A3(new_n234), .A4(new_n238), .ZN(new_n242));
  XOR2_X1   g041(.A(KEYINPUT27), .B(G183gat), .Z(new_n243));
  OR3_X1    g042(.A1(new_n243), .A2(new_n234), .A3(G190gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n241), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n218), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n247));
  OR3_X1    g046(.A1(new_n246), .A2(new_n247), .A3(KEYINPUT26), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n247), .B1(new_n246), .B2(KEYINPUT26), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n248), .A2(new_n249), .B1(KEYINPUT26), .B2(new_n246), .ZN(new_n250));
  AOI22_X1  g049(.A1(new_n250), .A2(new_n220), .B1(G183gat), .B2(G190gat), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT69), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n245), .A2(new_n254), .A3(new_n251), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n228), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  XOR2_X1   g055(.A(G113gat), .B(G120gat), .Z(new_n257));
  INV_X1    g056(.A(KEYINPUT1), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G127gat), .B(G134gat), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n262), .A2(KEYINPUT70), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT70), .B1(new_n262), .B2(new_n263), .ZN(new_n265));
  OR2_X1    g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n204), .B1(new_n256), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n228), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n245), .A2(new_n254), .A3(new_n251), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n254), .B1(new_n245), .B2(new_n251), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n266), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(KEYINPUT72), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT71), .B1(new_n271), .B2(new_n272), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n253), .A2(new_n255), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n276), .A2(new_n277), .A3(new_n266), .A4(new_n268), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n203), .B1(new_n274), .B2(new_n279), .ZN(new_n280));
  XOR2_X1   g079(.A(KEYINPUT73), .B(KEYINPUT33), .Z(new_n281));
  OAI21_X1  g080(.A(new_n202), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI22_X1  g081(.A1(new_n267), .A2(new_n273), .B1(new_n275), .B2(new_n278), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT32), .B1(new_n283), .B2(new_n203), .ZN(new_n284));
  XNOR2_X1  g083(.A(G15gat), .B(G43gat), .ZN(new_n285));
  INV_X1    g084(.A(G99gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(KEYINPUT75), .B(G71gat), .ZN(new_n288));
  XOR2_X1   g087(.A(new_n287), .B(new_n288), .Z(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n281), .ZN(new_n291));
  OAI211_X1 g090(.A(KEYINPUT74), .B(new_n291), .C1(new_n283), .C2(new_n203), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n282), .A2(new_n284), .A3(new_n290), .A4(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT34), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n283), .A2(new_n294), .A3(new_n203), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n294), .B1(new_n283), .B2(new_n203), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI221_X1 g096(.A(KEYINPUT32), .B1(new_n291), .B2(new_n289), .C1(new_n283), .C2(new_n203), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n293), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n297), .B1(new_n293), .B2(new_n298), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT36), .ZN(new_n301));
  NOR3_X1   g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n293), .A2(new_n298), .ZN(new_n303));
  INV_X1    g102(.A(new_n297), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n293), .A2(new_n297), .A3(new_n298), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT36), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(G78gat), .B(G106gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n308), .B(G22gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n309), .B(KEYINPUT86), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT76), .B(G197gat), .ZN(new_n312));
  INV_X1    g111(.A(G204gat), .ZN(new_n313));
  OR2_X1    g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT22), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT77), .B(G218gat), .ZN(new_n316));
  INV_X1    g115(.A(G211gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(new_n313), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n314), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(G211gat), .B(G218gat), .Z(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT78), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n320), .B(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT29), .ZN(new_n324));
  XOR2_X1   g123(.A(G155gat), .B(G162gat), .Z(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G141gat), .B(G148gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT80), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G155gat), .ZN(new_n330));
  INV_X1    g129(.A(G162gat), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT2), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G141gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n333), .A2(KEYINPUT80), .A3(G148gat), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n326), .A2(new_n329), .A3(new_n332), .A4(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(KEYINPUT79), .B(KEYINPUT2), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n325), .B1(new_n327), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n323), .B1(new_n324), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n320), .A2(new_n321), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(new_n324), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n320), .A2(new_n321), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n340), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n342), .B1(new_n338), .B2(new_n346), .ZN(new_n347));
  AND2_X1   g146(.A1(G228gat), .A2(G233gat), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT85), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(KEYINPUT31), .B(G50gat), .Z(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n342), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT3), .B1(new_n323), .B2(new_n324), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n354), .B(new_n348), .C1(new_n339), .C2(new_n355), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n351), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n353), .B1(new_n351), .B2(new_n356), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n311), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n351), .A2(new_n356), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(new_n352), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n351), .A2(new_n353), .A3(new_n356), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(new_n310), .A3(new_n362), .ZN(new_n363));
  AND2_X1   g162(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT37), .ZN(new_n365));
  INV_X1    g164(.A(G226gat), .ZN(new_n366));
  INV_X1    g165(.A(G233gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n368), .B(new_n268), .C1(new_n269), .C2(new_n270), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n252), .A2(new_n268), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n368), .A2(KEYINPUT29), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n323), .ZN(new_n374));
  INV_X1    g173(.A(new_n368), .ZN(new_n375));
  AOI211_X1 g174(.A(new_n375), .B(new_n228), .C1(new_n245), .C2(new_n251), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n323), .ZN(new_n378));
  INV_X1    g177(.A(new_n371), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n377), .B(new_n378), .C1(new_n256), .C2(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n365), .B1(new_n374), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G8gat), .B(G36gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(G64gat), .B(G92gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT88), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  AOI211_X1 g185(.A(new_n323), .B(new_n376), .C1(new_n271), .C2(new_n371), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n378), .B1(new_n369), .B2(new_n372), .ZN(new_n388));
  OAI21_X1  g187(.A(KEYINPUT37), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT88), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n390), .A3(new_n384), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n374), .A2(new_n380), .A3(new_n365), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n386), .A2(new_n391), .A3(KEYINPUT38), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n373), .A2(new_n378), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n377), .B1(new_n256), .B2(new_n379), .ZN(new_n395));
  OAI211_X1 g194(.A(new_n394), .B(KEYINPUT37), .C1(new_n378), .C2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n396), .A2(new_n384), .A3(new_n392), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT38), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n393), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n374), .A2(new_n380), .A3(new_n385), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT4), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n339), .B(new_n402), .C1(new_n264), .C2(new_n265), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n262), .A2(new_n263), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n338), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n403), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT82), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n338), .A2(KEYINPUT3), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n341), .A2(new_n404), .A3(new_n409), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n403), .B(KEYINPUT82), .C1(new_n402), .C2(new_n405), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n408), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G225gat), .A2(G233gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT81), .ZN(new_n414));
  OR3_X1    g213(.A1(new_n412), .A2(KEYINPUT5), .A3(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n338), .B(new_n404), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n414), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n414), .B1(new_n266), .B2(new_n339), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n418), .A2(new_n402), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n405), .B1(new_n410), .B2(KEYINPUT4), .ZN(new_n420));
  OAI211_X1 g219(.A(KEYINPUT5), .B(new_n417), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n415), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G1gat), .B(G29gat), .ZN(new_n423));
  INV_X1    g222(.A(G85gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT0), .B(G57gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  NAND2_X1  g226(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT84), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n427), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n431), .B1(new_n415), .B2(new_n421), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT84), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(KEYINPUT6), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n415), .A2(new_n431), .A3(new_n421), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n428), .A2(new_n429), .A3(new_n435), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n430), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n400), .A2(new_n401), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT30), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n401), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n374), .A2(new_n380), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n384), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n374), .A2(KEYINPUT30), .A3(new_n380), .A4(new_n385), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n440), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n445), .A2(new_n432), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n416), .A2(new_n414), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT87), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT87), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n412), .B2(new_n414), .ZN(new_n450));
  OAI211_X1 g249(.A(KEYINPUT39), .B(new_n448), .C1(new_n450), .C2(new_n447), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT39), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n412), .A2(new_n452), .A3(new_n414), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n431), .A3(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(KEYINPUT40), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n446), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n364), .B1(new_n438), .B2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT83), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n436), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n428), .A2(KEYINPUT83), .A3(new_n429), .A4(new_n435), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n459), .A2(new_n434), .A3(new_n430), .A4(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n359), .A2(new_n363), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n462), .A2(new_n463), .A3(new_n444), .ZN(new_n464));
  OAI22_X1  g263(.A1(new_n302), .A2(new_n307), .B1(new_n457), .B2(new_n464), .ZN(new_n465));
  XOR2_X1   g264(.A(KEYINPUT89), .B(KEYINPUT35), .Z(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n305), .A2(new_n306), .A3(new_n463), .A4(new_n467), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n468), .A2(new_n444), .A3(new_n437), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT35), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n299), .A2(new_n300), .A3(new_n364), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n462), .A2(new_n444), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n465), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(G8gat), .ZN(new_n475));
  OR2_X1    g274(.A1(KEYINPUT93), .A2(G1gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(KEYINPUT93), .A2(G1gat), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n476), .A2(KEYINPUT16), .A3(new_n477), .ZN(new_n478));
  XOR2_X1   g277(.A(G15gat), .B(G22gat), .Z(new_n479));
  OR2_X1    g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT94), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n475), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(G1gat), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(new_n482), .B(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT17), .ZN(new_n487));
  XNOR2_X1  g286(.A(G43gat), .B(G50gat), .ZN(new_n488));
  OR2_X1    g287(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n490));
  NAND2_X1  g289(.A1(G29gat), .A2(G36gat), .ZN(new_n491));
  OR3_X1    g290(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n489), .A2(new_n490), .A3(new_n491), .A4(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT92), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n492), .A2(KEYINPUT91), .A3(new_n493), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n497), .B(new_n491), .C1(KEYINPUT91), .C2(new_n493), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n498), .A2(KEYINPUT15), .A3(new_n488), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n486), .B1(new_n487), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n496), .A2(KEYINPUT17), .A3(new_n499), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n501), .A2(new_n502), .B1(new_n486), .B2(new_n500), .ZN(new_n503));
  NAND2_X1  g302(.A1(G229gat), .A2(G233gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n505), .B(KEYINPUT18), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n500), .B(new_n486), .ZN(new_n507));
  XOR2_X1   g306(.A(new_n504), .B(KEYINPUT13), .Z(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  XOR2_X1   g309(.A(G169gat), .B(G197gat), .Z(new_n511));
  XNOR2_X1  g310(.A(G113gat), .B(G141gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(KEYINPUT90), .B(KEYINPUT11), .Z(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  XOR2_X1   g314(.A(new_n515), .B(KEYINPUT12), .Z(new_n516));
  OR2_X1    g315(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT95), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n510), .A2(new_n516), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G57gat), .B(G64gat), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G71gat), .B(G78gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT21), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n486), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(new_n209), .ZN(new_n530));
  NAND2_X1  g329(.A1(G231gat), .A2(G233gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT96), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n530), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n526), .A2(new_n527), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(KEYINPUT97), .B(KEYINPUT19), .Z(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT98), .B(KEYINPUT20), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(G211gat), .ZN(new_n539));
  XOR2_X1   g338(.A(G127gat), .B(G155gat), .Z(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n537), .A2(new_n542), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n500), .A2(new_n487), .ZN(new_n546));
  NAND2_X1  g345(.A1(G85gat), .A2(G92gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT7), .ZN(new_n548));
  NAND2_X1  g347(.A1(G99gat), .A2(G106gat), .ZN(new_n549));
  INV_X1    g348(.A(G92gat), .ZN(new_n550));
  AOI22_X1  g349(.A1(KEYINPUT8), .A2(new_n549), .B1(new_n424), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G99gat), .B(G106gat), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n548), .B(new_n551), .C1(KEYINPUT99), .C2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(KEYINPUT99), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n553), .B(new_n554), .Z(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n546), .A2(new_n502), .A3(new_n556), .ZN(new_n557));
  AND2_X1   g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558));
  AOI22_X1  g357(.A1(new_n500), .A2(new_n555), .B1(KEYINPUT41), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G134gat), .B(G162gat), .Z(new_n561));
  XNOR2_X1  g360(.A(new_n560), .B(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(G190gat), .B(G218gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT100), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n558), .A2(KEYINPUT41), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n562), .B(new_n566), .Z(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(G230gat), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n569), .A2(new_n367), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n555), .B(new_n526), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT10), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OR3_X1    g372(.A1(new_n556), .A2(new_n526), .A3(new_n572), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n570), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n571), .A2(new_n569), .A3(new_n367), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G120gat), .B(G148gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(G176gat), .B(G204gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n577), .B(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  NOR3_X1   g381(.A1(new_n545), .A2(new_n568), .A3(new_n582), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n474), .A2(new_n521), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(new_n462), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n444), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT16), .B(G8gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n589), .B(KEYINPUT42), .Z(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(G8gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT101), .ZN(G1325gat));
  NOR2_X1   g392(.A1(new_n299), .A2(new_n300), .ZN(new_n594));
  AOI21_X1  g393(.A(G15gat), .B1(new_n584), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n301), .B1(new_n299), .B2(new_n300), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n305), .A2(KEYINPUT36), .A3(new_n306), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n584), .A2(G15gat), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n595), .B1(new_n599), .B2(new_n600), .ZN(G1326gat));
  NAND2_X1  g400(.A1(new_n584), .A2(new_n364), .ZN(new_n602));
  XNOR2_X1  g401(.A(KEYINPUT43), .B(G22gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(G1327gat));
  NAND2_X1  g403(.A1(new_n474), .A2(new_n568), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n545), .A2(new_n521), .A3(new_n581), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(G29gat), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n607), .A2(new_n608), .A3(new_n462), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT45), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT103), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n594), .A2(new_n472), .A3(new_n463), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT35), .ZN(new_n613));
  INV_X1    g412(.A(new_n437), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n471), .A2(new_n445), .A3(new_n614), .A4(new_n467), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n364), .A2(new_n461), .A3(new_n445), .ZN(new_n617));
  INV_X1    g416(.A(new_n401), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n618), .B1(new_n393), .B2(new_n399), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n619), .A2(new_n437), .B1(new_n446), .B2(new_n455), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n617), .B1(new_n620), .B2(new_n364), .ZN(new_n621));
  AND3_X1   g420(.A1(new_n598), .A2(new_n621), .A3(KEYINPUT102), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT102), .B1(new_n598), .B2(new_n621), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n616), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT44), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n624), .A2(new_n625), .A3(new_n568), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n605), .A2(KEYINPUT44), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n606), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n611), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI211_X1 g429(.A(KEYINPUT103), .B(new_n606), .C1(new_n626), .C2(new_n627), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(new_n461), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n633), .B(KEYINPUT104), .Z(new_n634));
  OAI21_X1  g433(.A(new_n610), .B1(new_n634), .B2(new_n608), .ZN(G1328gat));
  OAI21_X1  g434(.A(G36gat), .B1(new_n632), .B2(new_n445), .ZN(new_n636));
  INV_X1    g435(.A(new_n607), .ZN(new_n637));
  OR3_X1    g436(.A1(new_n637), .A2(G36gat), .A3(new_n445), .ZN(new_n638));
  AND2_X1   g437(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n639));
  NOR2_X1   g438(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI211_X1 g440(.A(new_n636), .B(new_n641), .C1(new_n639), .C2(new_n638), .ZN(G1329gat));
  NAND2_X1  g441(.A1(new_n628), .A2(new_n629), .ZN(new_n643));
  OAI21_X1  g442(.A(G43gat), .B1(new_n643), .B2(new_n598), .ZN(new_n644));
  INV_X1    g443(.A(G43gat), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n607), .A2(new_n645), .A3(new_n594), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n644), .A2(KEYINPUT47), .A3(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT106), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n625), .B1(new_n474), .B2(new_n568), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT102), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n465), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n598), .A2(new_n621), .A3(KEYINPUT102), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n567), .B1(new_n653), .B2(new_n616), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n649), .B1(new_n654), .B2(new_n625), .ZN(new_n655));
  OAI21_X1  g454(.A(KEYINPUT103), .B1(new_n655), .B2(new_n606), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n628), .A2(new_n611), .A3(new_n629), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n598), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n648), .B1(new_n658), .B2(new_n645), .ZN(new_n659));
  OAI211_X1 g458(.A(KEYINPUT106), .B(G43gat), .C1(new_n632), .C2(new_n598), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n659), .A2(new_n646), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT47), .ZN(new_n662));
  AND3_X1   g461(.A1(new_n661), .A2(KEYINPUT107), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(KEYINPUT107), .B1(new_n661), .B2(new_n662), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n647), .B1(new_n663), .B2(new_n664), .ZN(G1330gat));
  AOI21_X1  g464(.A(G50gat), .B1(new_n637), .B2(KEYINPUT110), .ZN(new_n666));
  OAI211_X1 g465(.A(new_n666), .B(new_n364), .C1(KEYINPUT110), .C2(new_n637), .ZN(new_n667));
  OAI21_X1  g466(.A(G50gat), .B1(new_n643), .B2(new_n463), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(KEYINPUT48), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(G50gat), .B1(new_n632), .B2(new_n463), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT109), .ZN(new_n671));
  OR2_X1    g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n672), .A2(new_n667), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT108), .B(KEYINPUT48), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n669), .B1(new_n674), .B2(new_n675), .ZN(G1331gat));
  INV_X1    g475(.A(new_n545), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n521), .A2(new_n581), .ZN(new_n678));
  AND4_X1   g477(.A1(new_n677), .A2(new_n624), .A3(new_n567), .A4(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n462), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT111), .B(G57gat), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(G1332gat));
  NAND2_X1  g481(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n679), .A2(new_n444), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT112), .ZN(new_n685));
  NOR2_X1   g484(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1333gat));
  AOI21_X1  g486(.A(G71gat), .B1(new_n679), .B2(new_n594), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n679), .A2(G71gat), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n688), .B1(new_n599), .B2(new_n689), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g490(.A1(new_n679), .A2(new_n364), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(G78gat), .ZN(G1335gat));
  INV_X1    g492(.A(new_n521), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n624), .A2(new_n694), .A3(new_n545), .A4(new_n568), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT51), .ZN(new_n696));
  OR2_X1    g495(.A1(new_n696), .A2(KEYINPUT113), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(KEYINPUT113), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n697), .A2(new_n424), .A3(new_n582), .A4(new_n698), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n628), .A2(new_n545), .A3(new_n678), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n700), .A2(new_n462), .ZN(new_n701));
  OAI22_X1  g500(.A1(new_n699), .A2(new_n461), .B1(new_n424), .B2(new_n701), .ZN(G1336gat));
  AOI21_X1  g501(.A(new_n550), .B1(new_n700), .B2(new_n444), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n695), .A2(KEYINPUT114), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT51), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n695), .A2(KEYINPUT114), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT115), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n709), .B(new_n710), .C1(new_n705), .C2(new_n695), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n445), .A2(G92gat), .A3(new_n581), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n703), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT52), .ZN(new_n714));
  INV_X1    g513(.A(new_n712), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n696), .B2(new_n715), .ZN(new_n716));
  OAI22_X1  g515(.A1(new_n713), .A2(new_n714), .B1(new_n703), .B2(new_n716), .ZN(G1337gat));
  NAND4_X1  g516(.A1(new_n697), .A2(new_n286), .A3(new_n582), .A4(new_n698), .ZN(new_n718));
  INV_X1    g517(.A(new_n594), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n700), .A2(new_n599), .ZN(new_n720));
  OAI22_X1  g519(.A1(new_n718), .A2(new_n719), .B1(new_n286), .B2(new_n720), .ZN(G1338gat));
  INV_X1    g520(.A(G106gat), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n722), .B1(new_n700), .B2(new_n364), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  XOR2_X1   g523(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n725));
  NOR3_X1   g524(.A1(new_n463), .A2(G106gat), .A3(new_n581), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n724), .B(new_n725), .C1(new_n696), .C2(new_n727), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n723), .B1(new_n711), .B2(new_n726), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT53), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(G1339gat));
  NOR2_X1   g530(.A1(new_n503), .A2(new_n504), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n507), .A2(new_n508), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n515), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n517), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n582), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n573), .A2(new_n574), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(new_n570), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT54), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT117), .ZN(new_n740));
  XNOR2_X1  g539(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n575), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n740), .A2(new_n580), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT55), .ZN(new_n744));
  OR3_X1    g543(.A1(new_n575), .A2(new_n576), .A3(new_n580), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n736), .B1(new_n746), .B2(new_n694), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n567), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n744), .A2(new_n745), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n749), .A2(new_n568), .A3(new_n735), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n751), .A2(new_n545), .B1(new_n694), .B2(new_n583), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n752), .A2(new_n719), .A3(new_n364), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n753), .A2(new_n462), .A3(new_n445), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n521), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G113gat), .ZN(G1340gat));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n582), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(G120gat), .ZN(G1341gat));
  NAND2_X1  g557(.A1(new_n754), .A2(new_n677), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g559(.A1(new_n754), .A2(new_n568), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(G134gat), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT56), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(G134gat), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n763), .A2(new_n764), .ZN(G1343gat));
  NOR2_X1   g564(.A1(new_n752), .A2(new_n463), .ZN(new_n766));
  OAI21_X1  g565(.A(KEYINPUT119), .B1(new_n766), .B2(KEYINPUT57), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT119), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT57), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n768), .B(new_n769), .C1(new_n752), .C2(new_n463), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n583), .A2(new_n694), .ZN(new_n771));
  INV_X1    g570(.A(new_n750), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n749), .A2(KEYINPUT120), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT120), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n521), .B1(new_n746), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n736), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n772), .B1(new_n776), .B2(new_n567), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n771), .B1(new_n777), .B2(new_n677), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n778), .A2(KEYINPUT57), .A3(new_n364), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n767), .A2(new_n770), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n599), .A2(new_n444), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n462), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(G141gat), .B1(new_n784), .B2(new_n694), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT121), .ZN(new_n786));
  INV_X1    g585(.A(new_n766), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n782), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n788), .A2(new_n333), .A3(new_n521), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n786), .A2(new_n790), .A3(KEYINPUT58), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT58), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n785), .B(new_n789), .C1(KEYINPUT121), .C2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(G1344gat));
  INV_X1    g593(.A(G148gat), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n788), .A2(new_n795), .A3(new_n582), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT59), .ZN(new_n797));
  AND2_X1   g596(.A1(new_n778), .A2(KEYINPUT122), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n364), .B1(new_n778), .B2(KEYINPUT122), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n769), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n766), .A2(KEYINPUT57), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(new_n582), .A3(new_n783), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n797), .B1(new_n803), .B2(G148gat), .ZN(new_n804));
  INV_X1    g603(.A(new_n784), .ZN(new_n805));
  AOI211_X1 g604(.A(KEYINPUT59), .B(new_n795), .C1(new_n805), .C2(new_n582), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n796), .B1(new_n804), .B2(new_n806), .ZN(G1345gat));
  AOI21_X1  g606(.A(G155gat), .B1(new_n788), .B2(new_n677), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n677), .A2(G155gat), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT123), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n808), .B1(new_n805), .B2(new_n810), .ZN(G1346gat));
  NAND3_X1  g610(.A1(new_n788), .A2(new_n331), .A3(new_n568), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT124), .ZN(new_n813));
  OAI21_X1  g612(.A(G162gat), .B1(new_n784), .B2(new_n567), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(G1347gat));
  NOR2_X1   g614(.A1(new_n462), .A2(new_n445), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n753), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n521), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n582), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g620(.A1(new_n817), .A2(new_n677), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n231), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n243), .B2(new_n822), .ZN(new_n824));
  XNOR2_X1  g623(.A(new_n824), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g624(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n826));
  XNOR2_X1  g625(.A(KEYINPUT61), .B(G190gat), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n817), .A2(new_n568), .ZN(new_n828));
  MUX2_X1   g627(.A(new_n826), .B(new_n827), .S(new_n828), .Z(G1351gat));
  NAND2_X1  g628(.A1(new_n598), .A2(new_n816), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n787), .A2(new_n830), .ZN(new_n831));
  XOR2_X1   g630(.A(KEYINPUT125), .B(G197gat), .Z(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(new_n521), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n830), .B1(new_n800), .B2(new_n801), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n834), .A2(new_n521), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n833), .B1(new_n835), .B2(new_n832), .ZN(G1352gat));
  XNOR2_X1  g635(.A(KEYINPUT126), .B(G204gat), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n831), .A2(new_n582), .A3(new_n837), .ZN(new_n838));
  XOR2_X1   g637(.A(new_n838), .B(KEYINPUT62), .Z(new_n839));
  AOI211_X1 g638(.A(new_n581), .B(new_n830), .C1(new_n800), .C2(new_n801), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n840), .B2(new_n837), .ZN(G1353gat));
  NAND3_X1  g640(.A1(new_n831), .A2(new_n317), .A3(new_n677), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT63), .ZN(new_n843));
  AOI211_X1 g642(.A(new_n843), .B(new_n317), .C1(new_n834), .C2(new_n677), .ZN(new_n844));
  INV_X1    g643(.A(new_n830), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n802), .A2(new_n677), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(KEYINPUT63), .B1(new_n846), .B2(G211gat), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n842), .B1(new_n844), .B2(new_n847), .ZN(G1354gat));
  AOI21_X1  g647(.A(G218gat), .B1(new_n831), .B2(new_n568), .ZN(new_n849));
  XOR2_X1   g648(.A(new_n849), .B(KEYINPUT127), .Z(new_n850));
  NOR2_X1   g649(.A1(new_n567), .A2(new_n316), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n850), .B1(new_n834), .B2(new_n851), .ZN(G1355gat));
endmodule


