

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732;

  XNOR2_X2 U369 ( .A(n554), .B(n553), .ZN(n731) );
  NOR2_X2 U370 ( .A1(G953), .A2(G237), .ZN(n386) );
  AND2_X1 U371 ( .A1(n504), .A2(n503), .ZN(n505) );
  XNOR2_X1 U372 ( .A(n526), .B(KEYINPUT0), .ZN(n546) );
  XNOR2_X1 U373 ( .A(n351), .B(G128), .ZN(n392) );
  XNOR2_X1 U374 ( .A(n477), .B(n476), .ZN(n691) );
  XNOR2_X1 U375 ( .A(n417), .B(n416), .ZN(n477) );
  XOR2_X2 U376 ( .A(n425), .B(n404), .Z(n717) );
  XNOR2_X2 U377 ( .A(n448), .B(n393), .ZN(n404) );
  XNOR2_X2 U378 ( .A(KEYINPUT68), .B(KEYINPUT3), .ZN(n389) );
  NOR2_X2 U379 ( .A1(n709), .A2(n566), .ZN(n548) );
  XNOR2_X2 U380 ( .A(n545), .B(KEYINPUT33), .ZN(n709) );
  XNOR2_X2 U381 ( .A(n563), .B(n478), .ZN(n569) );
  XNOR2_X1 U382 ( .A(n357), .B(n356), .ZN(n437) );
  XNOR2_X1 U383 ( .A(n392), .B(KEYINPUT4), .ZN(n448) );
  XNOR2_X1 U384 ( .A(n471), .B(n454), .ZN(n679) );
  INV_X1 U385 ( .A(KEYINPUT38), .ZN(n454) );
  XNOR2_X1 U386 ( .A(n534), .B(n533), .ZN(n572) );
  XNOR2_X1 U387 ( .A(n388), .B(KEYINPUT5), .ZN(n350) );
  XNOR2_X1 U388 ( .A(n390), .B(n389), .ZN(n438) );
  XNOR2_X1 U389 ( .A(G119), .B(G101), .ZN(n390) );
  XNOR2_X1 U390 ( .A(n365), .B(G146), .ZN(n446) );
  INV_X1 U391 ( .A(G125), .ZN(n365) );
  OR2_X1 U392 ( .A1(n679), .A2(n678), .ZN(n457) );
  XNOR2_X1 U393 ( .A(n404), .B(n347), .ZN(n593) );
  XNOR2_X1 U394 ( .A(n349), .B(n348), .ZN(n347) );
  XNOR2_X1 U395 ( .A(n387), .B(n391), .ZN(n348) );
  XNOR2_X1 U396 ( .A(n438), .B(n350), .ZN(n349) );
  INV_X1 U397 ( .A(G143), .ZN(n351) );
  XNOR2_X1 U398 ( .A(n364), .B(n363), .ZN(n367) );
  NOR2_X1 U399 ( .A1(n473), .A2(n679), .ZN(n455) );
  BUF_X1 U400 ( .A(n462), .Z(n563) );
  AND2_X1 U401 ( .A1(n477), .A2(n543), .ZN(n564) );
  BUF_X1 U402 ( .A(n546), .Z(n566) );
  NOR2_X1 U403 ( .A1(n723), .A2(G952), .ZN(n641) );
  NOR2_X1 U404 ( .A1(n710), .A2(n499), .ZN(n468) );
  XNOR2_X1 U405 ( .A(n456), .B(KEYINPUT106), .ZN(n730) );
  XNOR2_X1 U406 ( .A(n352), .B(KEYINPUT40), .ZN(n456) );
  OR2_X1 U407 ( .A1(n515), .A2(n496), .ZN(n352) );
  NOR2_X1 U408 ( .A1(n691), .A2(n490), .ZN(n663) );
  XNOR2_X1 U409 ( .A(n538), .B(n537), .ZN(n608) );
  NOR2_X1 U410 ( .A1(n572), .A2(n355), .ZN(n538) );
  XNOR2_X1 U411 ( .A(KEYINPUT103), .B(n496), .ZN(n654) );
  AND2_X1 U412 ( .A1(n517), .A2(KEYINPUT2), .ZN(n346) );
  AND2_X1 U413 ( .A1(n518), .A2(n517), .ZN(n721) );
  NAND2_X1 U414 ( .A1(n518), .A2(n346), .ZN(n520) );
  XNOR2_X1 U415 ( .A(n455), .B(KEYINPUT39), .ZN(n515) );
  BUF_X1 U416 ( .A(n610), .Z(n636) );
  XNOR2_X1 U417 ( .A(KEYINPUT24), .B(KEYINPUT92), .ZN(n353) );
  AND2_X1 U418 ( .A1(n589), .A2(n588), .ZN(G66) );
  OR2_X1 U419 ( .A1(n536), .A2(n535), .ZN(n355) );
  INV_X1 U420 ( .A(KEYINPUT86), .ZN(n541) );
  XNOR2_X1 U421 ( .A(G122), .B(G113), .ZN(n357) );
  INV_X1 U422 ( .A(KEYINPUT48), .ZN(n507) );
  XNOR2_X1 U423 ( .A(n437), .B(n360), .ZN(n364) );
  BUF_X1 U424 ( .A(n617), .Z(n667) );
  INV_X1 U425 ( .A(G469), .ZN(n414) );
  XNOR2_X1 U426 ( .A(n366), .B(G140), .ZN(n720) );
  INV_X1 U427 ( .A(KEYINPUT74), .ZN(n578) );
  XNOR2_X1 U428 ( .A(n486), .B(n485), .ZN(n497) );
  XNOR2_X1 U429 ( .A(n415), .B(n414), .ZN(n416) );
  BUF_X1 U430 ( .A(n599), .Z(n602) );
  INV_X1 U431 ( .A(KEYINPUT32), .ZN(n537) );
  XNOR2_X1 U432 ( .A(n461), .B(n460), .ZN(n710) );
  BUF_X1 U433 ( .A(n482), .Z(n471) );
  INV_X1 U434 ( .A(n641), .ZN(n588) );
  XNOR2_X1 U435 ( .A(KEYINPUT13), .B(G475), .ZN(n369) );
  INV_X1 U436 ( .A(G104), .ZN(n356) );
  XOR2_X1 U437 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n359) );
  XNOR2_X1 U438 ( .A(KEYINPUT97), .B(KEYINPUT11), .ZN(n358) );
  XNOR2_X1 U439 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U440 ( .A(G131), .B(G143), .Z(n362) );
  NAND2_X1 U441 ( .A1(G214), .A2(n386), .ZN(n361) );
  XNOR2_X1 U442 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U443 ( .A(n446), .B(KEYINPUT10), .ZN(n366) );
  XNOR2_X1 U444 ( .A(n367), .B(n720), .ZN(n611) );
  NOR2_X1 U445 ( .A1(G902), .A2(n611), .ZN(n368) );
  XNOR2_X1 U446 ( .A(n369), .B(n368), .ZN(n472) );
  INV_X1 U447 ( .A(n472), .ZN(n494) );
  INV_X2 U448 ( .A(G953), .ZN(n723) );
  NAND2_X1 U449 ( .A1(G234), .A2(n723), .ZN(n370) );
  XOR2_X1 U450 ( .A(KEYINPUT8), .B(n370), .Z(n423) );
  NAND2_X1 U451 ( .A1(n423), .A2(G217), .ZN(n373) );
  XOR2_X1 U452 ( .A(KEYINPUT99), .B(KEYINPUT9), .Z(n371) );
  XNOR2_X1 U453 ( .A(G116), .B(G107), .ZN(n440) );
  XNOR2_X1 U454 ( .A(n371), .B(n440), .ZN(n372) );
  XNOR2_X1 U455 ( .A(n373), .B(n372), .ZN(n378) );
  XOR2_X1 U456 ( .A(KEYINPUT7), .B(KEYINPUT100), .Z(n375) );
  XNOR2_X1 U457 ( .A(G134), .B(G122), .ZN(n374) );
  XNOR2_X1 U458 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U459 ( .A(n392), .B(n376), .ZN(n377) );
  XNOR2_X1 U460 ( .A(n378), .B(n377), .ZN(n633) );
  NOR2_X1 U461 ( .A1(G902), .A2(n633), .ZN(n379) );
  XOR2_X1 U462 ( .A(G478), .B(n379), .Z(n495) );
  OR2_X1 U463 ( .A1(n494), .A2(n495), .ZN(n496) );
  NAND2_X1 U464 ( .A1(G234), .A2(G237), .ZN(n380) );
  XNOR2_X1 U465 ( .A(n380), .B(KEYINPUT14), .ZN(n381) );
  XNOR2_X1 U466 ( .A(KEYINPUT72), .B(n381), .ZN(n382) );
  NAND2_X1 U467 ( .A1(G952), .A2(n382), .ZN(n708) );
  NOR2_X1 U468 ( .A1(n708), .A2(G953), .ZN(n523) );
  NAND2_X1 U469 ( .A1(G902), .A2(n382), .ZN(n521) );
  OR2_X1 U470 ( .A1(n723), .A2(n521), .ZN(n383) );
  NOR2_X1 U471 ( .A1(G900), .A2(n383), .ZN(n384) );
  NOR2_X1 U472 ( .A1(n523), .A2(n384), .ZN(n385) );
  XOR2_X1 U473 ( .A(KEYINPUT79), .B(n385), .Z(n463) );
  NAND2_X1 U474 ( .A1(n386), .A2(G210), .ZN(n388) );
  XOR2_X1 U475 ( .A(G116), .B(G146), .Z(n387) );
  XOR2_X1 U476 ( .A(G137), .B(G113), .Z(n391) );
  XNOR2_X1 U477 ( .A(G131), .B(G134), .ZN(n393) );
  INV_X1 U478 ( .A(G902), .ZN(n430) );
  NAND2_X1 U479 ( .A1(n593), .A2(n430), .ZN(n396) );
  XNOR2_X1 U480 ( .A(KEYINPUT95), .B(KEYINPUT70), .ZN(n394) );
  XNOR2_X1 U481 ( .A(n394), .B(G472), .ZN(n395) );
  XNOR2_X1 U482 ( .A(n396), .B(n395), .ZN(n462) );
  NOR2_X1 U483 ( .A1(G902), .A2(G237), .ZN(n398) );
  INV_X1 U484 ( .A(KEYINPUT73), .ZN(n397) );
  XNOR2_X1 U485 ( .A(n398), .B(n397), .ZN(n450) );
  INV_X1 U486 ( .A(G214), .ZN(n399) );
  OR2_X1 U487 ( .A1(n450), .A2(n399), .ZN(n401) );
  INV_X1 U488 ( .A(KEYINPUT90), .ZN(n400) );
  XNOR2_X1 U489 ( .A(n401), .B(n400), .ZN(n678) );
  NOR2_X1 U490 ( .A1(n462), .A2(n678), .ZN(n402) );
  XOR2_X1 U491 ( .A(KEYINPUT30), .B(n402), .Z(n403) );
  NOR2_X1 U492 ( .A1(n463), .A2(n403), .ZN(n436) );
  XOR2_X1 U493 ( .A(G137), .B(KEYINPUT66), .Z(n425) );
  XOR2_X1 U494 ( .A(G107), .B(G140), .Z(n406) );
  XNOR2_X1 U495 ( .A(G101), .B(G110), .ZN(n405) );
  XNOR2_X1 U496 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U497 ( .A(G146), .B(G104), .Z(n408) );
  NAND2_X1 U498 ( .A1(G227), .A2(n723), .ZN(n407) );
  XNOR2_X1 U499 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U500 ( .A(n410), .B(n409), .Z(n412) );
  XNOR2_X1 U501 ( .A(KEYINPUT75), .B(KEYINPUT76), .ZN(n411) );
  XNOR2_X1 U502 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U503 ( .A(n717), .B(n413), .ZN(n638) );
  NOR2_X1 U504 ( .A1(G902), .A2(n638), .ZN(n417) );
  INV_X1 U505 ( .A(KEYINPUT67), .ZN(n415) );
  XNOR2_X1 U506 ( .A(KEYINPUT15), .B(G902), .ZN(n582) );
  NAND2_X1 U507 ( .A1(G234), .A2(n582), .ZN(n418) );
  XNOR2_X1 U508 ( .A(KEYINPUT20), .B(n418), .ZN(n431) );
  NAND2_X1 U509 ( .A1(n431), .A2(G221), .ZN(n419) );
  XNOR2_X1 U510 ( .A(KEYINPUT21), .B(n419), .ZN(n687) );
  XOR2_X1 U511 ( .A(KEYINPUT94), .B(n687), .Z(n527) );
  XOR2_X1 U512 ( .A(KEYINPUT23), .B(G110), .Z(n421) );
  XNOR2_X1 U513 ( .A(G119), .B(G128), .ZN(n420) );
  XNOR2_X1 U514 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U515 ( .A(n422), .B(n720), .ZN(n429) );
  NAND2_X1 U516 ( .A1(G221), .A2(n423), .ZN(n424) );
  XNOR2_X1 U517 ( .A(n424), .B(n353), .ZN(n427) );
  XOR2_X1 U518 ( .A(n425), .B(KEYINPUT93), .Z(n426) );
  XNOR2_X1 U519 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U520 ( .A(n429), .B(n428), .ZN(n586) );
  NAND2_X1 U521 ( .A1(n586), .A2(n430), .ZN(n435) );
  NAND2_X1 U522 ( .A1(n431), .A2(G217), .ZN(n433) );
  INV_X1 U523 ( .A(KEYINPUT25), .ZN(n432) );
  XNOR2_X1 U524 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X2 U525 ( .A(n435), .B(n434), .ZN(n568) );
  NAND2_X1 U526 ( .A1(n527), .A2(n568), .ZN(n690) );
  INV_X1 U527 ( .A(n690), .ZN(n543) );
  NAND2_X1 U528 ( .A1(n436), .A2(n564), .ZN(n473) );
  XNOR2_X1 U529 ( .A(n438), .B(n437), .ZN(n442) );
  XNOR2_X1 U530 ( .A(KEYINPUT16), .B(G110), .ZN(n439) );
  XNOR2_X1 U531 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U532 ( .A(n442), .B(n441), .ZN(n627) );
  XNOR2_X1 U533 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n444) );
  NAND2_X1 U534 ( .A1(n723), .A2(G224), .ZN(n443) );
  XNOR2_X1 U535 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U536 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U537 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U538 ( .A(n627), .B(n449), .ZN(n599) );
  NAND2_X1 U539 ( .A1(n599), .A2(n582), .ZN(n453) );
  INV_X1 U540 ( .A(n450), .ZN(n451) );
  NAND2_X1 U541 ( .A1(n451), .A2(G210), .ZN(n452) );
  XNOR2_X1 U542 ( .A(n453), .B(n452), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n457), .B(KEYINPUT107), .ZN(n676) );
  NOR2_X1 U544 ( .A1(n472), .A2(n495), .ZN(n458) );
  XNOR2_X1 U545 ( .A(KEYINPUT101), .B(n458), .ZN(n681) );
  INV_X1 U546 ( .A(n681), .ZN(n459) );
  NAND2_X1 U547 ( .A1(n676), .A2(n459), .ZN(n461) );
  XOR2_X1 U548 ( .A(KEYINPUT41), .B(KEYINPUT108), .Z(n460) );
  INV_X1 U549 ( .A(n568), .ZN(n688) );
  NOR2_X1 U550 ( .A1(n687), .A2(n463), .ZN(n464) );
  NAND2_X1 U551 ( .A1(n688), .A2(n464), .ZN(n479) );
  NOR2_X1 U552 ( .A1(n563), .A2(n479), .ZN(n465) );
  XNOR2_X1 U553 ( .A(KEYINPUT28), .B(n465), .ZN(n466) );
  NAND2_X1 U554 ( .A1(n466), .A2(n477), .ZN(n499) );
  XNOR2_X1 U555 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n467) );
  XNOR2_X1 U556 ( .A(n468), .B(n467), .ZN(n732) );
  NAND2_X1 U557 ( .A1(n730), .A2(n732), .ZN(n470) );
  XOR2_X1 U558 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n469) );
  XNOR2_X1 U559 ( .A(n470), .B(n469), .ZN(n506) );
  INV_X1 U560 ( .A(n471), .ZN(n513) );
  NAND2_X1 U561 ( .A1(n472), .A2(n495), .ZN(n549) );
  NOR2_X1 U562 ( .A1(n549), .A2(n473), .ZN(n474) );
  NAND2_X1 U563 ( .A1(n513), .A2(n474), .ZN(n592) );
  NAND2_X1 U564 ( .A1(KEYINPUT47), .A2(KEYINPUT71), .ZN(n475) );
  NAND2_X1 U565 ( .A1(n592), .A2(n475), .ZN(n493) );
  INV_X1 U566 ( .A(KEYINPUT85), .ZN(n491) );
  INV_X1 U567 ( .A(KEYINPUT1), .ZN(n476) );
  INV_X1 U568 ( .A(KEYINPUT6), .ZN(n478) );
  NOR2_X1 U569 ( .A1(n569), .A2(n479), .ZN(n480) );
  XNOR2_X1 U570 ( .A(KEYINPUT104), .B(n480), .ZN(n481) );
  NAND2_X1 U571 ( .A1(n481), .A2(n654), .ZN(n509) );
  INV_X1 U572 ( .A(n509), .ZN(n487) );
  INV_X1 U573 ( .A(n482), .ZN(n484) );
  INV_X1 U574 ( .A(n678), .ZN(n483) );
  NAND2_X1 U575 ( .A1(n484), .A2(n483), .ZN(n486) );
  INV_X1 U576 ( .A(KEYINPUT88), .ZN(n485) );
  NAND2_X1 U577 ( .A1(n487), .A2(n497), .ZN(n489) );
  XOR2_X1 U578 ( .A(KEYINPUT36), .B(KEYINPUT87), .Z(n488) );
  XNOR2_X1 U579 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U580 ( .A(n491), .B(n663), .ZN(n492) );
  NOR2_X1 U581 ( .A1(n493), .A2(n492), .ZN(n504) );
  NOR2_X1 U582 ( .A1(KEYINPUT47), .A2(KEYINPUT71), .ZN(n502) );
  NAND2_X1 U583 ( .A1(n495), .A2(n494), .ZN(n659) );
  NAND2_X1 U584 ( .A1(n496), .A2(n659), .ZN(n675) );
  XNOR2_X1 U585 ( .A(n497), .B(KEYINPUT19), .ZN(n525) );
  BUF_X1 U586 ( .A(n525), .Z(n498) );
  NOR2_X1 U587 ( .A1(n499), .A2(n498), .ZN(n500) );
  XNOR2_X1 U588 ( .A(n500), .B(KEYINPUT78), .ZN(n653) );
  NAND2_X1 U589 ( .A1(n675), .A2(n653), .ZN(n501) );
  XNOR2_X1 U590 ( .A(n502), .B(n501), .ZN(n503) );
  NAND2_X1 U591 ( .A1(n506), .A2(n505), .ZN(n508) );
  XNOR2_X1 U592 ( .A(n508), .B(n507), .ZN(n518) );
  INV_X1 U593 ( .A(n691), .ZN(n544) );
  NOR2_X1 U594 ( .A1(n678), .A2(n509), .ZN(n510) );
  XNOR2_X1 U595 ( .A(n510), .B(KEYINPUT105), .ZN(n511) );
  NOR2_X1 U596 ( .A1(n544), .A2(n511), .ZN(n512) );
  XNOR2_X1 U597 ( .A(n512), .B(KEYINPUT43), .ZN(n514) );
  NOR2_X1 U598 ( .A1(n514), .A2(n513), .ZN(n591) );
  OR2_X1 U599 ( .A1(n659), .A2(n515), .ZN(n666) );
  INV_X1 U600 ( .A(n666), .ZN(n516) );
  NOR2_X1 U601 ( .A1(n591), .A2(n516), .ZN(n517) );
  INV_X1 U602 ( .A(KEYINPUT82), .ZN(n519) );
  XNOR2_X1 U603 ( .A(n520), .B(n519), .ZN(n577) );
  XNOR2_X1 U604 ( .A(G898), .B(KEYINPUT91), .ZN(n621) );
  NAND2_X1 U605 ( .A1(G953), .A2(n621), .ZN(n628) );
  NOR2_X1 U606 ( .A1(n521), .A2(n628), .ZN(n522) );
  NOR2_X1 U607 ( .A1(n523), .A2(n522), .ZN(n524) );
  OR2_X2 U608 ( .A1(n525), .A2(n524), .ZN(n526) );
  INV_X1 U609 ( .A(n546), .ZN(n531) );
  INV_X1 U610 ( .A(n527), .ZN(n528) );
  NOR2_X1 U611 ( .A1(n681), .A2(n528), .ZN(n529) );
  XNOR2_X1 U612 ( .A(n529), .B(KEYINPUT102), .ZN(n530) );
  NAND2_X1 U613 ( .A1(n531), .A2(n530), .ZN(n534) );
  INV_X1 U614 ( .A(KEYINPUT65), .ZN(n532) );
  XNOR2_X1 U615 ( .A(n532), .B(KEYINPUT22), .ZN(n533) );
  OR2_X1 U616 ( .A1(n691), .A2(n568), .ZN(n536) );
  XNOR2_X1 U617 ( .A(n569), .B(KEYINPUT77), .ZN(n535) );
  AND2_X1 U618 ( .A1(n563), .A2(n688), .ZN(n539) );
  NAND2_X1 U619 ( .A1(n691), .A2(n539), .ZN(n540) );
  OR2_X1 U620 ( .A1(n572), .A2(n540), .ZN(n590) );
  NAND2_X1 U621 ( .A1(n608), .A2(n590), .ZN(n542) );
  XNOR2_X1 U622 ( .A(n542), .B(n541), .ZN(n556) );
  NAND2_X1 U623 ( .A1(n544), .A2(n543), .ZN(n559) );
  NOR2_X1 U624 ( .A1(n569), .A2(n559), .ZN(n545) );
  XOR2_X1 U625 ( .A(KEYINPUT69), .B(KEYINPUT34), .Z(n547) );
  XNOR2_X1 U626 ( .A(n548), .B(n547), .ZN(n551) );
  INV_X1 U627 ( .A(n549), .ZN(n550) );
  NAND2_X1 U628 ( .A1(n551), .A2(n550), .ZN(n554) );
  INV_X1 U629 ( .A(KEYINPUT83), .ZN(n552) );
  XNOR2_X1 U630 ( .A(n552), .B(KEYINPUT35), .ZN(n553) );
  INV_X1 U631 ( .A(n731), .ZN(n555) );
  NAND2_X1 U632 ( .A1(n556), .A2(n555), .ZN(n558) );
  INV_X1 U633 ( .A(KEYINPUT44), .ZN(n557) );
  XNOR2_X1 U634 ( .A(n558), .B(n557), .ZN(n575) );
  INV_X1 U635 ( .A(n559), .ZN(n560) );
  INV_X1 U636 ( .A(n563), .ZN(n694) );
  NAND2_X1 U637 ( .A1(n560), .A2(n694), .ZN(n699) );
  OR2_X1 U638 ( .A1(n699), .A2(n566), .ZN(n562) );
  XOR2_X1 U639 ( .A(KEYINPUT31), .B(KEYINPUT96), .Z(n561) );
  XNOR2_X1 U640 ( .A(n562), .B(n561), .ZN(n660) );
  NAND2_X1 U641 ( .A1(n564), .A2(n563), .ZN(n565) );
  OR2_X1 U642 ( .A1(n566), .A2(n565), .ZN(n646) );
  NAND2_X1 U643 ( .A1(n660), .A2(n646), .ZN(n567) );
  NAND2_X1 U644 ( .A1(n567), .A2(n675), .ZN(n573) );
  AND2_X1 U645 ( .A1(n691), .A2(n568), .ZN(n570) );
  NAND2_X1 U646 ( .A1(n570), .A2(n569), .ZN(n571) );
  OR2_X1 U647 ( .A1(n572), .A2(n571), .ZN(n643) );
  AND2_X1 U648 ( .A1(n573), .A2(n643), .ZN(n574) );
  NAND2_X1 U649 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X2 U650 ( .A(n576), .B(KEYINPUT45), .ZN(n617) );
  NAND2_X1 U651 ( .A1(n577), .A2(n617), .ZN(n579) );
  XNOR2_X2 U652 ( .A(n579), .B(n578), .ZN(n673) );
  NAND2_X1 U653 ( .A1(n617), .A2(n721), .ZN(n581) );
  INV_X1 U654 ( .A(KEYINPUT2), .ZN(n580) );
  NAND2_X1 U655 ( .A1(n581), .A2(n580), .ZN(n584) );
  INV_X1 U656 ( .A(n582), .ZN(n583) );
  NAND2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X4 U658 ( .A1(n673), .A2(n585), .ZN(n610) );
  NAND2_X1 U659 ( .A1(n636), .A2(G217), .ZN(n587) );
  XNOR2_X1 U660 ( .A(n587), .B(n586), .ZN(n589) );
  XNOR2_X1 U661 ( .A(n590), .B(G110), .ZN(G12) );
  XOR2_X1 U662 ( .A(G140), .B(n591), .Z(G42) );
  XNOR2_X1 U663 ( .A(n592), .B(G143), .ZN(G45) );
  NAND2_X1 U664 ( .A1(n610), .A2(G472), .ZN(n595) );
  XOR2_X1 U665 ( .A(KEYINPUT62), .B(n593), .Z(n594) );
  XNOR2_X1 U666 ( .A(n595), .B(n594), .ZN(n596) );
  NOR2_X2 U667 ( .A1(n596), .A2(n641), .ZN(n598) );
  XNOR2_X1 U668 ( .A(KEYINPUT89), .B(KEYINPUT63), .ZN(n597) );
  XNOR2_X1 U669 ( .A(n598), .B(n597), .ZN(G57) );
  NAND2_X1 U670 ( .A1(n610), .A2(G210), .ZN(n604) );
  XNOR2_X1 U671 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n600) );
  XOR2_X1 U672 ( .A(n600), .B(KEYINPUT55), .Z(n601) );
  XNOR2_X1 U673 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U674 ( .A(n604), .B(n603), .ZN(n605) );
  NOR2_X2 U675 ( .A1(n605), .A2(n641), .ZN(n607) );
  XNOR2_X1 U676 ( .A(KEYINPUT84), .B(KEYINPUT56), .ZN(n606) );
  XNOR2_X1 U677 ( .A(n607), .B(n606), .ZN(G51) );
  BUF_X1 U678 ( .A(n608), .Z(n609) );
  XNOR2_X1 U679 ( .A(n609), .B(G119), .ZN(G21) );
  NAND2_X1 U680 ( .A1(n610), .A2(G475), .ZN(n613) );
  XOR2_X1 U681 ( .A(KEYINPUT59), .B(n611), .Z(n612) );
  XNOR2_X1 U682 ( .A(n613), .B(n612), .ZN(n614) );
  NOR2_X2 U683 ( .A1(n614), .A2(n641), .ZN(n616) );
  XNOR2_X1 U684 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n615) );
  XNOR2_X1 U685 ( .A(n616), .B(n615), .ZN(G60) );
  XOR2_X1 U686 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n626) );
  INV_X1 U687 ( .A(n667), .ZN(n618) );
  NOR2_X1 U688 ( .A1(n618), .A2(G953), .ZN(n623) );
  NAND2_X1 U689 ( .A1(G953), .A2(G224), .ZN(n619) );
  XOR2_X1 U690 ( .A(KEYINPUT61), .B(n619), .Z(n620) );
  NOR2_X1 U691 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U692 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U693 ( .A(n624), .B(KEYINPUT125), .ZN(n625) );
  XNOR2_X1 U694 ( .A(n626), .B(n625), .ZN(n632) );
  INV_X1 U695 ( .A(n627), .ZN(n630) );
  INV_X1 U696 ( .A(n628), .ZN(n629) );
  NOR2_X1 U697 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U698 ( .A(n632), .B(n631), .ZN(G69) );
  NAND2_X1 U699 ( .A1(n636), .A2(G478), .ZN(n634) );
  XNOR2_X1 U700 ( .A(n634), .B(n633), .ZN(n635) );
  NOR2_X1 U701 ( .A1(n635), .A2(n641), .ZN(G63) );
  NAND2_X1 U702 ( .A1(n636), .A2(G469), .ZN(n640) );
  XOR2_X1 U703 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n637) );
  XNOR2_X1 U704 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U705 ( .A(n640), .B(n639), .ZN(n642) );
  NOR2_X1 U706 ( .A1(n642), .A2(n641), .ZN(G54) );
  XNOR2_X1 U707 ( .A(G101), .B(n643), .ZN(G3) );
  INV_X1 U708 ( .A(n654), .ZN(n657) );
  NOR2_X1 U709 ( .A1(n646), .A2(n657), .ZN(n644) );
  XOR2_X1 U710 ( .A(KEYINPUT110), .B(n644), .Z(n645) );
  XNOR2_X1 U711 ( .A(G104), .B(n645), .ZN(G6) );
  NOR2_X1 U712 ( .A1(n646), .A2(n659), .ZN(n648) );
  XNOR2_X1 U713 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n647) );
  XNOR2_X1 U714 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U715 ( .A(G107), .B(n649), .ZN(G9) );
  XOR2_X1 U716 ( .A(G128), .B(KEYINPUT29), .Z(n652) );
  INV_X1 U717 ( .A(n659), .ZN(n650) );
  NAND2_X1 U718 ( .A1(n650), .A2(n653), .ZN(n651) );
  XNOR2_X1 U719 ( .A(n652), .B(n651), .ZN(G30) );
  XOR2_X1 U720 ( .A(G146), .B(KEYINPUT111), .Z(n656) );
  NAND2_X1 U721 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U722 ( .A(n656), .B(n655), .ZN(G48) );
  NOR2_X1 U723 ( .A1(n660), .A2(n657), .ZN(n658) );
  XOR2_X1 U724 ( .A(G113), .B(n658), .Z(G15) );
  NOR2_X1 U725 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U726 ( .A(KEYINPUT112), .B(n661), .Z(n662) );
  XNOR2_X1 U727 ( .A(G116), .B(n662), .ZN(G18) );
  XNOR2_X1 U728 ( .A(G125), .B(n663), .ZN(n664) );
  XNOR2_X1 U729 ( .A(n664), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U730 ( .A(G134), .B(KEYINPUT113), .Z(n665) );
  XNOR2_X1 U731 ( .A(n666), .B(n665), .ZN(G36) );
  XOR2_X1 U732 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n716) );
  XNOR2_X1 U733 ( .A(KEYINPUT2), .B(KEYINPUT80), .ZN(n668) );
  OR2_X1 U734 ( .A1(n667), .A2(n668), .ZN(n671) );
  NOR2_X1 U735 ( .A1(n721), .A2(n668), .ZN(n669) );
  XNOR2_X1 U736 ( .A(KEYINPUT81), .B(n669), .ZN(n670) );
  NAND2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  NOR2_X1 U738 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U739 ( .A1(G953), .A2(n674), .ZN(n714) );
  NAND2_X1 U740 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U741 ( .A(KEYINPUT117), .B(n677), .ZN(n683) );
  AND2_X1 U742 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U743 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U744 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U745 ( .A(n684), .B(KEYINPUT118), .ZN(n685) );
  NOR2_X1 U746 ( .A1(n709), .A2(n685), .ZN(n686) );
  XOR2_X1 U747 ( .A(KEYINPUT119), .B(n686), .Z(n705) );
  AND2_X1 U748 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U749 ( .A(KEYINPUT49), .B(n689), .ZN(n697) );
  XOR2_X1 U750 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n693) );
  NAND2_X1 U751 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U752 ( .A(n693), .B(n692), .ZN(n695) );
  NOR2_X1 U753 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X1 U754 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U755 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U756 ( .A(n700), .B(KEYINPUT51), .Z(n701) );
  XNOR2_X1 U757 ( .A(KEYINPUT115), .B(n701), .ZN(n702) );
  NOR2_X1 U758 ( .A1(n710), .A2(n702), .ZN(n703) );
  XNOR2_X1 U759 ( .A(KEYINPUT116), .B(n703), .ZN(n704) );
  NOR2_X1 U760 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U761 ( .A(n706), .B(KEYINPUT52), .ZN(n707) );
  NOR2_X1 U762 ( .A1(n708), .A2(n707), .ZN(n712) );
  NOR2_X1 U763 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U764 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U765 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U766 ( .A(n716), .B(n715), .ZN(G75) );
  XNOR2_X1 U767 ( .A(KEYINPUT127), .B(KEYINPUT126), .ZN(n718) );
  XNOR2_X1 U768 ( .A(n718), .B(n717), .ZN(n719) );
  XNOR2_X1 U769 ( .A(n720), .B(n719), .ZN(n725) );
  INV_X1 U770 ( .A(n725), .ZN(n722) );
  XNOR2_X1 U771 ( .A(n722), .B(n721), .ZN(n724) );
  NAND2_X1 U772 ( .A1(n724), .A2(n723), .ZN(n729) );
  XNOR2_X1 U773 ( .A(G227), .B(n725), .ZN(n726) );
  NAND2_X1 U774 ( .A1(n726), .A2(G900), .ZN(n727) );
  NAND2_X1 U775 ( .A1(n727), .A2(G953), .ZN(n728) );
  NAND2_X1 U776 ( .A1(n729), .A2(n728), .ZN(G72) );
  XNOR2_X1 U777 ( .A(G131), .B(n730), .ZN(G33) );
  XOR2_X1 U778 ( .A(G122), .B(n731), .Z(G24) );
  XNOR2_X1 U779 ( .A(G137), .B(n732), .ZN(G39) );
endmodule

