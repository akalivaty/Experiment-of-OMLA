//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 0 0 1 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n604, new_n605, new_n606, new_n607, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934;
  INV_X1    g000(.A(KEYINPUT67), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT2), .ZN(new_n188));
  INV_X1    g002(.A(G113), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n187), .A2(new_n188), .A3(new_n189), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n191));
  AOI22_X1  g005(.A1(new_n190), .A2(new_n191), .B1(KEYINPUT2), .B2(G113), .ZN(new_n192));
  XNOR2_X1  g006(.A(G116), .B(G119), .ZN(new_n193));
  OR2_X1    g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n190), .A2(new_n191), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT2), .A2(G113), .ZN(new_n196));
  AND4_X1   g010(.A1(KEYINPUT68), .A2(new_n195), .A3(new_n196), .A4(new_n193), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT68), .B1(new_n192), .B2(new_n193), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n194), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(new_n200), .A3(G143), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n202), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  AND2_X1   g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(KEYINPUT0), .A2(G128), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n201), .A2(new_n204), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n207), .A2(new_n210), .B1(new_n212), .B2(new_n208), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT69), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT11), .A2(G134), .ZN(new_n216));
  NOR2_X1   g030(.A1(KEYINPUT11), .A2(G134), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n216), .B1(new_n217), .B2(G137), .ZN(new_n218));
  INV_X1    g032(.A(G131), .ZN(new_n219));
  XNOR2_X1  g033(.A(KEYINPUT66), .B(G137), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n218), .B(new_n219), .C1(new_n220), .C2(new_n216), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(KEYINPUT11), .A2(G134), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n224), .A2(G137), .ZN(new_n225));
  INV_X1    g039(.A(G137), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(KEYINPUT66), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n223), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n219), .B1(new_n228), .B2(new_n218), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n215), .B1(new_n222), .B2(new_n229), .ZN(new_n230));
  OR2_X1    g044(.A1(KEYINPUT11), .A2(G134), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n223), .B1(new_n231), .B2(new_n226), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n226), .A2(KEYINPUT66), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n224), .A2(G137), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n216), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(G131), .B1(new_n232), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT69), .A3(new_n221), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n214), .B1(new_n230), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G128), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n207), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT1), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n212), .A2(new_n242), .A3(G128), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(G134), .A2(G137), .ZN(new_n245));
  OAI211_X1 g059(.A(G131), .B(new_n245), .C1(new_n220), .C2(G134), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n244), .A2(new_n221), .A3(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n199), .B1(new_n238), .B2(new_n247), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n236), .A2(KEYINPUT69), .A3(new_n221), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT69), .B1(new_n236), .B2(new_n221), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n213), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n199), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n244), .A2(new_n221), .A3(new_n246), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n248), .A2(KEYINPUT73), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT73), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n251), .A2(new_n256), .A3(new_n252), .A4(new_n253), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n255), .A2(KEYINPUT28), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n259));
  NOR3_X1   g073(.A1(new_n238), .A2(new_n199), .A3(new_n247), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n259), .B1(new_n260), .B2(KEYINPUT28), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n254), .A2(KEYINPUT71), .A3(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n264));
  INV_X1    g078(.A(G237), .ZN(new_n265));
  INV_X1    g079(.A(G953), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n266), .A3(G210), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n264), .B(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT26), .B(G101), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n271), .A2(KEYINPUT29), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n258), .A2(new_n261), .A3(new_n263), .A4(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G902), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT74), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n273), .A2(KEYINPUT74), .A3(new_n274), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n251), .A2(KEYINPUT30), .A3(new_n253), .ZN(new_n279));
  XNOR2_X1  g093(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n213), .B1(new_n222), .B2(new_n229), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n280), .B1(new_n247), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n279), .A2(new_n283), .A3(new_n199), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n254), .ZN(new_n285));
  AOI21_X1  g099(.A(KEYINPUT29), .B1(new_n285), .B2(new_n270), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n252), .B1(new_n281), .B2(new_n253), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT28), .B1(new_n260), .B2(new_n287), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n261), .A2(new_n288), .A3(new_n263), .A4(new_n271), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT72), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n286), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n277), .A2(new_n278), .A3(new_n291), .A4(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G472), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT75), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n284), .A2(new_n254), .A3(new_n271), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT31), .ZN(new_n298));
  OR2_X1    g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n298), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n261), .A2(new_n288), .A3(new_n263), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n270), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT32), .ZN(new_n305));
  NOR2_X1   g119(.A1(G472), .A2(G902), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n299), .A2(new_n300), .B1(new_n302), .B2(new_n270), .ZN(new_n308));
  INV_X1    g122(.A(new_n306), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT32), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT75), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n294), .A2(new_n312), .A3(G472), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n296), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(G110), .B(G122), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT4), .ZN(new_n317));
  INV_X1    g131(.A(G104), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT3), .B1(new_n318), .B2(G107), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n320));
  INV_X1    g134(.A(G107), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G104), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n318), .A2(G107), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n319), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT79), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(G101), .ZN(new_n326));
  INV_X1    g140(.A(G101), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n319), .A2(new_n322), .A3(new_n327), .A4(new_n323), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n317), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n326), .A2(new_n317), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n195), .A2(new_n196), .A3(new_n193), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT68), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n192), .A2(KEYINPUT68), .A3(new_n193), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI22_X1  g150(.A1(new_n330), .A2(new_n331), .B1(new_n336), .B2(new_n194), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n197), .A2(new_n198), .ZN(new_n338));
  INV_X1    g152(.A(G119), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G116), .ZN(new_n340));
  INV_X1    g154(.A(G116), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G119), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n342), .A3(KEYINPUT5), .ZN(new_n343));
  OR3_X1    g157(.A1(new_n341), .A2(KEYINPUT5), .A3(G119), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(G113), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT86), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n343), .A2(new_n344), .A3(KEYINPUT86), .A4(G113), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n323), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n318), .A2(G107), .ZN(new_n351));
  OAI21_X1  g165(.A(G101), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n328), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n338), .A2(new_n349), .A3(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n316), .B1(new_n337), .B2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n349), .ZN(new_n356));
  INV_X1    g170(.A(new_n353), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n336), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n331), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n199), .B1(new_n329), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n358), .A2(new_n360), .A3(new_n315), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n355), .A2(KEYINPUT6), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT6), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n363), .B(new_n316), .C1(new_n337), .C2(new_n354), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n244), .A2(G125), .ZN(new_n365));
  INV_X1    g179(.A(G125), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n213), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(G224), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n369), .A2(G953), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n368), .B(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n362), .A2(new_n364), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(KEYINPUT7), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n374), .B1(new_n367), .B2(KEYINPUT88), .ZN(new_n375));
  OR2_X1    g189(.A1(new_n368), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n315), .B(KEYINPUT87), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(KEYINPUT8), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n357), .B1(new_n356), .B2(new_n336), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n336), .A2(new_n357), .A3(new_n345), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n368), .A2(new_n375), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n376), .A2(new_n381), .A3(new_n361), .A4(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n373), .A2(new_n274), .A3(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(G210), .B1(G237), .B2(G902), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n373), .A2(new_n274), .A3(new_n385), .A4(new_n383), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(G214), .B1(G237), .B2(G902), .ZN(new_n391));
  XOR2_X1   g205(.A(new_n391), .B(KEYINPUT85), .Z(new_n392));
  NOR2_X1   g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  OAI211_X1 g207(.A(KEYINPUT80), .B(KEYINPUT1), .C1(new_n203), .C2(G146), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G128), .ZN(new_n395));
  AOI21_X1  g209(.A(KEYINPUT80), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n211), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT81), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI211_X1 g213(.A(KEYINPUT81), .B(new_n211), .C1(new_n395), .C2(new_n396), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n243), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n357), .ZN(new_n402));
  XOR2_X1   g216(.A(KEYINPUT82), .B(KEYINPUT10), .Z(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n213), .B1(new_n359), .B2(new_n329), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n244), .A2(KEYINPUT10), .A3(new_n357), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n249), .A2(new_n250), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n407), .A2(new_n409), .ZN(new_n411));
  XNOR2_X1  g225(.A(G110), .B(G140), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n266), .A2(G227), .ZN(new_n413));
  XOR2_X1   g227(.A(new_n412), .B(new_n413), .Z(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NOR3_X1   g229(.A1(new_n410), .A2(new_n411), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT12), .ZN(new_n418));
  AND3_X1   g232(.A1(new_n241), .A2(new_n353), .A3(new_n243), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n419), .B1(new_n401), .B2(new_n357), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n418), .B1(new_n420), .B2(new_n408), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT83), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n222), .A2(new_n229), .ZN(new_n424));
  OR3_X1    g238(.A1(new_n420), .A2(new_n418), .A3(new_n424), .ZN(new_n425));
  OAI211_X1 g239(.A(KEYINPUT83), .B(new_n418), .C1(new_n420), .C2(new_n408), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n423), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  OR2_X1    g241(.A1(new_n407), .A2(new_n409), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n415), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT84), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n417), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n414), .B1(new_n427), .B2(new_n428), .ZN(new_n433));
  OAI21_X1  g247(.A(KEYINPUT84), .B1(new_n433), .B2(new_n416), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n432), .A2(G469), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(G469), .A2(G902), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n427), .A2(new_n428), .A3(new_n414), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n415), .B1(new_n410), .B2(new_n411), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(G469), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(new_n274), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n435), .A2(new_n436), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G128), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(G143), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(G143), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(G134), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n447), .B(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G122), .ZN(new_n450));
  OAI21_X1  g264(.A(KEYINPUT14), .B1(new_n450), .B2(G116), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT92), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(G116), .ZN(new_n454));
  OR3_X1    g268(.A1(new_n450), .A2(KEYINPUT14), .A3(G116), .ZN(new_n455));
  OAI211_X1 g269(.A(KEYINPUT92), .B(KEYINPUT14), .C1(new_n450), .C2(G116), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n453), .A2(new_n454), .A3(new_n455), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G107), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT93), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G116), .B(G122), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n321), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n457), .A2(KEYINPUT93), .A3(G107), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n449), .A2(new_n460), .A3(new_n462), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n447), .A2(new_n448), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n461), .B(new_n321), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT91), .ZN(new_n467));
  OR3_X1    g281(.A1(new_n444), .A2(new_n467), .A3(KEYINPUT13), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n444), .A2(KEYINPUT13), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n467), .B1(new_n444), .B2(KEYINPUT13), .ZN(new_n470));
  AND4_X1   g284(.A1(new_n446), .A2(new_n468), .A3(new_n469), .A4(new_n470), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n465), .B(new_n466), .C1(new_n471), .C2(new_n448), .ZN(new_n472));
  XOR2_X1   g286(.A(KEYINPUT9), .B(G234), .Z(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(G217), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n474), .A2(new_n475), .A3(G953), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n464), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n476), .B1(new_n464), .B2(new_n472), .ZN(new_n478));
  OR2_X1    g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n274), .ZN(new_n480));
  INV_X1    g294(.A(G478), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT94), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(KEYINPUT15), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(KEYINPUT15), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n481), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n486), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n479), .A2(new_n274), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(G475), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n366), .A2(KEYINPUT16), .A3(G140), .ZN(new_n492));
  XNOR2_X1  g306(.A(G125), .B(G140), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n492), .B1(new_n493), .B2(KEYINPUT16), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(G146), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n494), .A2(G146), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n265), .A2(new_n266), .A3(G214), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(new_n203), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n500), .A2(KEYINPUT17), .A3(G131), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(G131), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n499), .B(G143), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n219), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n498), .B(new_n501), .C1(new_n505), .C2(KEYINPUT17), .ZN(new_n506));
  NAND2_X1  g320(.A1(KEYINPUT18), .A2(G131), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n500), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n493), .B(G146), .ZN(new_n509));
  OR2_X1    g323(.A1(new_n509), .A2(KEYINPUT89), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(KEYINPUT89), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n508), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(G113), .B(G122), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(new_n318), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n506), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n493), .A2(KEYINPUT90), .ZN(new_n517));
  XOR2_X1   g331(.A(new_n517), .B(KEYINPUT19), .Z(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n200), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n496), .B1(new_n502), .B2(new_n504), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n514), .B1(new_n521), .B2(new_n512), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n491), .B(new_n274), .C1(new_n516), .C2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT20), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n521), .A2(new_n512), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n515), .B1(new_n526), .B2(new_n514), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n527), .A2(KEYINPUT20), .A3(new_n491), .A4(new_n274), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n514), .B1(new_n506), .B2(new_n512), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n274), .B1(new_n516), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(G475), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n525), .A2(new_n528), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(G234), .A2(G237), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(G952), .A3(new_n266), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  XOR2_X1   g349(.A(KEYINPUT21), .B(G898), .Z(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n533), .A2(G902), .A3(G953), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n535), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n490), .A2(new_n532), .A3(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(G221), .B1(new_n474), .B2(G902), .ZN(new_n542));
  AND4_X1   g356(.A1(new_n393), .A2(new_n442), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n266), .A2(G221), .A3(G234), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(G137), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT78), .B(KEYINPUT22), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n443), .A2(G119), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(KEYINPUT76), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT23), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n339), .A2(G128), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT23), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n548), .A2(KEYINPUT76), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n550), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n551), .A2(new_n548), .ZN(new_n555));
  XOR2_X1   g369(.A(KEYINPUT24), .B(G110), .Z(new_n556));
  OAI22_X1  g370(.A1(new_n554), .A2(G110), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n493), .A2(new_n200), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(new_n495), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT77), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n554), .A2(G110), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n555), .A2(new_n556), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n561), .B(new_n562), .C1(new_n496), .C2(new_n497), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n559), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n560), .B1(new_n559), .B2(new_n563), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n547), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n547), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n559), .A3(new_n563), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT25), .B1(new_n569), .B2(G902), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n475), .B1(G234), .B2(new_n274), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT25), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n566), .A2(new_n572), .A3(new_n274), .A4(new_n568), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n571), .A2(G902), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n566), .A2(new_n568), .A3(new_n575), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n314), .A2(new_n543), .A3(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(G101), .ZN(G3));
  AND2_X1   g393(.A1(new_n442), .A2(new_n542), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n304), .A2(new_n274), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(G472), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n304), .A2(new_n306), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n580), .A2(new_n577), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n479), .A2(KEYINPUT33), .ZN(new_n587));
  OR3_X1    g401(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT33), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(G478), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(G478), .A2(G902), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n479), .A2(new_n481), .A3(new_n274), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n532), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n387), .A2(KEYINPUT95), .A3(new_n388), .ZN(new_n595));
  INV_X1    g409(.A(new_n392), .ZN(new_n596));
  OR2_X1    g410(.A1(new_n388), .A2(KEYINPUT95), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n540), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR3_X1   g414(.A1(new_n586), .A2(new_n594), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT34), .B(G104), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G6));
  NAND4_X1  g417(.A1(new_n490), .A2(new_n531), .A3(new_n525), .A4(new_n528), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n586), .A2(new_n600), .A3(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G107), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT96), .B(KEYINPUT35), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n606), .B(new_n607), .ZN(G9));
  OR2_X1    g422(.A1(new_n564), .A2(new_n565), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n547), .A2(KEYINPUT36), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(new_n575), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n574), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n543), .A2(new_n585), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G110), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT97), .B(KEYINPUT37), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G12));
  AND3_X1   g431(.A1(new_n442), .A2(new_n542), .A3(new_n598), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT98), .B(G900), .Z(new_n619));
  AOI21_X1  g433(.A(new_n535), .B1(new_n619), .B2(new_n539), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n604), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n314), .A2(new_n613), .A3(new_n618), .A4(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G128), .ZN(G30));
  INV_X1    g437(.A(new_n613), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n490), .A2(new_n532), .A3(new_n596), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT38), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n389), .B(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n626), .A2(new_n627), .ZN(new_n632));
  INV_X1    g446(.A(G472), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n255), .A2(new_n270), .A3(new_n257), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT99), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(G902), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n634), .A2(new_n635), .A3(new_n297), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n633), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(KEYINPUT100), .B1(new_n311), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n642));
  AOI211_X1 g456(.A(new_n642), .B(new_n639), .C1(new_n307), .C2(new_n310), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n631), .B(new_n632), .C1(new_n641), .C2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OR2_X1    g460(.A1(new_n641), .A2(new_n643), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n647), .A2(KEYINPUT102), .A3(new_n631), .A4(new_n632), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n620), .B(KEYINPUT39), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n580), .A2(KEYINPUT40), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n580), .A2(new_n650), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT40), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI22_X1  g468(.A1(new_n646), .A2(new_n648), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(new_n203), .ZN(G45));
  NOR2_X1   g470(.A1(new_n594), .A2(new_n620), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n314), .A2(new_n613), .A3(new_n618), .A4(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G146), .ZN(G48));
  NOR2_X1   g473(.A1(new_n600), .A2(new_n594), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n440), .B1(new_n439), .B2(new_n274), .ZN(new_n661));
  AOI211_X1 g475(.A(G469), .B(G902), .C1(new_n437), .C2(new_n438), .ZN(new_n662));
  INV_X1    g476(.A(new_n542), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT103), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n439), .A2(new_n274), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G469), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n668), .A2(new_n542), .A3(new_n441), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT103), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n314), .A2(new_n660), .A3(new_n577), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT41), .B(G113), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G15));
  NOR2_X1   g488(.A1(new_n600), .A2(new_n604), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n314), .A2(new_n577), .A3(new_n675), .A4(new_n671), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G116), .ZN(G18));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n678), .B1(new_n669), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n664), .A2(new_n598), .A3(KEYINPUT104), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n314), .A2(new_n682), .A3(new_n541), .A4(new_n613), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G119), .ZN(G21));
  NAND3_X1  g498(.A1(new_n625), .A2(new_n597), .A3(new_n595), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n540), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT105), .B(G472), .Z(new_n687));
  NAND2_X1  g501(.A1(new_n581), .A2(new_n687), .ZN(new_n688));
  AND3_X1   g502(.A1(new_n258), .A2(new_n261), .A3(new_n263), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n301), .B1(new_n689), .B2(new_n271), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n306), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n671), .A2(new_n686), .A3(new_n577), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G122), .ZN(G24));
  AND3_X1   g508(.A1(new_n688), .A2(new_n613), .A3(new_n691), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n682), .A2(new_n657), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G125), .ZN(G27));
  NAND2_X1  g511(.A1(new_n430), .A2(KEYINPUT107), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n433), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n698), .A2(G469), .A3(new_n417), .A4(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n436), .B(KEYINPUT106), .Z(new_n702));
  NAND3_X1  g516(.A1(new_n701), .A2(new_n441), .A3(new_n702), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n389), .A2(new_n392), .A3(new_n663), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n657), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n314), .A2(new_n577), .A3(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT42), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n314), .A2(KEYINPUT42), .A3(new_n577), .A4(new_n705), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G131), .ZN(G33));
  AND3_X1   g525(.A1(new_n314), .A2(new_n577), .A3(new_n621), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n703), .A2(new_n704), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G134), .ZN(G36));
  NAND4_X1  g529(.A1(new_n698), .A2(KEYINPUT45), .A3(new_n417), .A4(new_n700), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(G469), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT45), .B1(new_n432), .B2(new_n434), .ZN(new_n718));
  OAI211_X1 g532(.A(KEYINPUT46), .B(new_n702), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(KEYINPUT108), .A3(new_n441), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT108), .B1(new_n719), .B2(new_n441), .ZN(new_n722));
  OR2_X1    g536(.A1(new_n717), .A2(new_n718), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT46), .B1(new_n723), .B2(new_n702), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n725), .A2(new_n663), .A3(new_n649), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n592), .A2(new_n532), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT43), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n584), .A3(new_n613), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g545(.A(new_n731), .B(KEYINPUT109), .Z(new_n732));
  NAND2_X1  g546(.A1(new_n390), .A2(new_n596), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n729), .A2(new_n730), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n726), .A2(new_n732), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  XOR2_X1   g550(.A(KEYINPUT110), .B(G137), .Z(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G39));
  INV_X1    g552(.A(KEYINPUT47), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n739), .B1(new_n725), .B2(new_n663), .ZN(new_n740));
  INV_X1    g554(.A(new_n722), .ZN(new_n741));
  INV_X1    g555(.A(new_n724), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n742), .A3(new_n720), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(KEYINPUT47), .A3(new_n542), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  NOR4_X1   g559(.A1(new_n314), .A2(new_n577), .A3(new_n594), .A4(new_n620), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n734), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G140), .ZN(G42));
  INV_X1    g562(.A(G952), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n266), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT53), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n701), .A2(new_n702), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n685), .B1(new_n752), .B2(new_n441), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n613), .A2(new_n663), .A3(new_n620), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n753), .B(new_n754), .C1(new_n641), .C2(new_n643), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n622), .A2(new_n658), .A3(new_n696), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(KEYINPUT52), .ZN(new_n757));
  AOI22_X1  g571(.A1(new_n708), .A2(new_n709), .B1(new_n712), .B2(new_n713), .ZN(new_n758));
  AND4_X1   g572(.A1(new_n672), .A2(new_n683), .A3(new_n676), .A4(new_n693), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n490), .A2(new_n532), .A3(new_n620), .ZN(new_n760));
  AND3_X1   g574(.A1(new_n442), .A2(new_n542), .A3(new_n760), .ZN(new_n761));
  AND3_X1   g575(.A1(new_n314), .A2(new_n734), .A3(new_n761), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n705), .A2(new_n692), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n613), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n594), .A2(new_n604), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n765), .A2(new_n393), .A3(new_n599), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(new_n580), .A3(new_n577), .A4(new_n585), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n578), .A2(new_n614), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n758), .A2(new_n759), .A3(new_n764), .A4(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n751), .B1(new_n757), .B2(new_n770), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n294), .A2(new_n312), .A3(G472), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n312), .B1(new_n294), .B2(G472), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n624), .B1(new_n774), .B2(new_n311), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n775), .B(new_n618), .C1(new_n621), .C2(new_n657), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n776), .A2(KEYINPUT52), .A3(new_n696), .A4(new_n755), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n756), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n764), .A2(new_n710), .A3(new_n714), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n683), .A2(new_n672), .A3(new_n676), .A4(new_n693), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n768), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n780), .A2(new_n781), .A3(KEYINPUT53), .A4(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n771), .A2(KEYINPUT112), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT112), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n787), .B(new_n751), .C1(new_n757), .C2(new_n770), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n785), .A2(new_n786), .A3(KEYINPUT54), .A4(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n771), .A2(new_n790), .A3(new_n784), .ZN(new_n791));
  OAI211_X1 g605(.A(KEYINPUT114), .B(new_n751), .C1(new_n757), .C2(new_n770), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT113), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n785), .A2(KEYINPUT54), .A3(new_n788), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n789), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AND4_X1   g611(.A1(new_n577), .A2(new_n692), .A3(new_n728), .A4(new_n535), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n661), .A2(new_n662), .A3(new_n542), .ZN(new_n799));
  OAI211_X1 g613(.A(new_n734), .B(new_n798), .C1(new_n745), .C2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n647), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n669), .A2(new_n733), .A3(new_n534), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n577), .A3(new_n802), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n803), .A2(new_n532), .A3(new_n593), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n728), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT115), .Z(new_n806));
  INV_X1    g620(.A(KEYINPUT116), .ZN(new_n807));
  INV_X1    g621(.A(new_n695), .ZN(new_n808));
  OR3_X1    g622(.A1(new_n806), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n807), .B1(new_n806), .B2(new_n808), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n804), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n798), .A2(new_n392), .A3(new_n630), .A4(new_n664), .ZN(new_n812));
  XOR2_X1   g626(.A(new_n812), .B(KEYINPUT50), .Z(new_n813));
  NAND3_X1  g627(.A1(new_n800), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n803), .A2(new_n594), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n814), .A2(new_n815), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n314), .A2(new_n577), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n806), .A2(new_n819), .ZN(new_n820));
  OR2_X1    g634(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n820), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  AOI211_X1 g638(.A(new_n749), .B(G953), .C1(new_n798), .C2(new_n682), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n816), .A2(new_n817), .A3(new_n818), .A4(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n750), .B1(new_n797), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n661), .A2(new_n662), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT49), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n630), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT111), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n577), .A2(new_n596), .A3(new_n542), .ZN(new_n834));
  AOI211_X1 g648(.A(new_n831), .B(new_n832), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n727), .B1(new_n834), .B2(new_n833), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n830), .B2(new_n829), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n801), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n828), .A2(new_n838), .ZN(G75));
  NAND4_X1  g653(.A1(new_n791), .A2(G210), .A3(G902), .A4(new_n792), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT56), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n362), .A2(new_n364), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(new_n372), .ZN(new_n843));
  XNOR2_X1  g657(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n844));
  XOR2_X1   g658(.A(new_n843), .B(new_n844), .Z(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n840), .A2(new_n841), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n846), .B1(new_n840), .B2(new_n841), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n266), .A2(G952), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(G51));
  XOR2_X1   g664(.A(new_n702), .B(KEYINPUT57), .Z(new_n851));
  NOR2_X1   g665(.A1(new_n793), .A2(new_n794), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT54), .B1(new_n791), .B2(new_n792), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n439), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n723), .B(KEYINPUT119), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n791), .A2(G902), .A3(new_n792), .A4(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n849), .B1(new_n855), .B2(new_n857), .ZN(G54));
  INV_X1    g672(.A(KEYINPUT120), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n859), .A2(KEYINPUT58), .A3(G475), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n791), .A2(G902), .A3(new_n792), .A4(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n527), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n859), .B1(KEYINPUT58), .B2(G475), .ZN(new_n863));
  OR3_X1    g677(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n849), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n862), .B1(new_n861), .B2(new_n863), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(G60));
  AND2_X1   g681(.A1(new_n587), .A2(new_n588), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n590), .B(KEYINPUT59), .Z(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(new_n852), .B2(new_n853), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n865), .ZN(new_n872));
  INV_X1    g686(.A(new_n869), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n797), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n872), .B1(new_n874), .B2(new_n868), .ZN(G63));
  NAND2_X1  g689(.A1(G217), .A2(G902), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n876), .B(KEYINPUT60), .Z(new_n877));
  NAND3_X1  g691(.A1(new_n791), .A2(new_n792), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(new_n569), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n791), .A2(new_n611), .A3(new_n792), .A4(new_n877), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n879), .A2(new_n865), .A3(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n881), .A2(new_n882), .A3(KEYINPUT61), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT61), .B1(new_n881), .B2(new_n882), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(G66));
  OAI21_X1  g699(.A(G953), .B1(new_n537), .B2(new_n369), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n886), .B1(new_n783), .B2(G953), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT122), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n842), .B1(G898), .B2(new_n266), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n888), .B(new_n889), .ZN(G69));
  AND2_X1   g704(.A1(new_n747), .A2(new_n736), .ZN(new_n891));
  INV_X1    g705(.A(new_n758), .ZN(new_n892));
  INV_X1    g706(.A(new_n819), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n743), .A2(new_n893), .A3(new_n542), .A4(new_n650), .ZN(new_n894));
  OR3_X1    g708(.A1(new_n894), .A2(KEYINPUT125), .A3(new_n685), .ZN(new_n895));
  OAI21_X1  g709(.A(KEYINPUT125), .B1(new_n894), .B2(new_n685), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n892), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n622), .A2(new_n658), .A3(new_n696), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n891), .A2(new_n897), .A3(new_n266), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n279), .A2(new_n283), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n518), .B(KEYINPUT123), .Z(new_n901));
  XNOR2_X1  g715(.A(new_n900), .B(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(G900), .A2(G953), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n899), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n646), .A2(new_n648), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n654), .A2(new_n651), .ZN(new_n907));
  OAI211_X1 g721(.A(KEYINPUT62), .B(new_n898), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT62), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n776), .A2(new_n696), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n909), .B1(new_n655), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n652), .A2(new_n733), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n893), .A2(new_n913), .A3(new_n765), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n912), .A2(new_n747), .A3(new_n736), .A4(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(new_n266), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT124), .B1(new_n916), .B2(new_n902), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT126), .B1(new_n905), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(G227), .B1(new_n903), .B2(KEYINPUT126), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n266), .B1(new_n920), .B2(G900), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n918), .B(new_n921), .ZN(G72));
  XNOR2_X1  g736(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n633), .A2(new_n274), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n783), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n925), .B1(new_n915), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n927), .A2(new_n271), .A3(new_n285), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n285), .A2(new_n270), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n297), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n785), .A2(new_n788), .A3(new_n925), .A4(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n891), .A2(new_n897), .A3(new_n783), .A4(new_n898), .ZN(new_n933));
  AOI211_X1 g747(.A(new_n271), .B(new_n285), .C1(new_n933), .C2(new_n925), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n932), .A2(new_n934), .A3(new_n849), .ZN(G57));
endmodule


