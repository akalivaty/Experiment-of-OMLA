//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n985, new_n986, new_n987, new_n988,
    new_n989;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n202));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203));
  OR3_X1    g002(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n204));
  OAI21_X1  g003(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n205));
  INV_X1    g004(.A(G169gat), .ZN(new_n206));
  INV_X1    g005(.A(G176gat), .ZN(new_n207));
  OAI211_X1 g006(.A(new_n204), .B(new_n205), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT27), .B(G183gat), .ZN(new_n209));
  INV_X1    g008(.A(G190gat), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT28), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G183gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT27), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT27), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G183gat), .ZN(new_n215));
  AND4_X1   g014(.A1(KEYINPUT28), .A2(new_n213), .A3(new_n215), .A4(new_n210), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n203), .B(new_n208), .C1(new_n211), .C2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(new_n203), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n220));
  NAND3_X1  g019(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n223), .A2(new_n206), .A3(new_n207), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n206), .A2(new_n207), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n224), .B(new_n220), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n222), .A2(new_n227), .A3(KEYINPUT25), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT25), .B1(new_n222), .B2(new_n227), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n217), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G134gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT65), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G134gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n234), .A3(G127gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n231), .A2(G127gat), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G120gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G113gat), .ZN(new_n240));
  INV_X1    g039(.A(G113gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G120gat), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT1), .B1(new_n240), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(KEYINPUT66), .B1(new_n241), .B2(G120gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n246), .A2(new_n239), .A3(G113gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(new_n247), .A3(new_n242), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT1), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n249), .B1(new_n231), .B2(G127gat), .ZN(new_n250));
  INV_X1    g049(.A(G127gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n251), .A2(G134gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n238), .A2(new_n244), .B1(new_n248), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n248), .A2(new_n253), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT65), .B(G134gat), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n236), .B1(new_n258), .B2(G127gat), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n257), .B1(new_n259), .B2(new_n243), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT67), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n230), .A2(new_n256), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n222), .A2(new_n227), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT25), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n222), .A2(new_n227), .A3(KEYINPUT25), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n267), .A2(KEYINPUT67), .A3(new_n260), .A4(new_n217), .ZN(new_n268));
  INV_X1    g067(.A(G227gat), .ZN(new_n269));
  INV_X1    g068(.A(G233gat), .ZN(new_n270));
  NOR2_X1   g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n262), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G15gat), .B(G43gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(G71gat), .B(G99gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT33), .ZN(new_n276));
  OR2_X1    g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n272), .A2(KEYINPUT32), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT68), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT68), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n272), .A2(new_n280), .A3(KEYINPUT32), .A4(new_n277), .ZN(new_n281));
  AND2_X1   g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT34), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n262), .A2(new_n268), .ZN(new_n284));
  INV_X1    g083(.A(new_n271), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n283), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  AOI211_X1 g085(.A(KEYINPUT34), .B(new_n271), .C1(new_n262), .C2(new_n268), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n275), .B1(new_n272), .B2(KEYINPUT32), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n276), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n202), .B1(new_n282), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n279), .A2(new_n281), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n294), .A2(KEYINPUT69), .A3(new_n288), .A4(new_n291), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n279), .A2(new_n281), .B1(new_n290), .B2(new_n289), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(new_n288), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT36), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(KEYINPUT70), .A3(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n288), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n294), .A2(new_n291), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n288), .A2(new_n291), .ZN(new_n305));
  AOI22_X1  g104(.A1(new_n303), .A2(new_n304), .B1(new_n305), .B2(new_n294), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT36), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n298), .B1(new_n293), .B2(new_n295), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n308), .B1(new_n309), .B2(KEYINPUT36), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n302), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT38), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT29), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n230), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G226gat), .A2(G233gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n315), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n230), .A2(KEYINPUT71), .A3(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT71), .B1(new_n230), .B2(new_n317), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n316), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G197gat), .B(G204gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(G211gat), .A2(G218gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT22), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  OR2_X1    g124(.A1(G211gat), .A2(G218gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n322), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n322), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(new_n321), .A3(new_n324), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n320), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n327), .A2(new_n329), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n230), .A2(new_n317), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n316), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(KEYINPUT72), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT72), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n316), .A2(new_n336), .A3(new_n332), .A4(new_n333), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n331), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n312), .B1(new_n338), .B2(KEYINPUT37), .ZN(new_n339));
  XOR2_X1   g138(.A(G8gat), .B(G36gat), .Z(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(KEYINPUT73), .ZN(new_n341));
  XNOR2_X1  g140(.A(G64gat), .B(G92gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n341), .B(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n330), .A2(new_n320), .B1(new_n334), .B2(KEYINPUT72), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT37), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(new_n337), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n339), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n320), .A2(new_n332), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n316), .A2(new_n330), .A3(new_n333), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n349), .A2(KEYINPUT37), .A3(new_n350), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n344), .B(new_n351), .C1(new_n338), .C2(KEYINPUT37), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(new_n312), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(G1gat), .B(G29gat), .ZN(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(KEYINPUT0), .ZN(new_n356));
  XNOR2_X1  g155(.A(G57gat), .B(G85gat), .ZN(new_n357));
  XOR2_X1   g156(.A(new_n356), .B(new_n357), .Z(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  AND2_X1   g158(.A1(KEYINPUT78), .A2(G155gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(KEYINPUT78), .A2(G155gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(G162gat), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT2), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(G148gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT76), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT76), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(G148gat), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n366), .A2(new_n368), .A3(G141gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n365), .A2(G141gat), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT77), .ZN(new_n373));
  AND2_X1   g172(.A1(G155gat), .A2(G162gat), .ZN(new_n374));
  NOR2_X1   g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n373), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G155gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n363), .ZN(new_n378));
  NAND2_X1  g177(.A1(G155gat), .A2(G162gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(KEYINPUT77), .A3(new_n379), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n364), .A2(new_n372), .A3(new_n376), .A4(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT74), .B1(new_n374), .B2(new_n375), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT74), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n378), .A2(new_n383), .A3(new_n379), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT75), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n379), .A2(KEYINPUT2), .ZN(new_n387));
  INV_X1    g186(.A(G141gat), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n388), .A2(G148gat), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n387), .B1(new_n370), .B2(new_n389), .ZN(new_n390));
  AND3_X1   g189(.A1(new_n385), .A2(new_n386), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n386), .B1(new_n385), .B2(new_n390), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n381), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT3), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT79), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n248), .A2(new_n253), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n240), .A2(new_n242), .ZN(new_n397));
  AOI22_X1  g196(.A1(new_n235), .A2(new_n237), .B1(new_n397), .B2(new_n249), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n395), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n257), .B(KEYINPUT79), .C1(new_n259), .C2(new_n243), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n403), .B(new_n381), .C1(new_n391), .C2(new_n392), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n394), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n254), .B(new_n381), .C1(new_n391), .C2(new_n392), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G225gat), .A2(G233gat), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n374), .A2(new_n375), .A3(KEYINPUT74), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n383), .B1(new_n378), .B2(new_n379), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n390), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT75), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n385), .A2(new_n386), .A3(new_n390), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n415), .A2(KEYINPUT4), .A3(new_n381), .A4(new_n254), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n408), .A2(new_n409), .A3(new_n416), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n405), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT81), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n393), .A2(new_n399), .A3(new_n400), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n409), .B1(new_n420), .B2(new_n406), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT5), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n419), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(KEYINPUT76), .B(G148gat), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n370), .B1(new_n424), .B2(G141gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n376), .A2(new_n380), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n413), .A2(new_n414), .B1(new_n427), .B2(new_n364), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n406), .B1(new_n428), .B2(new_n401), .ZN(new_n429));
  INV_X1    g228(.A(new_n409), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n431), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n418), .B1(new_n423), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n407), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n428), .A2(new_n254), .A3(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT4), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n406), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NOR4_X1   g237(.A1(new_n405), .A2(new_n438), .A3(KEYINPUT5), .A4(new_n430), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n359), .B1(new_n433), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n394), .A2(new_n402), .A3(new_n404), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n441), .A2(new_n408), .A3(new_n409), .A4(new_n416), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT81), .B1(new_n431), .B2(KEYINPUT5), .ZN(new_n443));
  AOI211_X1 g242(.A(new_n419), .B(new_n422), .C1(new_n429), .C2(new_n430), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n405), .A2(new_n438), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n446), .A2(new_n422), .A3(new_n409), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n445), .A2(new_n358), .A3(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(KEYINPUT82), .B(KEYINPUT6), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n440), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n449), .ZN(new_n451));
  OAI211_X1 g250(.A(new_n359), .B(new_n451), .C1(new_n433), .C2(new_n439), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n331), .A2(new_n335), .A3(new_n337), .A4(new_n343), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n354), .A2(new_n450), .A3(new_n452), .A4(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(G228gat), .A2(G233gat), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n404), .A2(new_n313), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n330), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n403), .B1(new_n330), .B2(KEYINPUT29), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n393), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n456), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n332), .B1(new_n404), .B2(new_n313), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT3), .B1(new_n332), .B2(new_n313), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n428), .A2(new_n463), .ZN(new_n464));
  NOR3_X1   g263(.A1(new_n462), .A2(new_n464), .A3(new_n455), .ZN(new_n465));
  OAI21_X1  g264(.A(G22gat), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT29), .B1(new_n428), .B2(new_n403), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n456), .B(new_n460), .C1(new_n467), .C2(new_n332), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n455), .B1(new_n462), .B2(new_n464), .ZN(new_n469));
  INV_X1    g268(.A(G22gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  XNOR2_X1  g270(.A(G78gat), .B(G106gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(KEYINPUT31), .B(G50gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n466), .A2(KEYINPUT83), .A3(new_n471), .A4(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT83), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n478), .A2(new_n474), .B1(new_n466), .B2(new_n471), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT39), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n481), .B(new_n430), .C1(new_n405), .C2(new_n438), .ZN(new_n482));
  INV_X1    g281(.A(new_n438), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n409), .B1(new_n483), .B2(new_n441), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT39), .B1(new_n429), .B2(new_n430), .ZN(new_n485));
  OAI211_X1 g284(.A(new_n482), .B(new_n358), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT40), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n485), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n489), .B1(new_n446), .B2(new_n409), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n490), .A2(KEYINPUT40), .A3(new_n358), .A4(new_n482), .ZN(new_n491));
  AND3_X1   g290(.A1(new_n488), .A2(new_n440), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT30), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n453), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n345), .A2(KEYINPUT30), .A3(new_n337), .A4(new_n343), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n338), .A2(new_n344), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n480), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n450), .A2(new_n452), .ZN(new_n499));
  INV_X1    g298(.A(new_n497), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n454), .A2(new_n498), .B1(new_n501), .B2(new_n480), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT84), .ZN(new_n503));
  OAI22_X1  g302(.A1(new_n288), .A2(new_n297), .B1(new_n282), .B2(new_n292), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n503), .B1(new_n480), .B2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n497), .B1(new_n450), .B2(new_n452), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n478), .A2(new_n474), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n466), .A2(new_n471), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n475), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n510), .A2(new_n306), .A3(KEYINPUT84), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n505), .A2(new_n506), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT35), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n480), .A2(KEYINPUT35), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n506), .A2(new_n514), .A3(new_n309), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n311), .A2(new_n502), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G113gat), .B(G141gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(KEYINPUT85), .B(G197gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT11), .B(G169gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(new_n521), .B(KEYINPUT12), .Z(new_n522));
  INV_X1    g321(.A(KEYINPUT15), .ZN(new_n523));
  INV_X1    g322(.A(G50gat), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n523), .B1(G43gat), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(G43gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(G50gat), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT86), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT86), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n531), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT14), .ZN(new_n533));
  INV_X1    g332(.A(G29gat), .ZN(new_n534));
  INV_X1    g333(.A(G36gat), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n530), .A2(new_n532), .A3(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n534), .A2(new_n535), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n528), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n526), .A2(KEYINPUT87), .A3(G50gat), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT87), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(new_n526), .B2(G50gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n524), .A2(G43gat), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n523), .B(new_n540), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n538), .B1(new_n525), .B2(new_n527), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n536), .A2(KEYINPUT88), .ZN(new_n546));
  NOR3_X1   g345(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT88), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n529), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n544), .B(new_n545), .C1(new_n546), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n539), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G8gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n470), .A2(G15gat), .ZN(new_n553));
  INV_X1    g352(.A(G15gat), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(G22gat), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT16), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n553), .B(new_n555), .C1(new_n556), .C2(G1gat), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT89), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n552), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G15gat), .B(G22gat), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n557), .B1(G1gat), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  OAI221_X1 g361(.A(new_n557), .B1(new_n558), .B2(new_n552), .C1(G1gat), .C2(new_n560), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n551), .B(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G229gat), .A2(G233gat), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n566), .B(KEYINPUT13), .Z(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n564), .A2(KEYINPUT90), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT90), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n562), .A2(new_n570), .A3(new_n563), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT17), .ZN(new_n572));
  AND3_X1   g371(.A1(new_n539), .A2(new_n572), .A3(new_n550), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n572), .B1(new_n539), .B2(new_n550), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n569), .B(new_n571), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  AOI22_X1  g374(.A1(new_n551), .A2(new_n564), .B1(G229gat), .B2(G233gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(KEYINPUT18), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT18), .B1(new_n575), .B2(new_n576), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT91), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n568), .B(new_n577), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n578), .A2(new_n579), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n522), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT92), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n522), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n577), .A2(new_n568), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n578), .A2(new_n583), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n584), .A2(new_n585), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT93), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n582), .A2(new_n588), .A3(KEYINPUT93), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n516), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G71gat), .B(G78gat), .Z(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT9), .ZN(new_n598));
  INV_X1    g397(.A(G71gat), .ZN(new_n599));
  INV_X1    g398(.A(G78gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n598), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G57gat), .B(G64gat), .Z(new_n602));
  NAND3_X1  g401(.A1(new_n597), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n601), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(new_n596), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT21), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G127gat), .B(G155gat), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n608), .B(new_n609), .Z(new_n610));
  INV_X1    g409(.A(new_n606), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n564), .B1(new_n611), .B2(KEYINPUT21), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n610), .B(new_n612), .Z(new_n613));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT94), .ZN(new_n615));
  XOR2_X1   g414(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G183gat), .B(G211gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n613), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G120gat), .B(G148gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(G176gat), .B(G204gat), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n621), .B(new_n622), .Z(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(G230gat), .A2(G233gat), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(G85gat), .A2(G92gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT7), .ZN(new_n628));
  NAND2_X1  g427(.A1(G99gat), .A2(G106gat), .ZN(new_n629));
  INV_X1    g428(.A(G85gat), .ZN(new_n630));
  INV_X1    g429(.A(G92gat), .ZN(new_n631));
  AOI22_X1  g430(.A1(KEYINPUT8), .A2(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(G99gat), .B(G106gat), .Z(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n633), .A2(new_n634), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n606), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n628), .A2(new_n632), .ZN(new_n639));
  INV_X1    g438(.A(new_n634), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n641), .A2(new_n605), .A3(new_n603), .A4(new_n635), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n638), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n636), .A2(new_n637), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n645), .A2(KEYINPUT10), .A3(new_n611), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n626), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n625), .B1(new_n638), .B2(new_n642), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n624), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n649), .A2(KEYINPUT98), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(KEYINPUT98), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n648), .B(KEYINPUT97), .Z(new_n653));
  NOR2_X1   g452(.A1(new_n647), .A2(new_n624), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n657));
  XOR2_X1   g456(.A(G190gat), .B(G218gat), .Z(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(KEYINPUT95), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT96), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n661), .B1(new_n645), .B2(new_n551), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n573), .A2(new_n574), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n662), .B1(new_n663), .B2(new_n645), .ZN(new_n664));
  XNOR2_X1  g463(.A(G134gat), .B(G162gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n659), .A2(new_n660), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n668));
  INV_X1    g467(.A(G232gat), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n668), .B1(new_n669), .B2(new_n270), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n667), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n666), .B(new_n671), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n620), .A2(new_n656), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n595), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n674), .A2(new_n499), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT99), .B(G1gat), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1324gat));
  INV_X1    g476(.A(new_n674), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n497), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT16), .B(G8gat), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT42), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n679), .A2(G8gat), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n681), .A2(new_n682), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(G1325gat));
  XNOR2_X1  g485(.A(new_n311), .B(KEYINPUT100), .ZN(new_n687));
  OAI21_X1  g486(.A(G15gat), .B1(new_n674), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n309), .A2(new_n554), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n688), .B1(new_n674), .B2(new_n689), .ZN(G1326gat));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n510), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT43), .B(G22gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  AOI22_X1  g492(.A1(new_n650), .A2(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n694));
  AND4_X1   g493(.A1(new_n595), .A2(new_n620), .A3(new_n672), .A4(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n499), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(new_n534), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT45), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699));
  INV_X1    g498(.A(new_n672), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n699), .B1(new_n516), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n501), .A2(new_n480), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n454), .A2(new_n498), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n311), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n300), .A2(KEYINPUT35), .A3(new_n480), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n512), .A2(KEYINPUT35), .B1(new_n705), .B2(new_n506), .ZN(new_n706));
  OAI211_X1 g505(.A(KEYINPUT44), .B(new_n672), .C1(new_n704), .C2(new_n706), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n620), .ZN(new_n709));
  INV_X1    g508(.A(new_n589), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n709), .A2(new_n710), .A3(new_n656), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(G29gat), .B1(new_n712), .B2(new_n499), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n713), .ZN(G1328gat));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n500), .A2(G36gat), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n695), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT102), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G36gat), .B1(new_n712), .B2(new_n500), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n695), .A2(new_n716), .ZN(new_n721));
  AOI21_X1  g520(.A(KEYINPUT101), .B1(new_n721), .B2(KEYINPUT46), .ZN(new_n722));
  AND3_X1   g521(.A1(new_n721), .A2(KEYINPUT101), .A3(KEYINPUT46), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n719), .B(new_n720), .C1(new_n722), .C2(new_n723), .ZN(G1329gat));
  AND3_X1   g523(.A1(new_n695), .A2(new_n526), .A3(new_n309), .ZN(new_n725));
  INV_X1    g524(.A(new_n687), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n708), .A2(new_n726), .A3(new_n711), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n725), .B1(new_n727), .B2(G43gat), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729));
  OR2_X1    g528(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n712), .A2(new_n311), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(new_n526), .ZN(new_n732));
  OAI22_X1  g531(.A1(KEYINPUT47), .A2(new_n728), .B1(new_n730), .B2(new_n732), .ZN(G1330gat));
  NOR2_X1   g532(.A1(new_n510), .A2(G50gat), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT103), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n695), .A2(new_n735), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n701), .A2(new_n707), .A3(new_n480), .A4(new_n711), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G50gat), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(KEYINPUT48), .Z(G1331gat));
  NAND4_X1  g539(.A1(new_n700), .A2(new_n710), .A3(new_n709), .A4(new_n656), .ZN(new_n741));
  OR3_X1    g540(.A1(new_n516), .A2(KEYINPUT104), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT104), .B1(new_n516), .B2(new_n741), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n696), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g546(.A(KEYINPUT49), .B(G64gat), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n745), .A2(new_n497), .A3(new_n748), .ZN(new_n749));
  OAI22_X1  g548(.A1(new_n744), .A2(new_n500), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT105), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1333gat));
  OAI21_X1  g552(.A(G71gat), .B1(new_n744), .B2(new_n687), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n309), .A2(new_n599), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n754), .B1(new_n744), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT50), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n756), .B(new_n757), .ZN(G1334gat));
  NOR2_X1   g557(.A1(new_n744), .A2(new_n510), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n759), .B(new_n600), .ZN(G1335gat));
  NAND2_X1  g559(.A1(new_n502), .A2(new_n311), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n513), .A2(new_n515), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n709), .A2(new_n589), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n763), .A2(KEYINPUT51), .A3(new_n672), .A4(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT107), .ZN(new_n766));
  OR2_X1    g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n763), .A2(new_n672), .A3(new_n764), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT51), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n765), .A2(new_n766), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n767), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n772), .A2(new_n630), .A3(new_n696), .A4(new_n656), .ZN(new_n773));
  INV_X1    g572(.A(new_n764), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(new_n694), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n701), .A2(new_n707), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT106), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n701), .A2(new_n707), .A3(KEYINPUT106), .A4(new_n775), .ZN(new_n779));
  AND3_X1   g578(.A1(new_n778), .A2(new_n696), .A3(new_n779), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n773), .B1(new_n630), .B2(new_n780), .ZN(G1336gat));
  NOR3_X1   g580(.A1(new_n500), .A2(G92gat), .A3(new_n694), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n772), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  OAI21_X1  g583(.A(G92gat), .B1(new_n776), .B2(new_n500), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n778), .A2(new_n497), .A3(new_n779), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n765), .ZN(new_n788));
  AOI22_X1  g587(.A1(new_n787), .A2(G92gat), .B1(new_n788), .B2(new_n782), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n786), .B1(new_n789), .B2(new_n784), .ZN(G1337gat));
  NAND3_X1  g589(.A1(new_n778), .A2(new_n726), .A3(new_n779), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G99gat), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n300), .A2(G99gat), .A3(new_n694), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n772), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT108), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT108), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n792), .A2(new_n797), .A3(new_n794), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(G1338gat));
  NOR3_X1   g598(.A1(new_n510), .A2(G106gat), .A3(new_n694), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n772), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n802));
  OAI21_X1  g601(.A(G106gat), .B1(new_n776), .B2(new_n510), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n778), .A2(new_n480), .A3(new_n779), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n800), .B(KEYINPUT109), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n805), .A2(G106gat), .B1(new_n788), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n804), .B1(new_n807), .B2(new_n802), .ZN(G1339gat));
  NAND2_X1  g607(.A1(new_n644), .A2(new_n646), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n625), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n644), .A2(new_n626), .A3(new_n646), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(KEYINPUT54), .A3(new_n811), .ZN(new_n812));
  XOR2_X1   g611(.A(KEYINPUT110), .B(KEYINPUT54), .Z(new_n813));
  AOI21_X1  g612(.A(new_n623), .B1(new_n647), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n812), .A2(KEYINPUT55), .A3(new_n814), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n817), .A2(new_n655), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n589), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n551), .A2(new_n564), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n566), .B1(new_n575), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n565), .A2(new_n567), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n521), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n588), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n656), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n672), .B1(new_n820), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n819), .A2(new_n826), .A3(new_n672), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n620), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n673), .A2(new_n710), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n480), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT111), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n833), .A2(new_n834), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n499), .A2(new_n497), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n309), .ZN(new_n840));
  NOR4_X1   g639(.A1(new_n838), .A2(new_n241), .A3(new_n594), .A4(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n831), .A2(new_n832), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n505), .A2(new_n511), .ZN(new_n843));
  AND4_X1   g642(.A1(new_n696), .A2(new_n842), .A3(new_n500), .A4(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(G113gat), .B1(new_n844), .B2(new_n589), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n846), .B(KEYINPUT112), .ZN(G1340gat));
  AOI21_X1  g646(.A(G120gat), .B1(new_n844), .B2(new_n656), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n838), .A2(new_n840), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n694), .A2(new_n239), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(G1341gat));
  NAND3_X1  g650(.A1(new_n844), .A2(new_n251), .A3(new_n709), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n838), .A2(new_n620), .A3(new_n840), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n251), .ZN(G1342gat));
  NAND3_X1  g653(.A1(new_n844), .A2(new_n258), .A3(new_n672), .ZN(new_n855));
  XOR2_X1   g654(.A(new_n855), .B(KEYINPUT56), .Z(new_n856));
  INV_X1    g655(.A(KEYINPUT113), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n849), .A2(new_n672), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n857), .B1(new_n858), .B2(G134gat), .ZN(new_n859));
  AOI211_X1 g658(.A(KEYINPUT113), .B(new_n231), .C1(new_n849), .C2(new_n672), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n856), .B1(new_n859), .B2(new_n860), .ZN(G1343gat));
  NAND2_X1  g660(.A1(new_n311), .A2(new_n839), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(KEYINPUT114), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n582), .A2(new_n588), .A3(KEYINPUT93), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT93), .B1(new_n582), .B2(new_n588), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n819), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n672), .B1(new_n867), .B2(new_n827), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n620), .B1(new_n868), .B2(new_n830), .ZN(new_n869));
  AOI211_X1 g668(.A(new_n864), .B(new_n510), .C1(new_n869), .C2(new_n832), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT57), .B1(new_n842), .B2(new_n480), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n863), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(G141gat), .B1(new_n872), .B2(new_n594), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n842), .A2(new_n696), .A3(new_n500), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n726), .A2(new_n510), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n388), .A3(new_n593), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n873), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(G141gat), .B1(new_n872), .B2(new_n710), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n876), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n880), .A2(KEYINPUT115), .A3(KEYINPUT58), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT115), .B1(new_n880), .B2(KEYINPUT58), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n878), .B1(new_n881), .B2(new_n882), .ZN(G1344gat));
  NAND3_X1  g682(.A1(new_n875), .A2(new_n424), .A3(new_n656), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(KEYINPUT116), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n594), .A2(new_n673), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n510), .B1(new_n869), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT117), .B1(new_n887), .B2(KEYINPUT57), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT117), .ZN(new_n889));
  INV_X1    g688(.A(new_n886), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n694), .A2(new_n825), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n891), .B1(new_n593), .B2(new_n819), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n829), .B1(new_n892), .B2(new_n672), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n890), .B1(new_n893), .B2(new_n620), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n889), .B(new_n864), .C1(new_n894), .C2(new_n510), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n842), .A2(KEYINPUT57), .A3(new_n480), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n888), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n863), .A2(new_n656), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n365), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT118), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n424), .A2(KEYINPUT59), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n902), .B1(new_n872), .B2(new_n694), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n899), .A2(KEYINPUT118), .A3(new_n900), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n885), .B1(new_n904), .B2(new_n905), .ZN(G1345gat));
  NAND3_X1  g705(.A1(new_n875), .A2(new_n362), .A3(new_n709), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n872), .A2(new_n620), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(new_n362), .ZN(G1346gat));
  NAND3_X1  g708(.A1(new_n875), .A2(new_n363), .A3(new_n672), .ZN(new_n910));
  XOR2_X1   g709(.A(new_n910), .B(KEYINPUT119), .Z(new_n911));
  OAI21_X1  g710(.A(G162gat), .B1(new_n872), .B2(new_n700), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1347gat));
  NAND2_X1  g712(.A1(new_n843), .A2(new_n497), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n914), .A2(KEYINPUT120), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n696), .B1(new_n831), .B2(new_n832), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(KEYINPUT120), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n206), .B1(new_n918), .B2(new_n710), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n836), .A2(new_n837), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n696), .A2(new_n500), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(new_n300), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n593), .A2(G169gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n919), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT121), .Z(G1348gat));
  OAI21_X1  g726(.A(G176gat), .B1(new_n924), .B2(new_n694), .ZN(new_n928));
  INV_X1    g727(.A(new_n918), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(new_n207), .A3(new_n656), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(G1349gat));
  INV_X1    g730(.A(KEYINPUT122), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT60), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n709), .A2(new_n209), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n933), .B1(new_n918), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n920), .A2(new_n709), .A3(new_n923), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n936), .B2(G183gat), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n932), .A2(KEYINPUT60), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n937), .B(new_n938), .ZN(G1350gat));
  NAND3_X1  g738(.A1(new_n929), .A2(new_n210), .A3(new_n672), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n920), .A2(new_n672), .A3(new_n923), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT61), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n941), .A2(new_n942), .A3(G190gat), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n942), .B1(new_n941), .B2(G190gat), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(G1351gat));
  AND2_X1   g744(.A1(new_n311), .A2(KEYINPUT100), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n311), .A2(KEYINPUT100), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n497), .B(new_n480), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT123), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT123), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n687), .A2(new_n950), .A3(new_n497), .A4(new_n480), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n949), .A2(new_n916), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(G197gat), .B1(new_n952), .B2(new_n589), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n687), .A2(new_n921), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT124), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n897), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g755(.A1(new_n888), .A2(new_n895), .A3(KEYINPUT124), .A4(new_n896), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n593), .A2(G197gat), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n953), .B1(new_n958), .B2(new_n959), .ZN(G1352gat));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n961));
  INV_X1    g760(.A(G204gat), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n956), .A2(new_n957), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n954), .A2(new_n694), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n694), .A2(G204gat), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n949), .A2(new_n951), .A3(new_n916), .A4(new_n966), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n967), .B(KEYINPUT62), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n961), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT62), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n967), .B(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(new_n964), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n972), .B1(new_n956), .B2(new_n957), .ZN(new_n973));
  OAI211_X1 g772(.A(new_n971), .B(KEYINPUT125), .C1(new_n962), .C2(new_n973), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n969), .A2(new_n974), .ZN(G1353gat));
  OAI21_X1  g774(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n954), .A2(new_n620), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n976), .B1(new_n897), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n979));
  OR2_X1    g778(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n979), .ZN(new_n981));
  INV_X1    g780(.A(G211gat), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n952), .A2(new_n982), .A3(new_n709), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n980), .A2(new_n981), .A3(new_n983), .ZN(G1354gat));
  AOI21_X1  g783(.A(G218gat), .B1(new_n952), .B2(new_n672), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT127), .ZN(new_n986));
  OR2_X1    g785(.A1(new_n958), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n672), .A2(G218gat), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n988), .B1(new_n958), .B2(new_n986), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n985), .B1(new_n987), .B2(new_n989), .ZN(G1355gat));
endmodule


