//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 1 0 1 1 1 0 0 1 0 0 0 1 1 1 1 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:16 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n599, new_n600, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017;
  INV_X1    g000(.A(G953), .ZN(new_n187));
  NAND3_X1  g001(.A1(new_n187), .A2(G221), .A3(G234), .ZN(new_n188));
  OR2_X1    g002(.A1(new_n188), .A2(KEYINPUT73), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(KEYINPUT73), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT22), .B(G137), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n189), .A2(new_n192), .A3(new_n190), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT74), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(KEYINPUT74), .A3(new_n195), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G140), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT16), .ZN(new_n205));
  OR3_X1    g019(.A1(new_n203), .A2(KEYINPUT16), .A3(G140), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n205), .A2(new_n206), .A3(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G128), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n212), .B(G119), .C1(KEYINPUT72), .C2(KEYINPUT23), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT23), .ZN(new_n214));
  INV_X1    g028(.A(G119), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n214), .B1(new_n215), .B2(G128), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT72), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n217), .B1(new_n215), .B2(G128), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n213), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g033(.A(G119), .B(G128), .ZN(new_n220));
  XOR2_X1   g034(.A(KEYINPUT24), .B(G110), .Z(new_n221));
  AOI22_X1  g035(.A1(new_n219), .A2(G110), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n211), .A2(new_n222), .ZN(new_n223));
  OAI22_X1  g037(.A1(new_n219), .A2(G110), .B1(new_n220), .B2(new_n221), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n202), .A2(new_n204), .A3(new_n208), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n224), .A2(new_n210), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n200), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n223), .A2(new_n226), .A3(new_n196), .ZN(new_n229));
  AND2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XOR2_X1   g044(.A(KEYINPUT71), .B(G217), .Z(new_n231));
  INV_X1    g045(.A(G234), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(G902), .ZN(new_n233));
  INV_X1    g047(.A(G902), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n230), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n237), .B(KEYINPUT75), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n228), .A2(new_n234), .A3(new_n229), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n233), .B1(new_n239), .B2(KEYINPUT25), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n228), .A2(new_n241), .A3(new_n234), .A4(new_n229), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G137), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT11), .ZN(new_n246));
  INV_X1    g060(.A(G134), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT64), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT64), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G134), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n246), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  OR2_X1    g065(.A1(new_n245), .A2(KEYINPUT11), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n245), .A2(KEYINPUT11), .A3(G134), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(G131), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n246), .A2(new_n248), .A3(new_n250), .ZN(new_n256));
  INV_X1    g070(.A(G131), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n256), .A2(new_n257), .A3(new_n253), .A4(new_n252), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n255), .A2(KEYINPUT65), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n208), .A2(G143), .ZN(new_n260));
  INV_X1    g074(.A(G143), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G146), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n260), .A2(new_n262), .A3(KEYINPUT0), .A4(G128), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n260), .A2(new_n262), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT0), .B(G128), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n263), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n269), .B(G131), .C1(new_n251), .C2(new_n254), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n259), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n215), .A2(G116), .ZN(new_n272));
  INV_X1    g086(.A(G116), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G119), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  XOR2_X1   g089(.A(KEYINPUT2), .B(G113), .Z(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n272), .A2(new_n274), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT2), .B(G113), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n247), .A2(G137), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT64), .B(G134), .ZN(new_n284));
  OAI211_X1 g098(.A(KEYINPUT66), .B(new_n283), .C1(new_n284), .C2(G137), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n248), .A2(new_n250), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n245), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n285), .B(G131), .C1(KEYINPUT66), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n260), .A2(KEYINPUT1), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n264), .A2(new_n289), .A3(G128), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n260), .B(new_n262), .C1(KEYINPUT1), .C2(new_n212), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n288), .A2(new_n258), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n271), .A2(new_n282), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT68), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n271), .A2(new_n294), .A3(KEYINPUT68), .A4(new_n282), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n271), .A2(new_n294), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(new_n281), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT28), .ZN(new_n302));
  INV_X1    g116(.A(new_n295), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n303), .A2(KEYINPUT28), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(G237), .A2(G953), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G210), .ZN(new_n308));
  XOR2_X1   g122(.A(new_n308), .B(KEYINPUT27), .Z(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT26), .B(G101), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n309), .B(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n306), .A2(KEYINPUT69), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT69), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n304), .B1(new_n301), .B2(KEYINPUT28), .ZN(new_n314));
  INV_X1    g128(.A(new_n311), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT67), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n299), .A2(new_n317), .A3(KEYINPUT30), .ZN(new_n318));
  OR2_X1    g132(.A1(new_n317), .A2(KEYINPUT30), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(KEYINPUT30), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n271), .A2(new_n294), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n282), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n297), .A2(new_n298), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(KEYINPUT31), .B1(new_n324), .B2(new_n315), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT31), .ZN(new_n326));
  NOR4_X1   g140(.A1(new_n322), .A2(new_n323), .A3(new_n326), .A4(new_n311), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n312), .B(new_n316), .C1(new_n325), .C2(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(G472), .A2(G902), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT32), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT32), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n328), .A2(new_n332), .A3(new_n329), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n318), .A2(new_n321), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n281), .ZN(new_n336));
  INV_X1    g150(.A(new_n323), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(KEYINPUT29), .B1(new_n338), .B2(new_n311), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n314), .A2(new_n315), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n234), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n302), .A2(KEYINPUT70), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n305), .B1(new_n302), .B2(KEYINPUT70), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n315), .A2(KEYINPUT29), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(G472), .B1(new_n342), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n244), .B1(new_n334), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(G113), .B(G122), .ZN(new_n349));
  INV_X1    g163(.A(G104), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n349), .B(new_n350), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n307), .A2(G143), .A3(G214), .ZN(new_n352));
  AOI21_X1  g166(.A(G143), .B1(new_n307), .B2(G214), .ZN(new_n353));
  OAI211_X1 g167(.A(KEYINPUT18), .B(G131), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n202), .A2(new_n204), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G146), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n225), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n307), .A2(G214), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n261), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n307), .A2(G143), .A3(G214), .ZN(new_n360));
  NAND2_X1  g174(.A1(KEYINPUT18), .A2(G131), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n354), .A2(new_n357), .A3(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(G131), .B1(new_n352), .B2(new_n353), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n359), .A2(new_n257), .A3(new_n360), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT17), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  OAI211_X1 g181(.A(KEYINPUT17), .B(G131), .C1(new_n352), .C2(new_n353), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n209), .A2(new_n368), .A3(new_n210), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n351), .B(new_n363), .C1(new_n367), .C2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n373), .A2(new_n209), .A3(new_n210), .A4(new_n368), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n374), .A2(KEYINPUT81), .A3(new_n351), .A4(new_n363), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n364), .A2(new_n365), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT19), .ZN(new_n378));
  AOI21_X1  g192(.A(KEYINPUT19), .B1(new_n202), .B2(new_n204), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n208), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n377), .A2(new_n380), .A3(new_n210), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n351), .B1(new_n381), .B2(new_n363), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n376), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT20), .ZN(new_n385));
  NOR2_X1   g199(.A1(G475), .A2(G902), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT82), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n384), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n376), .A2(KEYINPUT82), .A3(new_n383), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n386), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n388), .B1(new_n392), .B2(KEYINPUT20), .ZN(new_n393));
  INV_X1    g207(.A(G475), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n374), .A2(new_n363), .ZN(new_n395));
  INV_X1    g209(.A(new_n351), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n376), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n394), .B1(new_n398), .B2(new_n234), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT83), .B1(new_n393), .B2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT83), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n398), .A2(new_n234), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G475), .ZN(new_n403));
  AOI21_X1  g217(.A(KEYINPUT82), .B1(new_n376), .B2(new_n383), .ZN(new_n404));
  AOI211_X1 g218(.A(new_n389), .B(new_n382), .C1(new_n372), .C2(new_n375), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n385), .B1(new_n406), .B2(new_n386), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n401), .B(new_n403), .C1(new_n407), .C2(new_n388), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n400), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT4), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n350), .A2(G107), .ZN(new_n411));
  NAND2_X1  g225(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NOR2_X1   g227(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n411), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G107), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(G104), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  OAI22_X1  g233(.A1(new_n350), .A2(G107), .B1(KEYINPUT77), .B2(KEYINPUT3), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n410), .B(G101), .C1(new_n416), .C2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G101), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n415), .A2(new_n423), .A3(new_n419), .A4(new_n420), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT4), .ZN(new_n425));
  INV_X1    g239(.A(new_n414), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n417), .A2(G104), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n418), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n423), .B1(new_n428), .B2(new_n415), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n268), .B(new_n422), .C1(new_n425), .C2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n259), .A2(new_n270), .ZN(new_n431));
  OAI21_X1  g245(.A(G101), .B1(new_n411), .B2(new_n418), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n293), .A2(KEYINPUT10), .A3(new_n424), .A4(new_n432), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n424), .A2(new_n291), .A3(new_n290), .A4(new_n432), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT10), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n430), .A2(new_n431), .A3(new_n433), .A4(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G110), .B(G140), .ZN(new_n438));
  INV_X1    g252(.A(G227), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(G953), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n438), .B(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n437), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n430), .A2(new_n433), .A3(new_n436), .ZN(new_n445));
  INV_X1    g259(.A(new_n431), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT78), .ZN(new_n449));
  INV_X1    g263(.A(new_n434), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n424), .A2(new_n432), .B1(new_n290), .B2(new_n291), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n270), .B(new_n259), .C1(new_n450), .C2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT12), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n449), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n453), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n424), .A2(new_n432), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n292), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n434), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n446), .A2(new_n458), .A3(KEYINPUT78), .A4(KEYINPUT12), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n454), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n460), .A2(new_n437), .ZN(new_n461));
  OAI211_X1 g275(.A(G469), .B(new_n448), .C1(new_n461), .C2(new_n442), .ZN(new_n462));
  INV_X1    g276(.A(G469), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n455), .A2(new_n459), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n443), .B1(new_n464), .B2(new_n454), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n442), .B1(new_n447), .B2(new_n437), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n463), .B(new_n234), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(G469), .A2(G902), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n462), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT9), .B(G234), .ZN(new_n470));
  OAI21_X1  g284(.A(G221), .B1(new_n470), .B2(G902), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n471), .B(KEYINPUT76), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n212), .A2(G143), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n212), .A2(G143), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n475), .B1(KEYINPUT13), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT84), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n247), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n475), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT13), .ZN(new_n481));
  OAI21_X1  g295(.A(KEYINPUT84), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n479), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n284), .A2(new_n480), .A3(new_n476), .ZN(new_n484));
  XNOR2_X1  g298(.A(G116), .B(G122), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(G107), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n417), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n484), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n273), .A2(KEYINPUT14), .A3(G122), .ZN(new_n491));
  OAI211_X1 g305(.A(G107), .B(new_n491), .C1(new_n486), .C2(KEYINPUT14), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n284), .B1(new_n480), .B2(new_n476), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n492), .B(new_n488), .C1(new_n484), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n470), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(new_n187), .A3(new_n231), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT85), .ZN(new_n499));
  INV_X1    g313(.A(new_n497), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n490), .A2(new_n494), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n498), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n495), .A2(KEYINPUT85), .A3(new_n497), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n234), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT15), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n505), .A3(G478), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(G478), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n502), .A2(new_n234), .A3(new_n503), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(G234), .A2(G237), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(G952), .A3(new_n187), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(G902), .A3(G953), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT21), .B(G898), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(G214), .B1(G237), .B2(G902), .ZN(new_n518));
  XNOR2_X1  g332(.A(G110), .B(G122), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(KEYINPUT8), .ZN(new_n520));
  INV_X1    g334(.A(G113), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n273), .A2(G119), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT5), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n272), .A2(new_n274), .A3(KEYINPUT5), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n275), .A2(new_n276), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n526), .A2(new_n424), .A3(new_n432), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n526), .B1(new_n424), .B2(new_n432), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n520), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n263), .B(G125), .C1(new_n265), .C2(new_n266), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n530), .B1(new_n292), .B2(G125), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n187), .A2(G224), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n531), .A2(new_n533), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT79), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n531), .A2(KEYINPUT79), .A3(new_n533), .ZN(new_n538));
  AND4_X1   g352(.A1(new_n529), .A2(new_n534), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n281), .B(new_n422), .C1(new_n425), .C2(new_n429), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n526), .A2(new_n424), .A3(new_n432), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n519), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(G902), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n541), .ZN(new_n544));
  INV_X1    g358(.A(new_n519), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(KEYINPUT6), .A3(new_n542), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT6), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n544), .A2(new_n548), .A3(new_n545), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n531), .B(new_n532), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n547), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(G210), .B1(G237), .B2(G902), .ZN(new_n552));
  OR2_X1    g366(.A1(new_n552), .A2(KEYINPUT80), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n543), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n553), .B1(new_n543), .B2(new_n551), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n517), .B(new_n518), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NOR4_X1   g370(.A1(new_n409), .A2(new_n474), .A3(new_n509), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n348), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(G101), .ZN(G3));
  NAND2_X1  g373(.A1(new_n328), .A2(new_n234), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G472), .ZN(new_n561));
  INV_X1    g375(.A(new_n474), .ZN(new_n562));
  INV_X1    g376(.A(new_n244), .ZN(new_n563));
  AND4_X1   g377(.A1(new_n330), .A2(new_n561), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT33), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n502), .A2(new_n565), .A3(new_n503), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n498), .A2(KEYINPUT33), .A3(new_n501), .ZN(new_n567));
  INV_X1    g381(.A(G478), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(G902), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n504), .A2(new_n568), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n570), .A2(KEYINPUT86), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT86), .B1(new_n570), .B2(new_n571), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(new_n400), .B2(new_n408), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n543), .A2(new_n551), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n552), .ZN(new_n577));
  INV_X1    g391(.A(new_n552), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n543), .A2(new_n551), .A3(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n577), .A2(new_n518), .A3(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(new_n516), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n564), .A2(new_n575), .A3(new_n581), .ZN(new_n582));
  XOR2_X1   g396(.A(KEYINPUT34), .B(G104), .Z(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(G6));
  NAND2_X1  g398(.A1(new_n403), .A2(KEYINPUT87), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT87), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n399), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n509), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n407), .ZN(new_n589));
  INV_X1    g403(.A(new_n386), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n404), .A2(new_n405), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n385), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n588), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n564), .A2(new_n581), .A3(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(KEYINPUT35), .B(G107), .Z(new_n595));
  XNOR2_X1  g409(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT88), .B(KEYINPUT89), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G9));
  INV_X1    g412(.A(KEYINPUT90), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n561), .A2(new_n330), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n200), .A2(KEYINPUT36), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(new_n227), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n236), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n603), .A2(new_n243), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n599), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n243), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n561), .A2(KEYINPUT90), .A3(new_n330), .A4(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n605), .A2(new_n557), .A3(new_n607), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT37), .B(G110), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G12));
  AND3_X1   g424(.A1(new_n328), .A2(new_n332), .A3(new_n329), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n332), .B1(new_n328), .B2(new_n329), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n347), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n588), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n589), .A2(new_n592), .ZN(new_n615));
  INV_X1    g429(.A(G900), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n514), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n511), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n614), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n474), .A2(new_n580), .A3(new_n604), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n613), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G128), .ZN(G30));
  INV_X1    g437(.A(new_n518), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n393), .A2(KEYINPUT83), .A3(new_n399), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n387), .B1(new_n591), .B2(new_n385), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n401), .B1(new_n626), .B2(new_n403), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n509), .B1(new_n625), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n554), .A2(new_n555), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(KEYINPUT38), .ZN(new_n630));
  OR4_X1    g444(.A1(new_n624), .A2(new_n628), .A3(new_n630), .A4(new_n606), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n324), .A2(new_n311), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n234), .B1(new_n301), .B2(new_n315), .ZN(new_n633));
  OAI21_X1  g447(.A(G472), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT91), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n635), .B1(new_n611), .B2(new_n612), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  OR3_X1    g451(.A1(new_n631), .A2(new_n637), .A3(KEYINPUT92), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT92), .B1(new_n631), .B2(new_n637), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n618), .B(KEYINPUT39), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n562), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(new_n641), .B(KEYINPUT40), .Z(new_n642));
  NAND3_X1  g456(.A1(new_n638), .A2(new_n639), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G143), .ZN(G45));
  INV_X1    g458(.A(new_n618), .ZN(new_n645));
  AOI211_X1 g459(.A(new_n645), .B(new_n574), .C1(new_n400), .C2(new_n408), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n613), .A2(new_n646), .A3(new_n621), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G146), .ZN(G48));
  OR2_X1    g462(.A1(new_n572), .A2(new_n573), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n466), .B1(new_n460), .B2(new_n444), .ZN(new_n650));
  OAI21_X1  g464(.A(G469), .B1(new_n650), .B2(G902), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n467), .A2(new_n651), .A3(new_n471), .ZN(new_n652));
  AND4_X1   g466(.A1(new_n409), .A2(new_n649), .A3(new_n581), .A4(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n613), .A3(new_n563), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT41), .B(G113), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(KEYINPUT93), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n654), .B(new_n656), .ZN(G15));
  AND3_X1   g471(.A1(new_n593), .A2(new_n581), .A3(new_n652), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n348), .A2(KEYINPUT94), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n613), .A2(new_n658), .A3(new_n563), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT94), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G116), .ZN(G18));
  NOR2_X1   g478(.A1(new_n604), .A2(new_n516), .ZN(new_n665));
  INV_X1    g479(.A(new_n509), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n400), .A2(new_n408), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n467), .A2(new_n651), .A3(new_n471), .ZN(new_n668));
  OAI21_X1  g482(.A(KEYINPUT95), .B1(new_n668), .B2(new_n580), .ZN(new_n669));
  AND3_X1   g483(.A1(new_n577), .A2(new_n518), .A3(new_n579), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT95), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n652), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n667), .B1(new_n669), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n613), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G119), .ZN(G21));
  INV_X1    g489(.A(KEYINPUT97), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n238), .A2(new_n676), .A3(new_n243), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n676), .B1(new_n238), .B2(new_n243), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n311), .B1(new_n343), .B2(new_n344), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n336), .A2(new_n337), .A3(new_n315), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n326), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n324), .A2(KEYINPUT31), .A3(new_n315), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n329), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n315), .B1(new_n302), .B2(new_n305), .ZN(new_n688));
  AOI22_X1  g502(.A1(new_n682), .A2(new_n683), .B1(new_n688), .B2(KEYINPUT69), .ZN(new_n689));
  AOI21_X1  g503(.A(G902), .B1(new_n689), .B2(new_n316), .ZN(new_n690));
  INV_X1    g504(.A(G472), .ZN(new_n691));
  OAI21_X1  g505(.A(KEYINPUT96), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT96), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n560), .A2(new_n693), .A3(G472), .ZN(new_n694));
  AOI211_X1 g508(.A(new_n679), .B(new_n687), .C1(new_n692), .C2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(KEYINPUT98), .B1(new_n409), .B2(new_n509), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT98), .ZN(new_n697));
  AOI211_X1 g511(.A(new_n697), .B(new_n666), .C1(new_n400), .C2(new_n408), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n581), .A2(new_n652), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n696), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n695), .A2(new_n700), .A3(KEYINPUT99), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT99), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n628), .A2(new_n697), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n409), .A2(KEYINPUT98), .A3(new_n509), .ZN(new_n704));
  INV_X1    g518(.A(new_n699), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n679), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n693), .B1(new_n560), .B2(G472), .ZN(new_n708));
  AOI211_X1 g522(.A(KEYINPUT96), .B(new_n691), .C1(new_n328), .C2(new_n234), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n707), .B(new_n686), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n702), .B1(new_n706), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n701), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G122), .ZN(G24));
  AOI21_X1  g527(.A(new_n687), .B1(new_n692), .B2(new_n694), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n672), .A2(new_n669), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n714), .A2(new_n606), .A3(new_n646), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G125), .ZN(G27));
  XNOR2_X1  g531(.A(new_n468), .B(KEYINPUT100), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n462), .A2(new_n467), .A3(new_n718), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n554), .A2(new_n555), .A3(new_n624), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n719), .A2(new_n720), .A3(new_n471), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n575), .A2(new_n618), .A3(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n722), .A2(KEYINPUT42), .A3(new_n613), .A4(new_n707), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n722), .A2(KEYINPUT101), .A3(new_n613), .A4(new_n563), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT42), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT101), .B1(new_n348), .B2(new_n722), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n723), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G131), .ZN(G33));
  OAI21_X1  g543(.A(new_n721), .B1(new_n619), .B2(KEYINPUT102), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT102), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n731), .B1(new_n593), .B2(new_n618), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n348), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G134), .ZN(G36));
  NOR2_X1   g549(.A1(new_n625), .A2(new_n627), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n649), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n737), .A2(KEYINPUT43), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(KEYINPUT43), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n600), .A2(new_n606), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT103), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n742), .A2(KEYINPUT103), .A3(new_n743), .ZN(new_n747));
  OR3_X1    g561(.A1(new_n740), .A2(new_n743), .A3(new_n741), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n448), .B1(new_n461), .B2(new_n442), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT45), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n463), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n750), .B2(new_n749), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(KEYINPUT46), .A3(new_n718), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n467), .ZN(new_n755));
  AOI21_X1  g569(.A(KEYINPUT46), .B1(new_n752), .B2(new_n718), .ZN(new_n756));
  OR3_X1    g570(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n471), .ZN(new_n758));
  INV_X1    g572(.A(new_n640), .ZN(new_n759));
  INV_X1    g573(.A(new_n720), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n746), .A2(new_n747), .A3(new_n748), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G137), .ZN(G39));
  NAND3_X1  g577(.A1(new_n757), .A2(KEYINPUT47), .A3(new_n471), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n765));
  NOR3_X1   g579(.A1(new_n754), .A2(new_n755), .A3(new_n756), .ZN(new_n766));
  INV_X1    g580(.A(new_n471), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n346), .ZN(new_n770));
  AOI21_X1  g584(.A(G902), .B1(new_n339), .B2(new_n340), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n691), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n772), .B1(new_n331), .B2(new_n333), .ZN(new_n773));
  AND4_X1   g587(.A1(new_n773), .A2(new_n244), .A3(new_n646), .A4(new_n720), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G140), .ZN(G42));
  NOR3_X1   g590(.A1(new_n740), .A2(new_n511), .A3(new_n710), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n467), .A2(new_n651), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n473), .ZN(new_n779));
  OAI211_X1 g593(.A(new_n720), .B(new_n777), .C1(new_n769), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n760), .A2(new_n668), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n738), .A2(new_n512), .A3(new_n739), .A4(new_n781), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n606), .B(new_n686), .C1(new_n708), .C2(new_n709), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n637), .A2(new_n563), .A3(new_n512), .A4(new_n781), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n736), .A2(new_n574), .ZN(new_n785));
  OAI22_X1  g599(.A1(new_n782), .A2(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n630), .A2(new_n624), .A3(new_n652), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n777), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT50), .B1(new_n777), .B2(new_n788), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n780), .B(new_n787), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT51), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT108), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n793), .A2(KEYINPUT108), .A3(new_n794), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n613), .A2(new_n707), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n782), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g615(.A(new_n801), .B(KEYINPUT48), .Z(new_n802));
  INV_X1    g616(.A(new_n575), .ZN(new_n803));
  OAI211_X1 g617(.A(G952), .B(new_n187), .C1(new_n784), .C2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n804), .B1(new_n777), .B2(new_n715), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n780), .A2(KEYINPUT51), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n789), .B(new_n790), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT109), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n786), .A2(new_n809), .ZN(new_n810));
  OAI221_X1 g624(.A(KEYINPUT109), .B1(new_n784), .B2(new_n785), .C1(new_n782), .C2(new_n783), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n807), .A2(new_n808), .A3(KEYINPUT110), .A4(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT110), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n780), .A2(KEYINPUT51), .A3(new_n810), .A4(new_n811), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n791), .A2(new_n792), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n806), .B1(new_n813), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n799), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT111), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n723), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n575), .A2(new_n721), .A3(new_n618), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n773), .A2(new_n823), .A3(new_n244), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT42), .B1(new_n824), .B2(KEYINPUT101), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n348), .A2(new_n722), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT101), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n822), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n409), .A2(new_n509), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n649), .B1(new_n408), .B2(new_n400), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n830), .A2(new_n831), .A3(new_n556), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n564), .A2(new_n832), .B1(new_n348), .B2(new_n557), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n585), .A2(new_n587), .ZN(new_n834));
  NOR4_X1   g648(.A1(new_n834), .A2(new_n604), .A3(new_n509), .A4(new_n645), .ZN(new_n835));
  AND4_X1   g649(.A1(new_n562), .A2(new_n835), .A3(new_n615), .A4(new_n720), .ZN(new_n836));
  AOI22_X1  g650(.A1(new_n348), .A2(new_n733), .B1(new_n613), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n714), .A2(new_n606), .A3(new_n722), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n833), .A2(new_n837), .A3(new_n838), .A4(new_n608), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n829), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT99), .B1(new_n695), .B2(new_n700), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n706), .A2(new_n710), .A3(new_n702), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n348), .A2(new_n653), .B1(new_n613), .B2(new_n673), .ZN(new_n844));
  AOI21_X1  g658(.A(KEYINPUT94), .B1(new_n348), .B2(new_n658), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n660), .A2(new_n661), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(KEYINPUT104), .B1(new_n843), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n654), .A2(new_n674), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n849), .B1(new_n662), .B2(new_n659), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT104), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n850), .A2(new_n712), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n696), .A2(new_n698), .ZN(new_n853));
  AND4_X1   g667(.A1(new_n471), .A2(new_n719), .A3(new_n604), .A4(new_n618), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n853), .A2(new_n670), .A3(new_n636), .A4(new_n854), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n613), .B(new_n621), .C1(new_n646), .C2(new_n620), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n855), .A2(new_n716), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n855), .A2(new_n716), .A3(KEYINPUT52), .A4(new_n856), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n840), .A2(new_n848), .A3(new_n852), .A4(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n832), .A2(new_n564), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n608), .A2(new_n558), .A3(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n867), .A2(KEYINPUT107), .A3(new_n838), .A4(new_n837), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT107), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n839), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  AND4_X1   g685(.A1(KEYINPUT53), .A2(new_n728), .A3(new_n712), .A4(new_n850), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n646), .A2(new_n715), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n856), .B1(new_n783), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n703), .A2(new_n670), .A3(new_n704), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n636), .A2(new_n854), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(KEYINPUT106), .B(new_n858), .C1(new_n874), .C2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT106), .B1(new_n857), .B2(new_n858), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n874), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n882), .A2(KEYINPUT105), .A3(KEYINPUT52), .A4(new_n855), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT105), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n860), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n871), .B(new_n872), .C1(new_n881), .C2(new_n886), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n864), .A2(new_n865), .A3(new_n887), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n881), .A2(new_n886), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n848), .A2(new_n852), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n889), .A2(new_n863), .A3(new_n890), .A4(new_n840), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n862), .A2(KEYINPUT53), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n888), .B1(new_n893), .B2(KEYINPUT54), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n799), .A2(new_n818), .A3(KEYINPUT111), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n821), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT112), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT112), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n821), .A2(new_n894), .A3(new_n898), .A4(new_n895), .ZN(new_n899));
  OR2_X1    g713(.A1(G952), .A2(G953), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n897), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n679), .A2(new_n472), .A3(new_n624), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n778), .A2(KEYINPUT49), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n778), .A2(KEYINPUT49), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n902), .A2(new_n630), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  OR3_X1    g719(.A1(new_n905), .A2(new_n636), .A3(new_n737), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n901), .A2(new_n906), .ZN(G75));
  NOR2_X1   g721(.A1(new_n187), .A2(G952), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n864), .A2(new_n887), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(new_n234), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n911), .A2(G210), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n547), .A2(new_n549), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n550), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT55), .Z(new_n915));
  OR2_X1    g729(.A1(KEYINPUT113), .A2(KEYINPUT114), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n912), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n911), .A2(KEYINPUT113), .A3(G210), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n909), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OR2_X1    g733(.A1(KEYINPUT114), .A2(KEYINPUT56), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n915), .B1(new_n912), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n908), .B1(new_n919), .B2(new_n921), .ZN(G51));
  INV_X1    g736(.A(new_n908), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n718), .B(KEYINPUT57), .Z(new_n924));
  AOI21_X1  g738(.A(new_n865), .B1(new_n864), .B2(new_n887), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n924), .B1(new_n888), .B2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n650), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n926), .A2(KEYINPUT115), .A3(new_n927), .ZN(new_n928));
  OR3_X1    g742(.A1(new_n910), .A2(new_n234), .A3(new_n752), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT115), .B1(new_n926), .B2(new_n927), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n923), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT116), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI211_X1 g748(.A(KEYINPUT116), .B(new_n923), .C1(new_n930), .C2(new_n931), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(G54));
  NAND3_X1  g750(.A1(new_n911), .A2(KEYINPUT58), .A3(G475), .ZN(new_n937));
  INV_X1    g751(.A(new_n406), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(new_n908), .ZN(G60));
  NAND2_X1  g755(.A1(new_n566), .A2(new_n567), .ZN(new_n942));
  NAND2_X1  g756(.A1(G478), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT59), .Z(new_n944));
  OAI21_X1  g758(.A(new_n942), .B1(new_n894), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(KEYINPUT117), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT117), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n947), .B(new_n942), .C1(new_n894), .C2(new_n944), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n888), .A2(new_n925), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n942), .A2(new_n944), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n908), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n946), .A2(new_n948), .A3(new_n951), .ZN(G63));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n953));
  NAND2_X1  g767(.A1(G217), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT118), .Z(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT60), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n910), .A2(new_n956), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n957), .A2(new_n230), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT119), .B1(new_n958), .B2(new_n923), .ZN(new_n959));
  OAI211_X1 g773(.A(KEYINPUT119), .B(new_n923), .C1(new_n957), .C2(new_n230), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n957), .A2(new_n602), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n953), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT120), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n958), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n958), .A2(new_n964), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n908), .A2(new_n953), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n966), .A2(new_n961), .A3(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n963), .B1(new_n965), .B2(new_n968), .ZN(G66));
  INV_X1    g783(.A(new_n515), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n187), .B1(new_n970), .B2(G224), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n890), .A2(new_n867), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n971), .B1(new_n972), .B2(new_n187), .ZN(new_n973));
  INV_X1    g787(.A(G898), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n913), .B1(new_n974), .B2(G953), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n973), .B(new_n975), .ZN(G69));
  NOR2_X1   g790(.A1(new_n378), .A2(new_n379), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n335), .B(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n728), .A2(new_n734), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT124), .ZN(new_n980));
  NOR4_X1   g794(.A1(new_n758), .A2(new_n759), .A3(new_n800), .A4(new_n875), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n769), .B2(new_n774), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n980), .A2(new_n762), .A3(new_n882), .A4(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n187), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n616), .A2(G953), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n985), .B(KEYINPUT123), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n978), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n643), .A2(new_n882), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(KEYINPUT62), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT62), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n643), .A2(new_n990), .A3(new_n882), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n830), .A2(new_n831), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n641), .A2(new_n760), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n348), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n775), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n762), .A2(new_n989), .A3(new_n991), .A4(new_n995), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(KEYINPUT121), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n187), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n987), .B1(new_n998), .B2(new_n978), .ZN(new_n999));
  OAI21_X1  g813(.A(G953), .B1(new_n439), .B2(new_n616), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n1000), .B1(new_n987), .B2(KEYINPUT122), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n999), .B(new_n1001), .Z(G72));
  NAND2_X1  g816(.A1(G472), .A2(G902), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT63), .Z(new_n1004));
  OAI21_X1  g818(.A(new_n1004), .B1(new_n997), .B2(new_n972), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n632), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n338), .A2(new_n311), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1007), .A2(new_n681), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1008), .A2(new_n1004), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT125), .Z(new_n1010));
  OAI21_X1  g824(.A(new_n1004), .B1(new_n983), .B2(new_n972), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n338), .A2(new_n315), .ZN(new_n1012));
  AOI22_X1  g826(.A1(new_n893), .A2(new_n1010), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1006), .A2(new_n1013), .A3(new_n923), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT126), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g830(.A1(new_n1006), .A2(KEYINPUT126), .A3(new_n923), .A4(new_n1013), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(G57));
endmodule


