

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  BUF_X1 U548 ( .A(n556), .Z(n557) );
  NAND2_X1 U549 ( .A1(n888), .A2(n516), .ZN(n751) );
  OR2_X1 U550 ( .A1(n750), .A2(n761), .ZN(n516) );
  AND2_X1 U551 ( .A1(n808), .A2(n798), .ZN(n517) );
  NAND2_X1 U552 ( .A1(n799), .A2(n517), .ZN(n518) );
  NOR2_X1 U553 ( .A1(n911), .A2(n706), .ZN(n693) );
  NOR2_X1 U554 ( .A1(G299), .A2(n700), .ZN(n697) );
  INV_X1 U555 ( .A(KEYINPUT90), .ZN(n672) );
  XNOR2_X1 U556 ( .A(n766), .B(n672), .ZN(n673) );
  NOR2_X1 U557 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U558 ( .A1(n673), .A2(n767), .ZN(n674) );
  INV_X1 U559 ( .A(n706), .ZN(n722) );
  NOR2_X1 U560 ( .A1(G651), .A2(n624), .ZN(n637) );
  INV_X1 U561 ( .A(KEYINPUT23), .ZN(n524) );
  OR2_X1 U562 ( .A1(n800), .A2(n518), .ZN(n815) );
  INV_X1 U563 ( .A(G2105), .ZN(n519) );
  NOR2_X1 U564 ( .A1(G2104), .A2(n519), .ZN(n1002) );
  NAND2_X1 U565 ( .A1(G125), .A2(n1002), .ZN(n521) );
  AND2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n1003) );
  NAND2_X1 U567 ( .A1(G113), .A2(n1003), .ZN(n520) );
  NAND2_X1 U568 ( .A1(n521), .A2(n520), .ZN(n529) );
  NOR2_X1 U569 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  XOR2_X2 U570 ( .A(KEYINPUT17), .B(n522), .Z(n1007) );
  NAND2_X1 U571 ( .A1(n1007), .A2(G137), .ZN(n527) );
  NAND2_X1 U572 ( .A1(n519), .A2(G2104), .ZN(n523) );
  XNOR2_X1 U573 ( .A(n523), .B(KEYINPUT65), .ZN(n556) );
  NAND2_X1 U574 ( .A1(G101), .A2(n556), .ZN(n525) );
  XNOR2_X1 U575 ( .A(n525), .B(n524), .ZN(n526) );
  NAND2_X1 U576 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U577 ( .A1(n529), .A2(n528), .ZN(G160) );
  XOR2_X1 U578 ( .A(KEYINPUT0), .B(G543), .Z(n624) );
  NAND2_X1 U579 ( .A1(n637), .A2(G53), .ZN(n531) );
  XOR2_X1 U580 ( .A(KEYINPUT66), .B(G651), .Z(n532) );
  NOR2_X1 U581 ( .A1(n624), .A2(n532), .ZN(n640) );
  NAND2_X1 U582 ( .A1(G78), .A2(n640), .ZN(n530) );
  NAND2_X1 U583 ( .A1(n531), .A2(n530), .ZN(n538) );
  NOR2_X1 U584 ( .A1(G651), .A2(G543), .ZN(n636) );
  NAND2_X1 U585 ( .A1(n636), .A2(G91), .ZN(n536) );
  NOR2_X1 U586 ( .A1(G543), .A2(n532), .ZN(n533) );
  XNOR2_X1 U587 ( .A(n533), .B(KEYINPUT1), .ZN(n534) );
  XNOR2_X1 U588 ( .A(KEYINPUT67), .B(n534), .ZN(n643) );
  NAND2_X1 U589 ( .A1(G65), .A2(n643), .ZN(n535) );
  NAND2_X1 U590 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U591 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U592 ( .A(n539), .B(KEYINPUT69), .ZN(G299) );
  NAND2_X1 U593 ( .A1(n636), .A2(G89), .ZN(n540) );
  XNOR2_X1 U594 ( .A(n540), .B(KEYINPUT4), .ZN(n542) );
  NAND2_X1 U595 ( .A1(G76), .A2(n640), .ZN(n541) );
  NAND2_X1 U596 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U597 ( .A(n543), .B(KEYINPUT5), .ZN(n548) );
  NAND2_X1 U598 ( .A1(n637), .A2(G51), .ZN(n545) );
  NAND2_X1 U599 ( .A1(G63), .A2(n643), .ZN(n544) );
  NAND2_X1 U600 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U601 ( .A(KEYINPUT6), .B(n546), .Z(n547) );
  NAND2_X1 U602 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U603 ( .A(n549), .B(KEYINPUT7), .Z(n887) );
  XNOR2_X1 U604 ( .A(n887), .B(KEYINPUT8), .ZN(G286) );
  NAND2_X1 U605 ( .A1(n636), .A2(G85), .ZN(n551) );
  NAND2_X1 U606 ( .A1(G60), .A2(n643), .ZN(n550) );
  NAND2_X1 U607 ( .A1(n551), .A2(n550), .ZN(n555) );
  NAND2_X1 U608 ( .A1(n637), .A2(G47), .ZN(n553) );
  NAND2_X1 U609 ( .A1(G72), .A2(n640), .ZN(n552) );
  NAND2_X1 U610 ( .A1(n553), .A2(n552), .ZN(n554) );
  OR2_X1 U611 ( .A1(n555), .A2(n554), .ZN(G290) );
  AND2_X1 U612 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U613 ( .A(G57), .ZN(G237) );
  INV_X1 U614 ( .A(G132), .ZN(G219) );
  INV_X1 U615 ( .A(G82), .ZN(G220) );
  INV_X1 U616 ( .A(G96), .ZN(G221) );
  NAND2_X1 U617 ( .A1(G138), .A2(n1007), .ZN(n559) );
  NAND2_X1 U618 ( .A1(G102), .A2(n557), .ZN(n558) );
  NAND2_X1 U619 ( .A1(n559), .A2(n558), .ZN(n563) );
  NAND2_X1 U620 ( .A1(G126), .A2(n1002), .ZN(n561) );
  NAND2_X1 U621 ( .A1(G114), .A2(n1003), .ZN(n560) );
  NAND2_X1 U622 ( .A1(n561), .A2(n560), .ZN(n562) );
  NOR2_X1 U623 ( .A1(n563), .A2(n562), .ZN(G164) );
  NAND2_X1 U624 ( .A1(G7), .A2(G661), .ZN(n564) );
  XNOR2_X1 U625 ( .A(n564), .B(KEYINPUT70), .ZN(n565) );
  XNOR2_X1 U626 ( .A(KEYINPUT10), .B(n565), .ZN(G223) );
  XNOR2_X1 U627 ( .A(KEYINPUT71), .B(G223), .ZN(n817) );
  NAND2_X1 U628 ( .A1(n817), .A2(G567), .ZN(n566) );
  XOR2_X1 U629 ( .A(KEYINPUT11), .B(n566), .Z(G234) );
  XOR2_X1 U630 ( .A(G860), .B(KEYINPUT74), .Z(n599) );
  XOR2_X1 U631 ( .A(KEYINPUT14), .B(KEYINPUT73), .Z(n568) );
  NAND2_X1 U632 ( .A1(G56), .A2(n643), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XOR2_X1 U634 ( .A(KEYINPUT72), .B(n569), .Z(n575) );
  NAND2_X1 U635 ( .A1(n636), .A2(G81), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(KEYINPUT12), .ZN(n572) );
  NAND2_X1 U637 ( .A1(G68), .A2(n640), .ZN(n571) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U639 ( .A(KEYINPUT13), .B(n573), .Z(n574) );
  NOR2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n637), .A2(G43), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n953) );
  OR2_X1 U643 ( .A1(n599), .A2(n953), .ZN(G153) );
  NAND2_X1 U644 ( .A1(n637), .A2(G52), .ZN(n579) );
  NAND2_X1 U645 ( .A1(G64), .A2(n643), .ZN(n578) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n585) );
  NAND2_X1 U647 ( .A1(G77), .A2(n640), .ZN(n580) );
  XNOR2_X1 U648 ( .A(n580), .B(KEYINPUT68), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G90), .A2(n636), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U651 ( .A(KEYINPUT9), .B(n583), .Z(n584) );
  NOR2_X1 U652 ( .A1(n585), .A2(n584), .ZN(G171) );
  INV_X1 U653 ( .A(G171), .ZN(G301) );
  NAND2_X1 U654 ( .A1(G868), .A2(G301), .ZN(n595) );
  NAND2_X1 U655 ( .A1(n636), .A2(G92), .ZN(n587) );
  NAND2_X1 U656 ( .A1(G66), .A2(n643), .ZN(n586) );
  NAND2_X1 U657 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U658 ( .A1(n637), .A2(G54), .ZN(n589) );
  NAND2_X1 U659 ( .A1(G79), .A2(n640), .ZN(n588) );
  NAND2_X1 U660 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U661 ( .A1(n591), .A2(n590), .ZN(n593) );
  XNOR2_X1 U662 ( .A(KEYINPUT75), .B(KEYINPUT15), .ZN(n592) );
  XOR2_X1 U663 ( .A(n593), .B(n592), .Z(n687) );
  INV_X1 U664 ( .A(G868), .ZN(n596) );
  NAND2_X1 U665 ( .A1(n687), .A2(n596), .ZN(n594) );
  NAND2_X1 U666 ( .A1(n595), .A2(n594), .ZN(G284) );
  NAND2_X1 U667 ( .A1(G286), .A2(G868), .ZN(n598) );
  NAND2_X1 U668 ( .A1(G299), .A2(n596), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n598), .A2(n597), .ZN(G297) );
  NAND2_X1 U670 ( .A1(n599), .A2(G559), .ZN(n600) );
  INV_X1 U671 ( .A(n687), .ZN(n954) );
  NAND2_X1 U672 ( .A1(n600), .A2(n954), .ZN(n601) );
  XNOR2_X1 U673 ( .A(n601), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U674 ( .A1(G868), .A2(n953), .ZN(n604) );
  NAND2_X1 U675 ( .A1(G868), .A2(n954), .ZN(n602) );
  NOR2_X1 U676 ( .A1(G559), .A2(n602), .ZN(n603) );
  NOR2_X1 U677 ( .A1(n604), .A2(n603), .ZN(G282) );
  NAND2_X1 U678 ( .A1(n1002), .A2(G123), .ZN(n605) );
  XNOR2_X1 U679 ( .A(n605), .B(KEYINPUT18), .ZN(n607) );
  NAND2_X1 U680 ( .A1(G111), .A2(n1003), .ZN(n606) );
  NAND2_X1 U681 ( .A1(n607), .A2(n606), .ZN(n611) );
  NAND2_X1 U682 ( .A1(G135), .A2(n1007), .ZN(n609) );
  NAND2_X1 U683 ( .A1(G99), .A2(n557), .ZN(n608) );
  NAND2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U685 ( .A1(n611), .A2(n610), .ZN(n991) );
  XNOR2_X1 U686 ( .A(n991), .B(G2096), .ZN(n612) );
  INV_X1 U687 ( .A(G2100), .ZN(n964) );
  NAND2_X1 U688 ( .A1(n612), .A2(n964), .ZN(G156) );
  NAND2_X1 U689 ( .A1(G559), .A2(n954), .ZN(n613) );
  XNOR2_X1 U690 ( .A(n613), .B(n953), .ZN(n653) );
  NOR2_X1 U691 ( .A1(n653), .A2(G860), .ZN(n622) );
  NAND2_X1 U692 ( .A1(G93), .A2(n636), .ZN(n615) );
  NAND2_X1 U693 ( .A1(G80), .A2(n640), .ZN(n614) );
  NAND2_X1 U694 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U695 ( .A(KEYINPUT76), .B(n616), .Z(n618) );
  NAND2_X1 U696 ( .A1(G67), .A2(n643), .ZN(n617) );
  NAND2_X1 U697 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U698 ( .A1(G55), .A2(n637), .ZN(n619) );
  XNOR2_X1 U699 ( .A(KEYINPUT77), .B(n619), .ZN(n620) );
  NOR2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n655) );
  INV_X1 U701 ( .A(n655), .ZN(n958) );
  XOR2_X1 U702 ( .A(n622), .B(n958), .Z(G145) );
  NAND2_X1 U703 ( .A1(G74), .A2(G651), .ZN(n623) );
  XNOR2_X1 U704 ( .A(n623), .B(KEYINPUT78), .ZN(n629) );
  NAND2_X1 U705 ( .A1(G49), .A2(n637), .ZN(n626) );
  NAND2_X1 U706 ( .A1(G87), .A2(n624), .ZN(n625) );
  NAND2_X1 U707 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U708 ( .A1(n643), .A2(n627), .ZN(n628) );
  NAND2_X1 U709 ( .A1(n629), .A2(n628), .ZN(G288) );
  NAND2_X1 U710 ( .A1(G88), .A2(n636), .ZN(n631) );
  NAND2_X1 U711 ( .A1(G75), .A2(n640), .ZN(n630) );
  NAND2_X1 U712 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U713 ( .A1(n637), .A2(G50), .ZN(n633) );
  NAND2_X1 U714 ( .A1(G62), .A2(n643), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U716 ( .A1(n635), .A2(n634), .ZN(G166) );
  INV_X1 U717 ( .A(G166), .ZN(G303) );
  NAND2_X1 U718 ( .A1(G86), .A2(n636), .ZN(n639) );
  NAND2_X1 U719 ( .A1(G48), .A2(n637), .ZN(n638) );
  NAND2_X1 U720 ( .A1(n639), .A2(n638), .ZN(n647) );
  NAND2_X1 U721 ( .A1(n640), .A2(G73), .ZN(n641) );
  XOR2_X1 U722 ( .A(KEYINPUT79), .B(n641), .Z(n642) );
  XNOR2_X1 U723 ( .A(n642), .B(KEYINPUT2), .ZN(n645) );
  NAND2_X1 U724 ( .A1(G61), .A2(n643), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n645), .A2(n644), .ZN(n646) );
  NOR2_X1 U726 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U727 ( .A(KEYINPUT80), .B(n648), .Z(G305) );
  XNOR2_X1 U728 ( .A(G288), .B(KEYINPUT19), .ZN(n650) );
  XOR2_X1 U729 ( .A(G303), .B(G305), .Z(n649) );
  XNOR2_X1 U730 ( .A(n650), .B(n649), .ZN(n651) );
  XOR2_X1 U731 ( .A(n651), .B(G290), .Z(n652) );
  XNOR2_X1 U732 ( .A(G299), .B(n652), .ZN(n957) );
  XNOR2_X1 U733 ( .A(n653), .B(n957), .ZN(n654) );
  NAND2_X1 U734 ( .A1(n654), .A2(G868), .ZN(n656) );
  XOR2_X1 U735 ( .A(n656), .B(n655), .Z(G295) );
  NAND2_X1 U736 ( .A1(G2084), .A2(G2078), .ZN(n657) );
  XOR2_X1 U737 ( .A(KEYINPUT20), .B(n657), .Z(n658) );
  NAND2_X1 U738 ( .A1(G2090), .A2(n658), .ZN(n660) );
  XOR2_X1 U739 ( .A(KEYINPUT21), .B(KEYINPUT81), .Z(n659) );
  XNOR2_X1 U740 ( .A(n660), .B(n659), .ZN(n661) );
  NAND2_X1 U741 ( .A1(G2072), .A2(n661), .ZN(G158) );
  XNOR2_X1 U742 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U743 ( .A1(G220), .A2(G219), .ZN(n662) );
  XOR2_X1 U744 ( .A(KEYINPUT22), .B(n662), .Z(n663) );
  NOR2_X1 U745 ( .A1(G218), .A2(n663), .ZN(n664) );
  XOR2_X1 U746 ( .A(KEYINPUT82), .B(n664), .Z(n665) );
  NOR2_X1 U747 ( .A1(G221), .A2(n665), .ZN(n666) );
  XNOR2_X1 U748 ( .A(KEYINPUT83), .B(n666), .ZN(n940) );
  NAND2_X1 U749 ( .A1(n940), .A2(G2106), .ZN(n670) );
  NAND2_X1 U750 ( .A1(G69), .A2(G120), .ZN(n667) );
  NOR2_X1 U751 ( .A1(G237), .A2(n667), .ZN(n668) );
  NAND2_X1 U752 ( .A1(G108), .A2(n668), .ZN(n941) );
  NAND2_X1 U753 ( .A1(n941), .A2(G567), .ZN(n669) );
  NAND2_X1 U754 ( .A1(n670), .A2(n669), .ZN(n1024) );
  NAND2_X1 U755 ( .A1(G483), .A2(G661), .ZN(n671) );
  NOR2_X1 U756 ( .A1(n1024), .A2(n671), .ZN(n819) );
  NAND2_X1 U757 ( .A1(n819), .A2(G36), .ZN(G176) );
  NAND2_X1 U758 ( .A1(G160), .A2(G40), .ZN(n766) );
  NOR2_X1 U759 ( .A1(G164), .A2(G1384), .ZN(n767) );
  XOR2_X2 U760 ( .A(n674), .B(KEYINPUT64), .Z(n706) );
  INV_X1 U761 ( .A(G1996), .ZN(n980) );
  NOR2_X1 U762 ( .A1(n722), .A2(n980), .ZN(n676) );
  INV_X1 U763 ( .A(KEYINPUT26), .ZN(n675) );
  NAND2_X1 U764 ( .A1(n676), .A2(n675), .ZN(n679) );
  INV_X1 U765 ( .A(n676), .ZN(n677) );
  NAND2_X1 U766 ( .A1(n677), .A2(KEYINPUT26), .ZN(n678) );
  NAND2_X1 U767 ( .A1(n679), .A2(n678), .ZN(n681) );
  NAND2_X1 U768 ( .A1(n722), .A2(G1341), .ZN(n680) );
  NAND2_X1 U769 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U770 ( .A1(n953), .A2(n682), .ZN(n689) );
  NAND2_X1 U771 ( .A1(G2067), .A2(n706), .ZN(n684) );
  NAND2_X1 U772 ( .A1(n722), .A2(G1348), .ZN(n683) );
  NAND2_X1 U773 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U774 ( .A(n685), .B(KEYINPUT94), .Z(n690) );
  INV_X1 U775 ( .A(n690), .ZN(n686) );
  NAND2_X1 U776 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U777 ( .A1(n689), .A2(n688), .ZN(n692) );
  NAND2_X1 U778 ( .A1(n690), .A2(n954), .ZN(n691) );
  NAND2_X1 U779 ( .A1(n692), .A2(n691), .ZN(n699) );
  XOR2_X1 U780 ( .A(G1956), .B(KEYINPUT92), .Z(n911) );
  XNOR2_X1 U781 ( .A(KEYINPUT93), .B(n693), .ZN(n696) );
  NAND2_X1 U782 ( .A1(G2072), .A2(n706), .ZN(n694) );
  XOR2_X1 U783 ( .A(KEYINPUT27), .B(n694), .Z(n695) );
  NAND2_X1 U784 ( .A1(n696), .A2(n695), .ZN(n700) );
  XOR2_X1 U785 ( .A(KEYINPUT95), .B(n697), .Z(n698) );
  NOR2_X1 U786 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U787 ( .A1(G299), .A2(n700), .ZN(n701) );
  XOR2_X1 U788 ( .A(KEYINPUT28), .B(n701), .Z(n702) );
  NOR2_X1 U789 ( .A1(n703), .A2(n702), .ZN(n705) );
  XNOR2_X1 U790 ( .A(KEYINPUT96), .B(KEYINPUT29), .ZN(n704) );
  XNOR2_X1 U791 ( .A(n705), .B(n704), .ZN(n710) );
  NOR2_X1 U792 ( .A1(G1961), .A2(n706), .ZN(n708) );
  XOR2_X1 U793 ( .A(G2078), .B(KEYINPUT25), .Z(n863) );
  NOR2_X1 U794 ( .A1(n722), .A2(n863), .ZN(n707) );
  NOR2_X1 U795 ( .A1(n708), .A2(n707), .ZN(n716) );
  OR2_X1 U796 ( .A1(G301), .A2(n716), .ZN(n709) );
  NAND2_X1 U797 ( .A1(n710), .A2(n709), .ZN(n721) );
  NAND2_X1 U798 ( .A1(n722), .A2(G8), .ZN(n761) );
  NOR2_X1 U799 ( .A1(G1966), .A2(n761), .ZN(n733) );
  NOR2_X1 U800 ( .A1(n722), .A2(G2084), .ZN(n711) );
  XOR2_X1 U801 ( .A(KEYINPUT91), .B(n711), .Z(n736) );
  INV_X1 U802 ( .A(n736), .ZN(n712) );
  NAND2_X1 U803 ( .A1(G8), .A2(n712), .ZN(n713) );
  NOR2_X1 U804 ( .A1(n733), .A2(n713), .ZN(n714) );
  XNOR2_X1 U805 ( .A(n714), .B(KEYINPUT30), .ZN(n715) );
  NAND2_X1 U806 ( .A1(n715), .A2(n887), .ZN(n718) );
  NAND2_X1 U807 ( .A1(n716), .A2(G301), .ZN(n717) );
  NAND2_X1 U808 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U809 ( .A(n719), .B(KEYINPUT31), .ZN(n720) );
  NAND2_X1 U810 ( .A1(n721), .A2(n720), .ZN(n731) );
  NAND2_X1 U811 ( .A1(n731), .A2(G286), .ZN(n727) );
  NOR2_X1 U812 ( .A1(n722), .A2(G2090), .ZN(n724) );
  NOR2_X1 U813 ( .A1(G1971), .A2(n761), .ZN(n723) );
  NOR2_X1 U814 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U815 ( .A1(n725), .A2(G303), .ZN(n726) );
  NAND2_X1 U816 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U817 ( .A(n728), .B(KEYINPUT98), .ZN(n729) );
  NAND2_X1 U818 ( .A1(n729), .A2(G8), .ZN(n730) );
  XNOR2_X1 U819 ( .A(KEYINPUT32), .B(n730), .ZN(n753) );
  INV_X1 U820 ( .A(KEYINPUT97), .ZN(n735) );
  INV_X1 U821 ( .A(n731), .ZN(n732) );
  XNOR2_X1 U822 ( .A(n735), .B(n734), .ZN(n738) );
  NAND2_X1 U823 ( .A1(G8), .A2(n736), .ZN(n737) );
  NAND2_X1 U824 ( .A1(n738), .A2(n737), .ZN(n754) );
  NAND2_X1 U825 ( .A1(G1976), .A2(G288), .ZN(n893) );
  INV_X1 U826 ( .A(n761), .ZN(n739) );
  NAND2_X1 U827 ( .A1(n893), .A2(n739), .ZN(n745) );
  INV_X1 U828 ( .A(n745), .ZN(n740) );
  AND2_X1 U829 ( .A1(n754), .A2(n740), .ZN(n741) );
  AND2_X1 U830 ( .A1(n753), .A2(n741), .ZN(n749) );
  NOR2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n895) );
  NOR2_X1 U832 ( .A1(G1971), .A2(G303), .ZN(n742) );
  XOR2_X1 U833 ( .A(n742), .B(KEYINPUT99), .Z(n743) );
  NOR2_X1 U834 ( .A1(n895), .A2(n743), .ZN(n744) );
  OR2_X1 U835 ( .A1(n745), .A2(n744), .ZN(n747) );
  INV_X1 U836 ( .A(KEYINPUT33), .ZN(n746) );
  NAND2_X1 U837 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U838 ( .A1(n749), .A2(n748), .ZN(n752) );
  XOR2_X1 U839 ( .A(G1981), .B(G305), .Z(n888) );
  NAND2_X1 U840 ( .A1(n895), .A2(KEYINPUT33), .ZN(n750) );
  NOR2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n765) );
  NAND2_X1 U842 ( .A1(n754), .A2(n753), .ZN(n757) );
  NOR2_X1 U843 ( .A1(G2090), .A2(G303), .ZN(n755) );
  NAND2_X1 U844 ( .A1(G8), .A2(n755), .ZN(n756) );
  NAND2_X1 U845 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U846 ( .A1(n758), .A2(n761), .ZN(n763) );
  NOR2_X1 U847 ( .A1(G1981), .A2(G305), .ZN(n759) );
  XOR2_X1 U848 ( .A(n759), .B(KEYINPUT24), .Z(n760) );
  OR2_X1 U849 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U850 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U851 ( .A1(n765), .A2(n764), .ZN(n800) );
  NOR2_X1 U852 ( .A1(n767), .A2(n766), .ZN(n813) );
  XNOR2_X1 U853 ( .A(KEYINPUT84), .B(G1986), .ZN(n768) );
  XNOR2_X1 U854 ( .A(n768), .B(G290), .ZN(n892) );
  NAND2_X1 U855 ( .A1(n813), .A2(n892), .ZN(n769) );
  XOR2_X1 U856 ( .A(KEYINPUT85), .B(n769), .Z(n799) );
  NAND2_X1 U857 ( .A1(G140), .A2(n1007), .ZN(n771) );
  NAND2_X1 U858 ( .A1(G104), .A2(n557), .ZN(n770) );
  NAND2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U860 ( .A(KEYINPUT34), .B(n772), .ZN(n777) );
  NAND2_X1 U861 ( .A1(G128), .A2(n1002), .ZN(n774) );
  NAND2_X1 U862 ( .A1(G116), .A2(n1003), .ZN(n773) );
  NAND2_X1 U863 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U864 ( .A(KEYINPUT35), .B(n775), .Z(n776) );
  NOR2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U866 ( .A(KEYINPUT36), .B(n778), .ZN(n1015) );
  XNOR2_X1 U867 ( .A(G2067), .B(KEYINPUT37), .ZN(n810) );
  NOR2_X1 U868 ( .A1(n1015), .A2(n810), .ZN(n842) );
  NAND2_X1 U869 ( .A1(n813), .A2(n842), .ZN(n808) );
  NAND2_X1 U870 ( .A1(n1003), .A2(G117), .ZN(n779) );
  XNOR2_X1 U871 ( .A(n779), .B(KEYINPUT86), .ZN(n781) );
  NAND2_X1 U872 ( .A1(G129), .A2(n1002), .ZN(n780) );
  NAND2_X1 U873 ( .A1(n781), .A2(n780), .ZN(n785) );
  NAND2_X1 U874 ( .A1(G105), .A2(n557), .ZN(n782) );
  XNOR2_X1 U875 ( .A(n782), .B(KEYINPUT38), .ZN(n783) );
  XNOR2_X1 U876 ( .A(n783), .B(KEYINPUT87), .ZN(n784) );
  NOR2_X1 U877 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U878 ( .A(n786), .B(KEYINPUT88), .ZN(n788) );
  NAND2_X1 U879 ( .A1(G141), .A2(n1007), .ZN(n787) );
  NAND2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n989) );
  AND2_X1 U881 ( .A1(n989), .A2(G1996), .ZN(n796) );
  NAND2_X1 U882 ( .A1(G131), .A2(n1007), .ZN(n790) );
  NAND2_X1 U883 ( .A1(G119), .A2(n1002), .ZN(n789) );
  NAND2_X1 U884 ( .A1(n790), .A2(n789), .ZN(n794) );
  NAND2_X1 U885 ( .A1(G95), .A2(n557), .ZN(n792) );
  NAND2_X1 U886 ( .A1(G107), .A2(n1003), .ZN(n791) );
  NAND2_X1 U887 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U888 ( .A1(n794), .A2(n793), .ZN(n990) );
  INV_X1 U889 ( .A(G1991), .ZN(n977) );
  NOR2_X1 U890 ( .A1(n990), .A2(n977), .ZN(n795) );
  NOR2_X1 U891 ( .A1(n796), .A2(n795), .ZN(n854) );
  INV_X1 U892 ( .A(n813), .ZN(n797) );
  NOR2_X1 U893 ( .A1(n854), .A2(n797), .ZN(n805) );
  XNOR2_X1 U894 ( .A(KEYINPUT89), .B(n805), .ZN(n798) );
  NOR2_X1 U895 ( .A1(n989), .A2(G1996), .ZN(n801) );
  XNOR2_X1 U896 ( .A(n801), .B(KEYINPUT100), .ZN(n851) );
  AND2_X1 U897 ( .A1(n977), .A2(n990), .ZN(n802) );
  XOR2_X1 U898 ( .A(KEYINPUT101), .B(n802), .Z(n847) );
  NOR2_X1 U899 ( .A1(G1986), .A2(G290), .ZN(n803) );
  NOR2_X1 U900 ( .A1(n847), .A2(n803), .ZN(n804) );
  NOR2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n806) );
  NOR2_X1 U902 ( .A1(n851), .A2(n806), .ZN(n807) );
  XNOR2_X1 U903 ( .A(KEYINPUT39), .B(n807), .ZN(n809) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U905 ( .A1(n1015), .A2(n810), .ZN(n844) );
  NAND2_X1 U906 ( .A1(n811), .A2(n844), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U909 ( .A(n816), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U910 ( .A(n887), .ZN(G168) );
  NAND2_X1 U911 ( .A1(G2106), .A2(n817), .ZN(G217) );
  AND2_X1 U912 ( .A1(G15), .A2(G2), .ZN(n818) );
  NAND2_X1 U913 ( .A1(G661), .A2(n818), .ZN(G259) );
  NAND2_X1 U914 ( .A1(G3), .A2(G1), .ZN(n820) );
  NAND2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n821) );
  XOR2_X1 U916 ( .A(KEYINPUT105), .B(n821), .Z(G188) );
  NAND2_X1 U918 ( .A1(G100), .A2(n557), .ZN(n823) );
  NAND2_X1 U919 ( .A1(G112), .A2(n1003), .ZN(n822) );
  NAND2_X1 U920 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U921 ( .A(n824), .B(KEYINPUT111), .ZN(n826) );
  NAND2_X1 U922 ( .A1(G136), .A2(n1007), .ZN(n825) );
  NAND2_X1 U923 ( .A1(n826), .A2(n825), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n1002), .A2(G124), .ZN(n827) );
  XOR2_X1 U925 ( .A(KEYINPUT44), .B(n827), .Z(n828) );
  NOR2_X1 U926 ( .A1(n829), .A2(n828), .ZN(G162) );
  NAND2_X1 U927 ( .A1(G139), .A2(n1007), .ZN(n831) );
  NAND2_X1 U928 ( .A1(G103), .A2(n557), .ZN(n830) );
  NAND2_X1 U929 ( .A1(n831), .A2(n830), .ZN(n837) );
  NAND2_X1 U930 ( .A1(G127), .A2(n1002), .ZN(n833) );
  NAND2_X1 U931 ( .A1(G115), .A2(n1003), .ZN(n832) );
  NAND2_X1 U932 ( .A1(n833), .A2(n832), .ZN(n834) );
  XOR2_X1 U933 ( .A(KEYINPUT114), .B(n834), .Z(n835) );
  XNOR2_X1 U934 ( .A(KEYINPUT47), .B(n835), .ZN(n836) );
  NOR2_X1 U935 ( .A1(n837), .A2(n836), .ZN(n997) );
  XOR2_X1 U936 ( .A(G2072), .B(n997), .Z(n839) );
  XOR2_X1 U937 ( .A(G164), .B(G2078), .Z(n838) );
  NOR2_X1 U938 ( .A1(n839), .A2(n838), .ZN(n840) );
  XOR2_X1 U939 ( .A(KEYINPUT50), .B(n840), .Z(n841) );
  NOR2_X1 U940 ( .A1(n842), .A2(n841), .ZN(n849) );
  XOR2_X1 U941 ( .A(G2084), .B(G160), .Z(n843) );
  NOR2_X1 U942 ( .A1(n991), .A2(n843), .ZN(n845) );
  NAND2_X1 U943 ( .A1(n845), .A2(n844), .ZN(n846) );
  NOR2_X1 U944 ( .A1(n847), .A2(n846), .ZN(n848) );
  NAND2_X1 U945 ( .A1(n849), .A2(n848), .ZN(n856) );
  XOR2_X1 U946 ( .A(G2090), .B(G162), .Z(n850) );
  NOR2_X1 U947 ( .A1(n851), .A2(n850), .ZN(n852) );
  XOR2_X1 U948 ( .A(KEYINPUT51), .B(n852), .Z(n853) );
  NAND2_X1 U949 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U950 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U951 ( .A(KEYINPUT52), .B(n857), .ZN(n858) );
  INV_X1 U952 ( .A(KEYINPUT55), .ZN(n882) );
  NAND2_X1 U953 ( .A1(n858), .A2(n882), .ZN(n859) );
  NAND2_X1 U954 ( .A1(n859), .A2(G29), .ZN(n860) );
  XNOR2_X1 U955 ( .A(KEYINPUT118), .B(n860), .ZN(n861) );
  NAND2_X1 U956 ( .A1(n861), .A2(G11), .ZN(n886) );
  XNOR2_X1 U957 ( .A(G2090), .B(G35), .ZN(n877) );
  XOR2_X1 U958 ( .A(G32), .B(G1996), .Z(n870) );
  XOR2_X1 U959 ( .A(G2072), .B(G33), .Z(n865) );
  XOR2_X1 U960 ( .A(KEYINPUT120), .B(G27), .Z(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n864) );
  NAND2_X1 U962 ( .A1(n865), .A2(n864), .ZN(n868) );
  XOR2_X1 U963 ( .A(KEYINPUT119), .B(G2067), .Z(n866) );
  XNOR2_X1 U964 ( .A(G26), .B(n866), .ZN(n867) );
  NOR2_X1 U965 ( .A1(n868), .A2(n867), .ZN(n869) );
  NAND2_X1 U966 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U967 ( .A(KEYINPUT121), .B(n871), .ZN(n872) );
  NAND2_X1 U968 ( .A1(n872), .A2(G28), .ZN(n874) );
  XOR2_X1 U969 ( .A(G25), .B(n977), .Z(n873) );
  NOR2_X1 U970 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U971 ( .A(KEYINPUT53), .B(n875), .ZN(n876) );
  NOR2_X1 U972 ( .A1(n877), .A2(n876), .ZN(n880) );
  XOR2_X1 U973 ( .A(G2084), .B(G34), .Z(n878) );
  XNOR2_X1 U974 ( .A(KEYINPUT54), .B(n878), .ZN(n879) );
  NAND2_X1 U975 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U976 ( .A(n882), .B(n881), .Z(n883) );
  NOR2_X1 U977 ( .A1(G29), .A2(n883), .ZN(n884) );
  XNOR2_X1 U978 ( .A(KEYINPUT122), .B(n884), .ZN(n885) );
  NOR2_X1 U979 ( .A1(n886), .A2(n885), .ZN(n938) );
  XOR2_X1 U980 ( .A(G1966), .B(n887), .Z(n889) );
  NAND2_X1 U981 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U982 ( .A(KEYINPUT57), .B(n890), .Z(n908) );
  XNOR2_X1 U983 ( .A(G1341), .B(n953), .ZN(n891) );
  NOR2_X1 U984 ( .A1(n892), .A2(n891), .ZN(n899) );
  XOR2_X1 U985 ( .A(G303), .B(G1971), .Z(n894) );
  NAND2_X1 U986 ( .A1(n894), .A2(n893), .ZN(n896) );
  NOR2_X1 U987 ( .A1(n896), .A2(n895), .ZN(n897) );
  XOR2_X1 U988 ( .A(KEYINPUT123), .B(n897), .Z(n898) );
  NAND2_X1 U989 ( .A1(n899), .A2(n898), .ZN(n905) );
  XOR2_X1 U990 ( .A(G301), .B(G1961), .Z(n903) );
  XOR2_X1 U991 ( .A(n954), .B(G1348), .Z(n901) );
  XNOR2_X1 U992 ( .A(G299), .B(G1956), .ZN(n900) );
  NOR2_X1 U993 ( .A1(n901), .A2(n900), .ZN(n902) );
  NAND2_X1 U994 ( .A1(n903), .A2(n902), .ZN(n904) );
  NOR2_X1 U995 ( .A1(n905), .A2(n904), .ZN(n906) );
  XOR2_X1 U996 ( .A(KEYINPUT124), .B(n906), .Z(n907) );
  NOR2_X1 U997 ( .A1(n908), .A2(n907), .ZN(n910) );
  XOR2_X1 U998 ( .A(KEYINPUT56), .B(G16), .Z(n909) );
  NOR2_X1 U999 ( .A1(n910), .A2(n909), .ZN(n935) );
  XNOR2_X1 U1000 ( .A(n911), .B(G20), .ZN(n915) );
  XNOR2_X1 U1001 ( .A(G1341), .B(G19), .ZN(n913) );
  XNOR2_X1 U1002 ( .A(G1981), .B(G6), .ZN(n912) );
  NOR2_X1 U1003 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1004 ( .A1(n915), .A2(n914), .ZN(n918) );
  XOR2_X1 U1005 ( .A(KEYINPUT59), .B(G1348), .Z(n916) );
  XNOR2_X1 U1006 ( .A(G4), .B(n916), .ZN(n917) );
  NOR2_X1 U1007 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1008 ( .A(KEYINPUT60), .B(n919), .ZN(n923) );
  XNOR2_X1 U1009 ( .A(G1966), .B(G21), .ZN(n921) );
  XNOR2_X1 U1010 ( .A(G1961), .B(G5), .ZN(n920) );
  NOR2_X1 U1011 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1012 ( .A1(n923), .A2(n922), .ZN(n930) );
  XNOR2_X1 U1013 ( .A(G1986), .B(G24), .ZN(n925) );
  XNOR2_X1 U1014 ( .A(G1971), .B(G22), .ZN(n924) );
  NOR2_X1 U1015 ( .A1(n925), .A2(n924), .ZN(n927) );
  XOR2_X1 U1016 ( .A(G1976), .B(G23), .Z(n926) );
  NAND2_X1 U1017 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1018 ( .A(KEYINPUT58), .B(n928), .ZN(n929) );
  NOR2_X1 U1019 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1020 ( .A(KEYINPUT61), .B(n931), .Z(n933) );
  XOR2_X1 U1021 ( .A(G16), .B(KEYINPUT125), .Z(n932) );
  NOR2_X1 U1022 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1023 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1024 ( .A(n936), .B(KEYINPUT126), .ZN(n937) );
  NAND2_X1 U1025 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1026 ( .A(KEYINPUT62), .B(n939), .Z(G311) );
  XNOR2_X1 U1027 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1028 ( .A(G120), .ZN(G236) );
  INV_X1 U1029 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1030 ( .A1(n941), .A2(n940), .ZN(G325) );
  INV_X1 U1031 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U1032 ( .A(G2446), .B(G1348), .ZN(n950) );
  XNOR2_X1 U1033 ( .A(G2430), .B(G2451), .ZN(n948) );
  XOR2_X1 U1034 ( .A(G2454), .B(G2427), .Z(n943) );
  XNOR2_X1 U1035 ( .A(KEYINPUT102), .B(G2435), .ZN(n942) );
  XNOR2_X1 U1036 ( .A(n943), .B(n942), .ZN(n944) );
  XOR2_X1 U1037 ( .A(n944), .B(G2438), .Z(n946) );
  XNOR2_X1 U1038 ( .A(G1341), .B(G2443), .ZN(n945) );
  XNOR2_X1 U1039 ( .A(n946), .B(n945), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(n948), .B(n947), .ZN(n949) );
  XNOR2_X1 U1041 ( .A(n950), .B(n949), .ZN(n951) );
  NAND2_X1 U1042 ( .A1(n951), .A2(G14), .ZN(n952) );
  XOR2_X1 U1043 ( .A(KEYINPUT103), .B(n952), .Z(n1020) );
  XOR2_X1 U1044 ( .A(KEYINPUT104), .B(n1020), .Z(G401) );
  XNOR2_X1 U1045 ( .A(n953), .B(KEYINPUT116), .ZN(n956) );
  XOR2_X1 U1046 ( .A(G301), .B(n954), .Z(n955) );
  XNOR2_X1 U1047 ( .A(n956), .B(n955), .ZN(n961) );
  XOR2_X1 U1048 ( .A(n958), .B(n957), .Z(n959) );
  XOR2_X1 U1049 ( .A(G286), .B(n959), .Z(n960) );
  XNOR2_X1 U1050 ( .A(n961), .B(n960), .ZN(n962) );
  NOR2_X1 U1051 ( .A1(G37), .A2(n962), .ZN(n963) );
  XOR2_X1 U1052 ( .A(KEYINPUT117), .B(n963), .Z(G397) );
  XNOR2_X1 U1053 ( .A(KEYINPUT43), .B(n964), .ZN(n966) );
  XNOR2_X1 U1054 ( .A(G2090), .B(G2678), .ZN(n965) );
  XNOR2_X1 U1055 ( .A(n966), .B(n965), .ZN(n970) );
  XOR2_X1 U1056 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n968) );
  XNOR2_X1 U1057 ( .A(G2067), .B(KEYINPUT42), .ZN(n967) );
  XNOR2_X1 U1058 ( .A(n968), .B(n967), .ZN(n969) );
  XOR2_X1 U1059 ( .A(n970), .B(n969), .Z(n972) );
  XNOR2_X1 U1060 ( .A(G2072), .B(G2096), .ZN(n971) );
  XNOR2_X1 U1061 ( .A(n972), .B(n971), .ZN(n974) );
  XOR2_X1 U1062 ( .A(G2084), .B(G2078), .Z(n973) );
  XNOR2_X1 U1063 ( .A(n974), .B(n973), .ZN(G227) );
  XOR2_X1 U1064 ( .A(KEYINPUT108), .B(G1976), .Z(n976) );
  XNOR2_X1 U1065 ( .A(G1961), .B(G1956), .ZN(n975) );
  XNOR2_X1 U1066 ( .A(n976), .B(n975), .ZN(n988) );
  XOR2_X1 U1067 ( .A(G2474), .B(KEYINPUT41), .Z(n979) );
  XOR2_X1 U1068 ( .A(n977), .B(G1966), .Z(n978) );
  XNOR2_X1 U1069 ( .A(n979), .B(n978), .ZN(n984) );
  XOR2_X1 U1070 ( .A(KEYINPUT109), .B(G1981), .Z(n982) );
  XOR2_X1 U1071 ( .A(n980), .B(G1971), .Z(n981) );
  XNOR2_X1 U1072 ( .A(n982), .B(n981), .ZN(n983) );
  XOR2_X1 U1073 ( .A(n984), .B(n983), .Z(n986) );
  XNOR2_X1 U1074 ( .A(G1986), .B(KEYINPUT110), .ZN(n985) );
  XNOR2_X1 U1075 ( .A(n986), .B(n985), .ZN(n987) );
  XNOR2_X1 U1076 ( .A(n988), .B(n987), .ZN(G229) );
  XOR2_X1 U1077 ( .A(n990), .B(n989), .Z(n992) );
  XNOR2_X1 U1078 ( .A(n992), .B(n991), .ZN(n996) );
  XOR2_X1 U1079 ( .A(KEYINPUT113), .B(KEYINPUT115), .Z(n994) );
  XNOR2_X1 U1080 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(n994), .B(n993), .ZN(n995) );
  XOR2_X1 U1082 ( .A(n996), .B(n995), .Z(n1001) );
  XNOR2_X1 U1083 ( .A(G160), .B(G162), .ZN(n998) );
  XNOR2_X1 U1084 ( .A(n998), .B(n997), .ZN(n999) );
  XNOR2_X1 U1085 ( .A(G164), .B(n999), .ZN(n1000) );
  XNOR2_X1 U1086 ( .A(n1001), .B(n1000), .ZN(n1014) );
  NAND2_X1 U1087 ( .A1(G130), .A2(n1002), .ZN(n1005) );
  NAND2_X1 U1088 ( .A1(G118), .A2(n1003), .ZN(n1004) );
  NAND2_X1 U1089 ( .A1(n1005), .A2(n1004), .ZN(n1012) );
  NAND2_X1 U1090 ( .A1(n557), .A2(G106), .ZN(n1006) );
  XNOR2_X1 U1091 ( .A(n1006), .B(KEYINPUT112), .ZN(n1009) );
  NAND2_X1 U1092 ( .A1(G142), .A2(n1007), .ZN(n1008) );
  NAND2_X1 U1093 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1094 ( .A(n1010), .B(KEYINPUT45), .Z(n1011) );
  NOR2_X1 U1095 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1096 ( .A(n1014), .B(n1013), .Z(n1016) );
  XOR2_X1 U1097 ( .A(n1016), .B(n1015), .Z(n1017) );
  NOR2_X1 U1098 ( .A1(G37), .A2(n1017), .ZN(G395) );
  NOR2_X1 U1099 ( .A1(G227), .A2(G229), .ZN(n1018) );
  XOR2_X1 U1100 ( .A(KEYINPUT49), .B(n1018), .Z(n1019) );
  NAND2_X1 U1101 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1102 ( .A1(G397), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1103 ( .A1(G395), .A2(n1024), .ZN(n1022) );
  NAND2_X1 U1104 ( .A1(n1023), .A2(n1022), .ZN(G225) );
  INV_X1 U1105 ( .A(G225), .ZN(G308) );
  INV_X1 U1106 ( .A(n1024), .ZN(G319) );
  INV_X1 U1107 ( .A(G108), .ZN(G238) );
endmodule

