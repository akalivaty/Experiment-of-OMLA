//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962;
  INV_X1    g000(.A(G140), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G125), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(KEYINPUT16), .ZN(new_n189));
  INV_X1    g003(.A(G125), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n187), .B1(new_n190), .B2(KEYINPUT73), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT73), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(G125), .A3(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n189), .B1(new_n194), .B2(KEYINPUT16), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT74), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n190), .A2(G140), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n188), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n197), .B1(new_n200), .B2(new_n201), .ZN(new_n202));
  NOR3_X1   g016(.A1(new_n199), .A2(KEYINPUT74), .A3(G146), .ZN(new_n203));
  OR2_X1    g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G128), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G119), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(G128), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(G119), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n208), .B(KEYINPUT72), .ZN(new_n209));
  XOR2_X1   g023(.A(KEYINPUT24), .B(G110), .Z(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n208), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT23), .B1(new_n205), .B2(G119), .ZN(new_n215));
  NOR3_X1   g029(.A1(new_n214), .A2(G110), .A3(new_n215), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n196), .B(new_n204), .C1(new_n212), .C2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n195), .B(new_n201), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(G110), .B1(new_n214), .B2(new_n215), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n219), .B(new_n220), .C1(new_n211), .C2(new_n209), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G953), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(G221), .A3(G234), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n224), .B(KEYINPUT22), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n225), .B(G137), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n222), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n217), .A2(new_n221), .A3(new_n226), .ZN(new_n229));
  INV_X1    g043(.A(G902), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT25), .ZN(new_n232));
  INV_X1    g046(.A(G217), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n233), .B1(G234), .B2(new_n230), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT25), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n228), .A2(new_n229), .A3(new_n235), .A4(new_n230), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n232), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n228), .A2(new_n229), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n234), .A2(G902), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AND2_X1   g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G472), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT11), .ZN(new_n243));
  INV_X1    g057(.A(G134), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n243), .B1(new_n244), .B2(G137), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(G137), .ZN(new_n246));
  INV_X1    g060(.A(G137), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT11), .A3(G134), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n245), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n249), .A2(G131), .ZN(new_n250));
  INV_X1    g064(.A(G131), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n245), .A2(new_n248), .A3(new_n251), .A4(new_n246), .ZN(new_n252));
  OR2_X1    g066(.A1(new_n252), .A2(KEYINPUT64), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(KEYINPUT64), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n250), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n201), .A2(G143), .ZN(new_n256));
  INV_X1    g070(.A(G143), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G146), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n259), .B1(KEYINPUT0), .B2(G128), .ZN(new_n260));
  OR2_X1    g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  NAND2_X1  g075(.A1(KEYINPUT0), .A2(G128), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n256), .A2(new_n258), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT65), .B1(new_n255), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n249), .A2(G131), .ZN(new_n266));
  AND2_X1   g080(.A1(new_n252), .A2(KEYINPUT64), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n252), .A2(KEYINPUT64), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n264), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT65), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT1), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n273), .B1(G143), .B2(new_n201), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n259), .B1(new_n207), .B2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n256), .A2(new_n258), .A3(new_n273), .A4(G128), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n246), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n244), .A2(G137), .ZN(new_n279));
  OAI21_X1  g093(.A(G131), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n277), .B(new_n280), .C1(new_n267), .C2(new_n268), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT67), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n253), .A2(new_n254), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n284), .A2(KEYINPUT67), .A3(new_n277), .A4(new_n280), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n265), .A2(new_n272), .A3(new_n283), .A4(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT30), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  XOR2_X1   g102(.A(G116), .B(G119), .Z(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT2), .B(G113), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n289), .B(new_n290), .ZN(new_n291));
  OAI211_X1 g105(.A(new_n281), .B(KEYINPUT30), .C1(new_n255), .C2(new_n264), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n288), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT31), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n269), .A2(new_n270), .ZN(new_n295));
  INV_X1    g109(.A(new_n291), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n296), .A3(new_n281), .ZN(new_n297));
  XOR2_X1   g111(.A(KEYINPUT26), .B(G101), .Z(new_n298));
  INV_X1    g112(.A(G237), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(new_n223), .A3(G210), .ZN(new_n300));
  XNOR2_X1  g114(.A(new_n298), .B(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n301), .B(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n293), .A2(new_n294), .A3(new_n297), .A4(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n286), .A2(new_n291), .ZN(new_n306));
  INV_X1    g120(.A(new_n297), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT28), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT28), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n297), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n306), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n303), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n305), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n292), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n314), .B1(new_n286), .B2(new_n287), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n307), .B1(new_n315), .B2(new_n291), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n294), .B1(new_n316), .B2(new_n304), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n242), .B(new_n230), .C1(new_n313), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT32), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n293), .A2(new_n297), .A3(new_n304), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT31), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n321), .A2(new_n305), .A3(new_n312), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT32), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n322), .A2(new_n323), .A3(new_n242), .A4(new_n230), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT69), .B1(new_n316), .B2(new_n304), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n306), .A2(new_n308), .A3(new_n310), .ZN(new_n327));
  AOI21_X1  g141(.A(KEYINPUT29), .B1(new_n327), .B2(new_n304), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT69), .ZN(new_n329));
  AOI211_X1 g143(.A(new_n296), .B(new_n314), .C1(new_n286), .C2(new_n287), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n329), .B(new_n303), .C1(new_n330), .C2(new_n307), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n326), .A2(new_n328), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n296), .B1(new_n295), .B2(new_n281), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT28), .B1(new_n307), .B2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n297), .A2(KEYINPUT70), .A3(new_n309), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT70), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n310), .A2(new_n336), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n304), .A2(KEYINPUT29), .ZN(new_n339));
  AOI21_X1  g153(.A(G902), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n332), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(KEYINPUT71), .B1(new_n341), .B2(G472), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT71), .ZN(new_n343));
  AOI211_X1 g157(.A(new_n343), .B(new_n242), .C1(new_n332), .C2(new_n340), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n325), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G104), .ZN(new_n346));
  INV_X1    g160(.A(G107), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT76), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G107), .ZN(new_n350));
  AOI211_X1 g164(.A(KEYINPUT3), .B(new_n346), .C1(new_n348), .C2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT3), .B1(new_n346), .B2(G107), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n346), .A2(G107), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(G101), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n348), .A2(new_n350), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(G104), .ZN(new_n358));
  INV_X1    g172(.A(G101), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n358), .B(new_n359), .C1(new_n353), .C2(new_n352), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n355), .A2(new_n360), .A3(KEYINPUT4), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT4), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n362), .B(G101), .C1(new_n351), .C2(new_n354), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n270), .A3(new_n363), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n356), .A2(G104), .ZN(new_n365));
  OAI21_X1  g179(.A(G101), .B1(new_n365), .B2(new_n353), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n259), .B1(new_n274), .B2(new_n205), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n276), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n360), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n360), .A2(new_n366), .A3(KEYINPUT10), .A4(new_n277), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n364), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n269), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n364), .A2(new_n371), .A3(new_n255), .A4(new_n372), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g190(.A(G110), .B(G140), .ZN(new_n377));
  AND2_X1   g191(.A1(new_n223), .A2(G227), .ZN(new_n378));
  XOR2_X1   g192(.A(new_n377), .B(new_n378), .Z(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT78), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT78), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n376), .A2(new_n383), .A3(new_n380), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n375), .A2(new_n379), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n360), .A2(new_n366), .ZN(new_n387));
  INV_X1    g201(.A(new_n277), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n255), .B1(new_n389), .B2(new_n369), .ZN(new_n390));
  AND2_X1   g204(.A1(new_n390), .A2(KEYINPUT12), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(KEYINPUT12), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n386), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n382), .A2(new_n384), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G469), .ZN(new_n395));
  OR2_X1    g209(.A1(new_n395), .A2(KEYINPUT77), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(KEYINPUT77), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n394), .A2(new_n230), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n375), .B1(new_n391), .B2(new_n392), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n380), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n386), .A2(new_n374), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n230), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G469), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  XOR2_X1   g219(.A(KEYINPUT9), .B(G234), .Z(new_n406));
  XNOR2_X1  g220(.A(new_n406), .B(KEYINPUT75), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G221), .B1(new_n408), .B2(G902), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(G214), .B1(G237), .B2(G902), .ZN(new_n411));
  INV_X1    g225(.A(G952), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(G953), .ZN(new_n413));
  NAND2_X1  g227(.A1(G234), .A2(G237), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(KEYINPUT95), .ZN(new_n416));
  XOR2_X1   g230(.A(KEYINPUT21), .B(G898), .Z(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(G902), .A3(G953), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n416), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  XOR2_X1   g233(.A(G110), .B(G122), .Z(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n361), .A2(new_n291), .A3(new_n363), .ZN(new_n422));
  INV_X1    g236(.A(G113), .ZN(new_n423));
  XNOR2_X1  g237(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n424));
  INV_X1    g238(.A(G116), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(G119), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n423), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n427), .B1(new_n289), .B2(new_n424), .ZN(new_n428));
  OR2_X1    g242(.A1(new_n289), .A2(new_n290), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n360), .A2(new_n428), .A3(new_n366), .A4(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n421), .B1(new_n422), .B2(new_n430), .ZN(new_n431));
  OR2_X1    g245(.A1(new_n431), .A2(KEYINPUT6), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n422), .A2(new_n430), .A3(new_n421), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT80), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT80), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n422), .A2(new_n435), .A3(new_n430), .A4(new_n421), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n431), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT6), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n432), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n388), .A2(G125), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n264), .A2(new_n190), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n223), .A2(G224), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n443), .B(KEYINPUT81), .ZN(new_n444));
  XOR2_X1   g258(.A(new_n442), .B(new_n444), .Z(new_n445));
  NAND2_X1  g259(.A1(new_n439), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G210), .B1(G237), .B2(G902), .ZN(new_n447));
  XOR2_X1   g261(.A(KEYINPUT82), .B(KEYINPUT8), .Z(new_n448));
  XNOR2_X1  g262(.A(new_n420), .B(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n428), .A2(new_n429), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n387), .A2(new_n450), .ZN(new_n451));
  XOR2_X1   g265(.A(new_n451), .B(KEYINPUT83), .Z(new_n452));
  INV_X1    g266(.A(KEYINPUT5), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n427), .B1(new_n453), .B2(new_n289), .ZN(new_n454));
  AND4_X1   g268(.A1(new_n429), .A2(new_n360), .A3(new_n366), .A4(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n449), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n444), .A2(KEYINPUT7), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n440), .B2(new_n441), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n442), .A2(KEYINPUT7), .A3(new_n444), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n434), .A2(new_n436), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(G902), .B1(new_n456), .B2(new_n460), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n446), .A2(new_n447), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n447), .B1(new_n446), .B2(new_n461), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n411), .B(new_n419), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n410), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G478), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT94), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n467), .A2(KEYINPUT15), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(KEYINPUT15), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n466), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NOR3_X1   g286(.A1(new_n408), .A2(new_n233), .A3(G953), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(KEYINPUT88), .B1(new_n205), .B2(G143), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT88), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(new_n257), .A3(G128), .ZN(new_n477));
  AND2_X1   g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT89), .ZN(new_n479));
  AND2_X1   g293(.A1(KEYINPUT66), .A2(G128), .ZN(new_n480));
  NOR2_X1   g294(.A1(KEYINPUT66), .A2(G128), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n479), .B(G143), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(G143), .B1(new_n480), .B2(new_n481), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT89), .ZN(new_n484));
  AOI211_X1 g298(.A(KEYINPUT90), .B(new_n478), .C1(new_n482), .C2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT90), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n484), .A2(new_n482), .ZN(new_n487));
  INV_X1    g301(.A(new_n478), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n244), .B1(new_n485), .B2(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n478), .B(KEYINPUT13), .ZN(new_n491));
  INV_X1    g305(.A(new_n487), .ZN(new_n492));
  OAI21_X1  g306(.A(G134), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n425), .A2(G122), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n425), .A2(G122), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(new_n348), .A3(new_n350), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n356), .A2(new_n495), .A3(new_n496), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n490), .A2(new_n493), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT91), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT91), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n490), .A2(new_n503), .A3(new_n493), .A4(new_n500), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT93), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n494), .B1(KEYINPUT14), .B2(new_n496), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n507), .B(KEYINPUT92), .C1(KEYINPUT14), .C2(new_n496), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n508), .B(G107), .C1(KEYINPUT92), .C2(new_n507), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n479), .B1(new_n207), .B2(G143), .ZN(new_n510));
  INV_X1    g324(.A(new_n482), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n488), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT90), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n487), .A2(new_n486), .A3(new_n488), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n515), .A2(new_n244), .ZN(new_n516));
  AOI21_X1  g330(.A(G134), .B1(new_n513), .B2(new_n514), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n499), .B(new_n509), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n505), .A2(new_n506), .A3(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n506), .B1(new_n505), .B2(new_n518), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n474), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n500), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n522), .B1(new_n515), .B2(new_n244), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n503), .B1(new_n523), .B2(new_n493), .ZN(new_n524));
  INV_X1    g338(.A(new_n504), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n518), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT93), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n505), .A2(new_n506), .A3(new_n518), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(new_n473), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n521), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n472), .B1(new_n530), .B2(new_n230), .ZN(new_n531));
  AOI211_X1 g345(.A(G902), .B(new_n471), .C1(new_n521), .C2(new_n529), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT86), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n194), .A2(KEYINPUT19), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n534), .B1(KEYINPUT19), .B2(new_n200), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n201), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n536), .A2(new_n196), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n299), .A2(new_n223), .A3(G214), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n257), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n299), .A2(new_n223), .A3(G143), .A4(G214), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(G131), .ZN(new_n542));
  OR3_X1    g356(.A1(new_n194), .A2(KEYINPUT84), .A3(new_n201), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT84), .B1(new_n194), .B2(new_n201), .ZN(new_n544));
  OAI211_X1 g358(.A(new_n543), .B(new_n544), .C1(new_n202), .C2(new_n203), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT85), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n539), .A2(new_n546), .A3(new_n540), .ZN(new_n547));
  NAND2_X1  g361(.A1(KEYINPUT18), .A2(G131), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n547), .B(new_n548), .ZN(new_n549));
  AOI22_X1  g363(.A1(new_n537), .A2(new_n542), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(G113), .B(G122), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(new_n346), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n533), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n552), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n545), .A2(new_n549), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n542), .A2(new_n536), .A3(new_n196), .ZN(new_n557));
  OAI211_X1 g371(.A(KEYINPUT86), .B(new_n554), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n541), .A2(KEYINPUT17), .A3(G131), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n218), .B(new_n559), .C1(KEYINPUT17), .C2(new_n542), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n560), .A2(new_n555), .A3(new_n552), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n553), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(G475), .A2(G902), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n563), .B(KEYINPUT87), .Z(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT20), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n561), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n552), .B1(new_n560), .B2(new_n555), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n230), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(G475), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n562), .A2(KEYINPUT20), .A3(new_n564), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n567), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n531), .A2(new_n532), .A3(new_n573), .ZN(new_n574));
  AND4_X1   g388(.A1(new_n241), .A2(new_n345), .A3(new_n465), .A4(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(new_n359), .ZN(G3));
  NAND2_X1  g390(.A1(new_n446), .A2(new_n461), .ZN(new_n577));
  INV_X1    g391(.A(new_n447), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT97), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n446), .A2(new_n447), .A3(new_n461), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n411), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n463), .B2(KEYINPUT97), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n567), .A2(new_n571), .A3(new_n572), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT33), .ZN(new_n588));
  NOR3_X1   g402(.A1(new_n519), .A2(new_n520), .A3(new_n474), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n473), .B1(new_n527), .B2(new_n528), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n521), .A2(KEYINPUT33), .A3(new_n529), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n466), .A2(G902), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n230), .B1(new_n589), .B2(new_n590), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n466), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n587), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n586), .A2(new_n597), .A3(new_n419), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n230), .B1(new_n313), .B2(new_n317), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(G472), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(KEYINPUT96), .A3(new_n318), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT96), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n599), .A2(new_n602), .A3(G472), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n409), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n605), .B1(new_n398), .B2(new_n404), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n604), .A2(new_n241), .A3(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n598), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT34), .B(G104), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G6));
  NAND2_X1  g424(.A1(new_n595), .A2(new_n471), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n530), .A2(new_n230), .A3(new_n472), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n586), .A2(new_n613), .A3(new_n587), .A4(new_n419), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n614), .A2(new_n607), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT35), .B(G107), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G9));
  NOR2_X1   g431(.A1(new_n227), .A2(KEYINPUT36), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n222), .B(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n239), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n237), .A2(new_n620), .ZN(new_n621));
  AND4_X1   g435(.A1(new_n574), .A2(new_n465), .A3(new_n604), .A4(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT37), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G110), .ZN(G12));
  NOR2_X1   g438(.A1(new_n585), .A2(new_n410), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n418), .A2(G900), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n626), .B(KEYINPUT98), .Z(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n416), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT99), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n587), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n631), .B1(new_n611), .B2(new_n612), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n625), .A2(new_n345), .A3(new_n621), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(G128), .ZN(G30));
  INV_X1    g448(.A(new_n621), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n303), .B1(new_n307), .B2(new_n333), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n320), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n242), .B1(new_n637), .B2(new_n230), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(KEYINPUT100), .B1(new_n325), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT100), .ZN(new_n641));
  AOI211_X1 g455(.A(new_n641), .B(new_n638), .C1(new_n319), .C2(new_n324), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n635), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n629), .B(KEYINPUT39), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n606), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n646), .A2(KEYINPUT40), .ZN(new_n647));
  OR2_X1    g461(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n587), .B1(new_n611), .B2(new_n612), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n649), .B(new_n411), .C1(new_n646), .C2(KEYINPUT40), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n579), .A2(new_n581), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT38), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(new_n653));
  OR3_X1    g467(.A1(new_n648), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT101), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G143), .ZN(G45));
  AOI211_X1 g470(.A(new_n587), .B(new_n629), .C1(new_n594), .C2(new_n596), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n657), .A2(new_n625), .A3(new_n345), .A4(new_n621), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT102), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G146), .ZN(G48));
  AND3_X1   g474(.A1(new_n382), .A2(new_n384), .A3(new_n393), .ZN(new_n661));
  OAI21_X1  g475(.A(G469), .B1(new_n661), .B2(G902), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n662), .A2(new_n398), .A3(new_n409), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n345), .A2(new_n241), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n598), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT41), .B(G113), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G15));
  NOR2_X1   g482(.A1(new_n614), .A2(new_n665), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(new_n425), .ZN(G18));
  INV_X1    g484(.A(new_n419), .ZN(new_n671));
  NOR3_X1   g485(.A1(new_n613), .A2(new_n573), .A3(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n585), .A2(new_n663), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n672), .A2(new_n673), .A3(new_n345), .A4(new_n621), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G119), .ZN(G21));
  NAND2_X1  g489(.A1(new_n613), .A2(new_n573), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n582), .A2(new_n419), .A3(new_n584), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n676), .A2(new_n677), .A3(new_n663), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n305), .B1(new_n304), .B2(new_n338), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n242), .B(new_n230), .C1(new_n679), .C2(new_n317), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n241), .A2(new_n600), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT103), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G122), .ZN(G24));
  AND3_X1   g498(.A1(new_n600), .A2(new_n621), .A3(new_n680), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n657), .A2(new_n673), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G125), .ZN(G27));
  NAND2_X1  g501(.A1(new_n345), .A2(new_n241), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT104), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n594), .A2(new_n596), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n690), .A2(KEYINPUT42), .A3(new_n573), .A4(new_n630), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n579), .A2(new_n411), .A3(new_n581), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n606), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n345), .A2(new_n696), .A3(new_n241), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n689), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT42), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n410), .A2(new_n692), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n345), .A2(new_n700), .A3(new_n241), .ZN(new_n701));
  INV_X1    g515(.A(new_n657), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n699), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n698), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT105), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G131), .ZN(G33));
  INV_X1    g520(.A(new_n701), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n632), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G134), .ZN(G36));
  INV_X1    g523(.A(KEYINPUT45), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n402), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n400), .A2(KEYINPUT45), .A3(new_n401), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(G469), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(G469), .A2(G902), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n713), .A2(KEYINPUT46), .A3(new_n714), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(new_n398), .A3(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n409), .A3(new_n645), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n587), .A2(KEYINPUT106), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n573), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n690), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(KEYINPUT43), .B1(new_n594), .B2(new_n596), .ZN(new_n726));
  AOI22_X1  g540(.A1(new_n725), .A2(KEYINPUT43), .B1(new_n726), .B2(new_n587), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n727), .A2(new_n603), .A3(new_n601), .A4(new_n621), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n720), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n730), .B(new_n693), .C1(new_n729), .C2(new_n728), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G137), .ZN(G39));
  NAND2_X1  g546(.A1(new_n719), .A2(new_n409), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT47), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n719), .A2(KEYINPUT47), .A3(new_n409), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n692), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OR2_X1    g551(.A1(new_n342), .A2(new_n344), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n702), .A2(new_n241), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n737), .A2(new_n325), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT107), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G140), .ZN(G42));
  INV_X1    g556(.A(KEYINPUT117), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n597), .A2(new_n600), .A3(new_n630), .A4(new_n680), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n745), .B1(new_n531), .B2(new_n532), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n611), .A2(KEYINPUT111), .A3(new_n612), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n345), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n744), .B1(new_n749), .B2(new_n631), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(new_n621), .A3(new_n700), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n704), .A2(new_n708), .A3(new_n751), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n674), .B1(new_n614), .B2(new_n665), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT103), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n681), .B(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n586), .A2(new_n649), .A3(new_n419), .A4(new_n664), .ZN(new_n756));
  OAI22_X1  g570(.A1(new_n755), .A2(new_n756), .B1(new_n665), .B2(new_n598), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT109), .B1(new_n753), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n665), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n690), .A2(new_n573), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n677), .ZN(new_n761));
  AOI22_X1  g575(.A1(new_n759), .A2(new_n761), .B1(new_n678), .B2(new_n682), .ZN(new_n762));
  INV_X1    g576(.A(new_n669), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n762), .A2(new_n763), .A3(new_n764), .A4(new_n674), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n752), .B1(new_n758), .B2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n767), .B1(new_n760), .B2(new_n464), .ZN(new_n768));
  INV_X1    g582(.A(new_n464), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n746), .A2(new_n769), .A3(new_n747), .A4(new_n587), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n597), .A2(KEYINPUT110), .A3(new_n769), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n768), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n607), .ZN(new_n773));
  AOI211_X1 g587(.A(new_n622), .B(new_n575), .C1(new_n772), .C2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n658), .A2(new_n633), .A3(new_n686), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n586), .A2(new_n606), .A3(new_n630), .A4(new_n649), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n643), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT52), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n633), .A2(new_n686), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n606), .A2(new_n630), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n676), .A2(new_n585), .A3(new_n780), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n781), .B(new_n635), .C1(new_n640), .C2(new_n642), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n779), .A2(new_n782), .A3(new_n783), .A4(new_n658), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n774), .A2(new_n778), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT53), .B1(new_n766), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n774), .A2(new_n778), .A3(new_n784), .ZN(new_n787));
  AOI22_X1  g601(.A1(new_n698), .A2(new_n703), .B1(new_n632), .B2(new_n707), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n753), .A2(new_n757), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n789), .A3(KEYINPUT53), .A4(new_n751), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n786), .A2(KEYINPUT54), .A3(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n765), .A2(new_n758), .ZN(new_n795));
  AND3_X1   g609(.A1(new_n704), .A2(new_n708), .A3(new_n751), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n794), .B1(new_n797), .B2(new_n787), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n766), .A2(KEYINPUT53), .A3(new_n785), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n793), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(KEYINPUT112), .B1(new_n792), .B2(new_n800), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n797), .A2(new_n794), .A3(new_n787), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT54), .B1(new_n802), .B2(new_n786), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n804));
  INV_X1    g618(.A(new_n791), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n798), .A2(new_n805), .A3(new_n793), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n801), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n697), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n696), .B1(new_n345), .B2(new_n241), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n663), .A2(new_n692), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n813));
  INV_X1    g627(.A(new_n416), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n813), .B1(new_n727), .B2(new_n814), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n594), .A2(new_n596), .B1(new_n721), .B2(new_n723), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT43), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI211_X1 g632(.A(KEYINPUT43), .B(new_n573), .C1(new_n594), .C2(new_n596), .ZN(new_n819));
  NOR4_X1   g633(.A1(new_n818), .A2(new_n819), .A3(KEYINPUT113), .A4(new_n416), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n811), .B(new_n812), .C1(new_n815), .C2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n690), .A2(new_n817), .A3(new_n587), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n824), .B(new_n814), .C1(new_n817), .C2(new_n816), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT113), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n725), .A2(KEYINPUT43), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n827), .A2(new_n813), .A3(new_n814), .A4(new_n824), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(KEYINPUT115), .A3(new_n811), .A4(new_n812), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n823), .A2(KEYINPUT48), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n640), .A2(new_n642), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n832), .A2(new_n241), .A3(new_n814), .A4(new_n812), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n833), .A2(new_n760), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n831), .A2(new_n413), .A3(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n823), .A2(KEYINPUT48), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n829), .A2(new_n586), .A3(new_n664), .A4(new_n682), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT114), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n755), .B1(new_n826), .B2(new_n828), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(KEYINPUT114), .A3(new_n586), .A4(new_n664), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n835), .A2(KEYINPUT116), .A3(new_n837), .A4(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n843), .A2(new_n831), .A3(new_n413), .A4(new_n834), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n845), .B1(new_n846), .B2(new_n836), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n653), .A2(new_n583), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n841), .A2(new_n664), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT50), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n841), .A2(KEYINPUT50), .A3(new_n664), .A4(new_n849), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n662), .A2(new_n398), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n735), .B(new_n736), .C1(new_n409), .C2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n841), .A2(new_n693), .A3(new_n856), .ZN(new_n857));
  OR3_X1    g671(.A1(new_n833), .A2(new_n573), .A3(new_n690), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n829), .A2(new_n685), .A3(new_n812), .ZN(new_n859));
  AND3_X1   g673(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n854), .A2(new_n860), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n861), .A2(KEYINPUT51), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(KEYINPUT51), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n848), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n743), .B1(new_n808), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n412), .A2(new_n223), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n844), .A2(new_n847), .B1(new_n862), .B2(new_n863), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n868), .A2(KEYINPUT117), .A3(new_n807), .A4(new_n801), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n816), .B1(KEYINPUT49), .B2(new_n855), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(KEYINPUT49), .B2(new_n855), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n241), .A2(new_n409), .A3(new_n411), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT108), .Z(new_n874));
  NAND4_X1  g688(.A1(new_n872), .A2(new_n653), .A3(new_n832), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n870), .A2(new_n875), .ZN(G75));
  NOR2_X1   g690(.A1(new_n786), .A2(new_n791), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(new_n230), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(G210), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT56), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n439), .B(new_n445), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n881), .B(KEYINPUT55), .Z(new_n882));
  AND3_X1   g696(.A1(new_n879), .A2(new_n880), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n882), .B1(new_n879), .B2(new_n880), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n223), .A2(G952), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(G51));
  OAI21_X1  g700(.A(KEYINPUT54), .B1(new_n786), .B2(new_n791), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n887), .A2(new_n806), .A3(KEYINPUT118), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n798), .A2(new_n805), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(new_n890), .A3(KEYINPUT54), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n714), .B(KEYINPUT57), .Z(new_n892));
  NAND3_X1  g706(.A1(new_n888), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n661), .B(KEYINPUT119), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OR3_X1    g709(.A1(new_n877), .A2(new_n230), .A3(new_n713), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n885), .B1(new_n895), .B2(new_n896), .ZN(G54));
  NAND3_X1  g711(.A1(new_n878), .A2(KEYINPUT58), .A3(G475), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(new_n562), .ZN(new_n899));
  INV_X1    g713(.A(new_n885), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(G60));
  AND2_X1   g715(.A1(new_n591), .A2(new_n592), .ZN(new_n902));
  NAND2_X1  g716(.A1(G478), .A2(G902), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT59), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n888), .A2(new_n902), .A3(new_n891), .A4(new_n904), .ZN(new_n905));
  AND3_X1   g719(.A1(new_n905), .A2(KEYINPUT120), .A3(new_n900), .ZN(new_n906));
  AOI21_X1  g720(.A(KEYINPUT120), .B1(new_n905), .B2(new_n900), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n902), .B1(new_n808), .B2(new_n904), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(G63));
  NAND2_X1  g723(.A1(G217), .A2(G902), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT60), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n619), .B(KEYINPUT121), .Z(new_n913));
  NAND3_X1  g727(.A1(new_n889), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n900), .ZN(new_n915));
  OAI21_X1  g729(.A(KEYINPUT61), .B1(new_n915), .B2(KEYINPUT122), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n877), .A2(new_n911), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n900), .B(new_n914), .C1(new_n917), .C2(new_n238), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n916), .B(new_n918), .ZN(G66));
  NAND2_X1  g733(.A1(new_n795), .A2(new_n774), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n223), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n223), .B1(new_n417), .B2(G224), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n921), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n439), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(G898), .B2(new_n223), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n926), .B(new_n928), .ZN(G69));
  NAND3_X1  g743(.A1(new_n654), .A2(new_n658), .A3(new_n779), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT62), .Z(new_n931));
  AND2_X1   g745(.A1(new_n741), .A2(new_n731), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n760), .B1(new_n748), .B2(new_n573), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n707), .A2(new_n645), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n223), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n315), .B(new_n535), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT124), .Z(new_n938));
  NAND2_X1  g752(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(G900), .A2(G953), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n809), .A2(new_n810), .A3(new_n720), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n676), .A2(new_n585), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n775), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n932), .A2(new_n788), .A3(new_n943), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n937), .B(new_n940), .C1(new_n944), .C2(G953), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n939), .A2(KEYINPUT125), .A3(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n223), .B1(G227), .B2(G900), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n947), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n939), .A2(KEYINPUT125), .A3(new_n949), .A4(new_n945), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(G72));
  NAND2_X1  g765(.A1(G472), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT63), .Z(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n935), .B2(new_n920), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n316), .B(KEYINPUT126), .Z(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n954), .A2(new_n304), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n953), .B1(new_n944), .B2(new_n920), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n958), .A2(new_n303), .A3(new_n955), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n326), .A2(new_n320), .A3(new_n331), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n798), .B2(new_n799), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n953), .ZN(new_n962));
  AND4_X1   g776(.A1(new_n900), .A2(new_n957), .A3(new_n959), .A4(new_n962), .ZN(G57));
endmodule


