

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768;

  INV_X1 U375 ( .A(n620), .ZN(n698) );
  XNOR2_X1 U376 ( .A(n752), .B(n576), .ZN(n725) );
  INV_X1 U377 ( .A(G953), .ZN(n755) );
  XNOR2_X1 U378 ( .A(n515), .B(n473), .ZN(n688) );
  XNOR2_X2 U379 ( .A(n518), .B(n517), .ZN(n548) );
  XNOR2_X2 U380 ( .A(n496), .B(n495), .ZN(n518) );
  NOR2_X2 U381 ( .A1(n724), .A2(G953), .ZN(n383) );
  XNOR2_X2 U382 ( .A(n528), .B(G472), .ZN(n620) );
  NOR2_X1 U383 ( .A1(n688), .A2(n689), .ZN(n693) );
  NAND2_X1 U384 ( .A1(n381), .A2(n462), .ZN(n746) );
  AND2_X1 U385 ( .A1(n478), .A2(n476), .ZN(n754) );
  INV_X1 U386 ( .A(n692), .ZN(n581) );
  XNOR2_X1 U387 ( .A(G146), .B(KEYINPUT4), .ZN(n388) );
  INV_X1 U388 ( .A(KEYINPUT32), .ZN(n352) );
  NAND2_X1 U389 ( .A1(n746), .A2(n456), .ZN(n385) );
  AND2_X1 U390 ( .A1(n462), .A2(n659), .ZN(n458) );
  NOR2_X1 U391 ( .A1(n376), .A2(n664), .ZN(n375) );
  NOR2_X1 U392 ( .A1(n688), .A2(n578), .ZN(n664) );
  XNOR2_X1 U393 ( .A(n470), .B(KEYINPUT35), .ZN(n766) );
  OR2_X1 U394 ( .A1(n767), .A2(n763), .ZN(n438) );
  AND2_X1 U395 ( .A1(n414), .A2(n413), .ZN(n412) );
  NOR2_X1 U396 ( .A1(n707), .A2(n689), .ZN(n566) );
  XNOR2_X1 U397 ( .A(n472), .B(n548), .ZN(n752) );
  XNOR2_X2 U398 ( .A(n524), .B(n529), .ZN(n433) );
  XNOR2_X1 U399 ( .A(n388), .B(KEYINPUT69), .ZN(n520) );
  XNOR2_X1 U400 ( .A(n353), .B(n352), .ZN(n768) );
  NOR2_X1 U401 ( .A1(n580), .A2(n365), .ZN(n353) );
  BUF_X1 U402 ( .A(n671), .Z(n354) );
  BUF_X1 U403 ( .A(n372), .Z(n355) );
  XNOR2_X2 U404 ( .A(n433), .B(n431), .ZN(n739) );
  XNOR2_X2 U405 ( .A(n483), .B(G119), .ZN(n524) );
  XNOR2_X2 U406 ( .A(G116), .B(KEYINPUT3), .ZN(n483) );
  NAND2_X1 U407 ( .A1(n725), .A2(G469), .ZN(n393) );
  AND2_X1 U408 ( .A1(n766), .A2(KEYINPUT44), .ZN(n376) );
  NAND2_X1 U409 ( .A1(n398), .A2(n396), .ZN(n401) );
  NAND2_X1 U410 ( .A1(n397), .A2(KEYINPUT1), .ZN(n396) );
  INV_X1 U411 ( .A(n407), .ZN(n397) );
  XNOR2_X1 U412 ( .A(n505), .B(n504), .ZN(n753) );
  XOR2_X1 U413 ( .A(G128), .B(KEYINPUT64), .Z(n496) );
  AND2_X1 U414 ( .A1(n393), .A2(n407), .ZN(n389) );
  XOR2_X1 U415 ( .A(G146), .B(n753), .Z(n535) );
  INV_X1 U416 ( .A(G134), .ZN(n517) );
  XNOR2_X1 U417 ( .A(n435), .B(n586), .ZN(n722) );
  NOR2_X1 U418 ( .A1(n585), .A2(n594), .ZN(n435) );
  NOR2_X1 U419 ( .A1(n596), .A2(n709), .ZN(n597) );
  NAND2_X1 U420 ( .A1(n358), .A2(n648), .ZN(n441) );
  NAND2_X1 U421 ( .A1(G902), .A2(G469), .ZN(n407) );
  XOR2_X1 U422 ( .A(G107), .B(G122), .Z(n540) );
  NOR2_X1 U423 ( .A1(n467), .A2(KEYINPUT45), .ZN(n463) );
  NAND2_X1 U424 ( .A1(n391), .A2(n390), .ZN(n692) );
  NOR2_X1 U425 ( .A1(n401), .A2(n402), .ZN(n391) );
  NAND2_X1 U426 ( .A1(n392), .A2(n404), .ZN(n390) );
  NOR2_X1 U427 ( .A1(n764), .A2(n477), .ZN(n476) );
  XNOR2_X1 U428 ( .A(n479), .B(KEYINPUT48), .ZN(n478) );
  INV_X1 U429 ( .A(n686), .ZN(n477) );
  XNOR2_X1 U430 ( .A(n507), .B(n509), .ZN(n445) );
  XNOR2_X1 U431 ( .A(n506), .B(n508), .ZN(n444) );
  XOR2_X1 U432 ( .A(KEYINPUT9), .B(KEYINPUT98), .Z(n542) );
  XNOR2_X1 U433 ( .A(KEYINPUT7), .B(KEYINPUT97), .ZN(n541) );
  XNOR2_X1 U434 ( .A(n540), .B(n424), .ZN(n544) );
  XNOR2_X1 U435 ( .A(G116), .B(KEYINPUT99), .ZN(n424) );
  XNOR2_X1 U436 ( .A(n533), .B(n360), .ZN(n534) );
  INV_X1 U437 ( .A(n660), .ZN(n417) );
  XNOR2_X1 U438 ( .A(n520), .B(n387), .ZN(n472) );
  XNOR2_X1 U439 ( .A(n519), .B(G137), .ZN(n387) );
  INV_X1 U440 ( .A(G131), .ZN(n519) );
  XOR2_X1 U441 ( .A(G140), .B(KEYINPUT76), .Z(n571) );
  XNOR2_X1 U442 ( .A(n447), .B(KEYINPUT104), .ZN(n651) );
  XNOR2_X1 U443 ( .A(n581), .B(KEYINPUT89), .ZN(n641) );
  XNOR2_X1 U444 ( .A(n637), .B(n421), .ZN(n638) );
  INV_X1 U445 ( .A(KEYINPUT107), .ZN(n421) );
  NAND2_X1 U446 ( .A1(n565), .A2(n415), .ZN(n413) );
  XNOR2_X1 U447 ( .A(G478), .B(n549), .ZN(n589) );
  XNOR2_X1 U448 ( .A(n620), .B(KEYINPUT6), .ZN(n613) );
  XNOR2_X1 U449 ( .A(n514), .B(n516), .ZN(n473) );
  AND2_X1 U450 ( .A1(n418), .A2(n382), .ZN(n420) );
  AND2_X1 U451 ( .A1(n720), .A2(n359), .ZN(n382) );
  NAND2_X1 U452 ( .A1(n400), .A2(n406), .ZN(n405) );
  NOR2_X1 U453 ( .A1(n403), .A2(n400), .ZN(n399) );
  NOR2_X1 U454 ( .A1(G953), .A2(G237), .ZN(n532) );
  NAND2_X1 U455 ( .A1(n597), .A2(KEYINPUT86), .ZN(n468) );
  INV_X1 U456 ( .A(n655), .ZN(n705) );
  NAND2_X1 U457 ( .A1(G237), .A2(G234), .ZN(n557) );
  NAND2_X1 U458 ( .A1(n395), .A2(KEYINPUT1), .ZN(n394) );
  INV_X1 U459 ( .A(n405), .ZN(n395) );
  AND2_X1 U460 ( .A1(n393), .A2(n367), .ZN(n392) );
  XOR2_X1 U461 ( .A(KEYINPUT93), .B(KEYINPUT20), .Z(n513) );
  AND2_X1 U462 ( .A1(n439), .A2(n437), .ZN(n479) );
  XNOR2_X1 U463 ( .A(n438), .B(n657), .ZN(n437) );
  XNOR2_X1 U464 ( .A(G122), .B(G143), .ZN(n530) );
  XOR2_X1 U465 ( .A(KEYINPUT11), .B(G131), .Z(n531) );
  XNOR2_X1 U466 ( .A(G902), .B(KEYINPUT15), .ZN(n660) );
  XOR2_X1 U467 ( .A(KEYINPUT18), .B(KEYINPUT77), .Z(n489) );
  XNOR2_X1 U468 ( .A(KEYINPUT17), .B(KEYINPUT90), .ZN(n488) );
  OR2_X1 U469 ( .A1(G902), .A2(G237), .ZN(n553) );
  INV_X1 U470 ( .A(KEYINPUT0), .ZN(n415) );
  NOR2_X1 U471 ( .A1(n565), .A2(n415), .ZN(n410) );
  NAND2_X1 U472 ( .A1(n692), .A2(n693), .ZN(n594) );
  XNOR2_X1 U473 ( .A(n540), .B(n432), .ZN(n431) );
  INV_X1 U474 ( .A(KEYINPUT16), .ZN(n432) );
  AND2_X1 U475 ( .A1(n754), .A2(KEYINPUT2), .ZN(n456) );
  OR2_X1 U476 ( .A1(n754), .A2(KEYINPUT2), .ZN(n459) );
  XNOR2_X1 U477 ( .A(n475), .B(n474), .ZN(n658) );
  INV_X1 U478 ( .A(KEYINPUT39), .ZN(n474) );
  XNOR2_X1 U479 ( .A(n446), .B(KEYINPUT80), .ZN(n644) );
  XNOR2_X1 U480 ( .A(n539), .B(n538), .ZN(n590) );
  NAND2_X1 U481 ( .A1(n622), .A2(n693), .ZN(n591) );
  XNOR2_X1 U482 ( .A(n442), .B(n535), .ZN(n737) );
  XNOR2_X1 U483 ( .A(n443), .B(n511), .ZN(n442) );
  XNOR2_X1 U484 ( .A(n445), .B(n444), .ZN(n443) );
  XNOR2_X1 U485 ( .A(n547), .B(n422), .ZN(n734) );
  XNOR2_X1 U486 ( .A(n548), .B(n546), .ZN(n422) );
  XNOR2_X1 U487 ( .A(G107), .B(G104), .ZN(n574) );
  XNOR2_X1 U488 ( .A(n573), .B(n572), .ZN(n575) );
  XNOR2_X1 U489 ( .A(n656), .B(KEYINPUT40), .ZN(n767) );
  AND2_X1 U490 ( .A1(n658), .A2(n678), .ZN(n656) );
  XNOR2_X1 U491 ( .A(n640), .B(n423), .ZN(n642) );
  XNOR2_X1 U492 ( .A(KEYINPUT88), .B(KEYINPUT36), .ZN(n423) );
  NOR2_X1 U493 ( .A1(n722), .A2(n592), .ZN(n587) );
  OR2_X1 U494 ( .A1(n613), .A2(n580), .ZN(n568) );
  XNOR2_X1 U495 ( .A(n750), .B(n426), .ZN(G69) );
  XNOR2_X1 U496 ( .A(n751), .B(KEYINPUT125), .ZN(n426) );
  INV_X1 U497 ( .A(KEYINPUT60), .ZN(n427) );
  INV_X1 U498 ( .A(KEYINPUT118), .ZN(n419) );
  XOR2_X1 U499 ( .A(n622), .B(KEYINPUT103), .Z(n356) );
  NOR2_X1 U500 ( .A1(n698), .A2(n579), .ZN(n357) );
  AND2_X1 U501 ( .A1(n643), .A2(n683), .ZN(n358) );
  XNOR2_X1 U502 ( .A(KEYINPUT117), .B(n723), .ZN(n359) );
  AND2_X1 U503 ( .A1(n532), .A2(G214), .ZN(n360) );
  AND2_X1 U504 ( .A1(n553), .A2(G210), .ZN(n361) );
  XNOR2_X1 U505 ( .A(KEYINPUT79), .B(n613), .ZN(n362) );
  AND2_X1 U506 ( .A1(n375), .A2(n460), .ZN(n363) );
  XNOR2_X1 U507 ( .A(KEYINPUT28), .B(n621), .ZN(n364) );
  NAND2_X1 U508 ( .A1(n362), .A2(n582), .ZN(n365) );
  INV_X1 U509 ( .A(KEYINPUT1), .ZN(n403) );
  AND2_X1 U510 ( .A1(n532), .A2(G210), .ZN(n366) );
  AND2_X1 U511 ( .A1(n407), .A2(n403), .ZN(n367) );
  INV_X1 U512 ( .A(G902), .ZN(n406) );
  XOR2_X1 U513 ( .A(n663), .B(n662), .Z(n368) );
  XOR2_X1 U514 ( .A(n503), .B(n502), .Z(n369) );
  XNOR2_X1 U515 ( .A(KEYINPUT59), .B(KEYINPUT66), .ZN(n370) );
  XOR2_X1 U516 ( .A(KEYINPUT56), .B(KEYINPUT120), .Z(n371) );
  NAND2_X1 U517 ( .A1(n411), .A2(n410), .ZN(n409) );
  NOR2_X1 U518 ( .A1(n647), .A2(n709), .ZN(n440) );
  NAND2_X1 U519 ( .A1(n554), .A2(n704), .ZN(n372) );
  NAND2_X1 U520 ( .A1(n554), .A2(n704), .ZN(n639) );
  AND2_X2 U521 ( .A1(n416), .A2(n429), .ZN(n373) );
  AND2_X2 U522 ( .A1(n416), .A2(n429), .ZN(n736) );
  NOR2_X1 U523 ( .A1(n654), .A2(n655), .ZN(n475) );
  XNOR2_X1 U524 ( .A(n372), .B(n555), .ZN(n374) );
  XNOR2_X1 U525 ( .A(n639), .B(n555), .ZN(n623) );
  NAND2_X1 U526 ( .A1(n373), .A2(G210), .ZN(n455) );
  NAND2_X1 U527 ( .A1(n736), .A2(G217), .ZN(n436) );
  NAND2_X1 U528 ( .A1(n736), .A2(G472), .ZN(n450) );
  NAND2_X1 U529 ( .A1(n449), .A2(n461), .ZN(n448) );
  XNOR2_X1 U530 ( .A(n450), .B(n368), .ZN(n449) );
  NAND2_X1 U531 ( .A1(n481), .A2(n461), .ZN(n480) );
  XNOR2_X1 U532 ( .A(n436), .B(n482), .ZN(n481) );
  OR2_X1 U533 ( .A1(n725), .A2(n405), .ZN(n404) );
  OR2_X1 U534 ( .A1(n651), .A2(n374), .ZN(n446) );
  INV_X1 U535 ( .A(n738), .ZN(n461) );
  NAND2_X1 U536 ( .A1(n378), .A2(n377), .ZN(n469) );
  NAND2_X1 U537 ( .A1(n380), .A2(n363), .ZN(n377) );
  NAND2_X1 U538 ( .A1(n379), .A2(KEYINPUT86), .ZN(n378) );
  NAND2_X1 U539 ( .A1(n380), .A2(n375), .ZN(n379) );
  XNOR2_X2 U540 ( .A(n484), .B(n584), .ZN(n380) );
  NAND2_X1 U541 ( .A1(n381), .A2(n458), .ZN(n457) );
  AND2_X2 U542 ( .A1(n465), .A2(n466), .ZN(n381) );
  NAND2_X2 U543 ( .A1(n412), .A2(n409), .ZN(n384) );
  NAND2_X1 U544 ( .A1(n384), .A2(n566), .ZN(n567) );
  XNOR2_X2 U545 ( .A(n567), .B(KEYINPUT22), .ZN(n580) );
  XNOR2_X1 U546 ( .A(n383), .B(KEYINPUT53), .ZN(G75) );
  XNOR2_X1 U547 ( .A(n384), .B(n434), .ZN(n592) );
  NAND2_X1 U548 ( .A1(n700), .A2(n384), .ZN(n595) );
  AND2_X2 U549 ( .A1(n385), .A2(n417), .ZN(n416) );
  NAND2_X1 U550 ( .A1(n429), .A2(n385), .ZN(n418) );
  XNOR2_X2 U551 ( .A(n386), .B(n361), .ZN(n554) );
  NAND2_X1 U552 ( .A1(n552), .A2(n660), .ZN(n386) );
  NAND2_X1 U553 ( .A1(n404), .A2(n389), .ZN(n622) );
  NOR2_X1 U554 ( .A1(n725), .A2(n394), .ZN(n402) );
  NAND2_X1 U555 ( .A1(n725), .A2(n399), .ZN(n398) );
  INV_X1 U556 ( .A(G469), .ZN(n400) );
  XNOR2_X1 U557 ( .A(n408), .B(n491), .ZN(n569) );
  XNOR2_X2 U558 ( .A(G101), .B(KEYINPUT67), .ZN(n408) );
  XNOR2_X1 U559 ( .A(n408), .B(KEYINPUT5), .ZN(n526) );
  INV_X1 U560 ( .A(n374), .ZN(n411) );
  NAND2_X1 U561 ( .A1(n623), .A2(n415), .ZN(n414) );
  XNOR2_X1 U562 ( .A(n420), .B(n419), .ZN(n724) );
  NAND2_X1 U563 ( .A1(n612), .A2(n613), .ZN(n637) );
  XNOR2_X1 U564 ( .A(n425), .B(n523), .ZN(n525) );
  XNOR2_X1 U565 ( .A(n524), .B(n366), .ZN(n425) );
  NAND2_X1 U566 ( .A1(n485), .A2(n461), .ZN(n428) );
  XNOR2_X1 U567 ( .A(n428), .B(n427), .ZN(G60) );
  INV_X1 U568 ( .A(n469), .ZN(n464) );
  AND2_X2 U569 ( .A1(n457), .A2(n459), .ZN(n429) );
  XNOR2_X1 U570 ( .A(n430), .B(n583), .ZN(n599) );
  NAND2_X1 U571 ( .A1(n671), .A2(n768), .ZN(n430) );
  NAND2_X1 U572 ( .A1(n464), .A2(n463), .ZN(n462) );
  XNOR2_X1 U573 ( .A(n452), .B(KEYINPUT100), .ZN(n451) );
  INV_X1 U574 ( .A(KEYINPUT92), .ZN(n434) );
  NAND2_X1 U575 ( .A1(n602), .A2(n468), .ZN(n467) );
  NOR2_X1 U576 ( .A1(n441), .A2(n440), .ZN(n439) );
  NAND2_X1 U577 ( .A1(n364), .A2(n356), .ZN(n447) );
  XNOR2_X1 U578 ( .A(n448), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U579 ( .A1(n451), .A2(n357), .ZN(n671) );
  NOR2_X2 U580 ( .A1(n580), .A2(n692), .ZN(n452) );
  XNOR2_X1 U581 ( .A(n453), .B(n371), .ZN(G51) );
  NAND2_X1 U582 ( .A1(n454), .A2(n461), .ZN(n453) );
  XNOR2_X1 U583 ( .A(n455), .B(n369), .ZN(n454) );
  NOR2_X1 U584 ( .A1(n597), .A2(KEYINPUT86), .ZN(n460) );
  NAND2_X1 U585 ( .A1(n469), .A2(KEYINPUT45), .ZN(n465) );
  NAND2_X1 U586 ( .A1(n467), .A2(KEYINPUT45), .ZN(n466) );
  NAND2_X1 U587 ( .A1(n471), .A2(n626), .ZN(n470) );
  XNOR2_X1 U588 ( .A(n587), .B(KEYINPUT34), .ZN(n471) );
  NAND2_X1 U589 ( .A1(n631), .A2(n632), .ZN(n654) );
  XNOR2_X1 U590 ( .A(n480), .B(KEYINPUT123), .ZN(G66) );
  INV_X1 U591 ( .A(n737), .ZN(n482) );
  INV_X1 U592 ( .A(n554), .ZN(n616) );
  XNOR2_X1 U593 ( .A(n499), .B(n500), .ZN(n552) );
  NAND2_X1 U594 ( .A1(n599), .A2(KEYINPUT44), .ZN(n484) );
  XNOR2_X1 U595 ( .A(n487), .B(n486), .ZN(n485) );
  XNOR2_X1 U596 ( .A(n732), .B(n370), .ZN(n486) );
  NAND2_X1 U597 ( .A1(n736), .A2(G475), .ZN(n487) );
  BUF_X1 U598 ( .A(n552), .Z(n501) );
  INV_X1 U599 ( .A(KEYINPUT87), .ZN(n583) );
  INV_X1 U600 ( .A(n569), .ZN(n573) );
  INV_X1 U601 ( .A(n613), .ZN(n585) );
  INV_X1 U602 ( .A(KEYINPUT19), .ZN(n555) );
  INV_X1 U603 ( .A(G143), .ZN(n495) );
  XNOR2_X1 U604 ( .A(n575), .B(n574), .ZN(n576) );
  INV_X1 U605 ( .A(n661), .ZN(n663) );
  XNOR2_X1 U606 ( .A(KEYINPUT13), .B(G475), .ZN(n538) );
  NOR2_X1 U607 ( .A1(G952), .A2(n755), .ZN(n738) );
  XOR2_X1 U608 ( .A(KEYINPUT119), .B(KEYINPUT54), .Z(n503) );
  XOR2_X1 U609 ( .A(G104), .B(G113), .Z(n529) );
  XNOR2_X1 U610 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U611 ( .A(n739), .B(n490), .ZN(n500) );
  XNOR2_X1 U612 ( .A(G110), .B(KEYINPUT71), .ZN(n491) );
  XNOR2_X1 U613 ( .A(n569), .B(KEYINPUT78), .ZN(n494) );
  AND2_X1 U614 ( .A1(G224), .A2(n755), .ZN(n492) );
  XNOR2_X1 U615 ( .A(n520), .B(n492), .ZN(n493) );
  XNOR2_X1 U616 ( .A(n494), .B(n493), .ZN(n498) );
  XNOR2_X1 U617 ( .A(G125), .B(n518), .ZN(n497) );
  XNOR2_X1 U618 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U619 ( .A(n501), .B(KEYINPUT55), .ZN(n502) );
  XOR2_X1 U620 ( .A(G125), .B(KEYINPUT70), .Z(n505) );
  XNOR2_X1 U621 ( .A(G140), .B(KEYINPUT10), .ZN(n504) );
  XOR2_X1 U622 ( .A(G110), .B(G137), .Z(n507) );
  XNOR2_X1 U623 ( .A(G119), .B(G128), .ZN(n506) );
  XOR2_X1 U624 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n509) );
  XNOR2_X1 U625 ( .A(KEYINPUT75), .B(KEYINPUT83), .ZN(n508) );
  NAND2_X1 U626 ( .A1(G234), .A2(n755), .ZN(n510) );
  XOR2_X1 U627 ( .A(KEYINPUT8), .B(n510), .Z(n545) );
  NAND2_X1 U628 ( .A1(G221), .A2(n545), .ZN(n511) );
  NOR2_X1 U629 ( .A1(n737), .A2(G902), .ZN(n515) );
  NAND2_X1 U630 ( .A1(G234), .A2(n660), .ZN(n512) );
  XNOR2_X1 U631 ( .A(n513), .B(n512), .ZN(n550) );
  NAND2_X1 U632 ( .A1(n550), .A2(G217), .ZN(n514) );
  XOR2_X1 U633 ( .A(KEYINPUT25), .B(KEYINPUT74), .Z(n516) );
  XOR2_X1 U634 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n522) );
  XNOR2_X1 U635 ( .A(G113), .B(KEYINPUT73), .ZN(n521) );
  XNOR2_X1 U636 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U637 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U638 ( .A(n752), .B(n527), .ZN(n661) );
  NOR2_X1 U639 ( .A1(n661), .A2(G902), .ZN(n528) );
  XNOR2_X1 U640 ( .A(n529), .B(KEYINPUT12), .ZN(n537) );
  XNOR2_X1 U641 ( .A(n531), .B(n530), .ZN(n533) );
  XNOR2_X1 U642 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U643 ( .A(n537), .B(n536), .ZN(n732) );
  NOR2_X1 U644 ( .A1(G902), .A2(n732), .ZN(n539) );
  INV_X1 U645 ( .A(n590), .ZN(n588) );
  XNOR2_X1 U646 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U647 ( .A(n544), .B(n543), .Z(n547) );
  NAND2_X1 U648 ( .A1(G217), .A2(n545), .ZN(n546) );
  NOR2_X1 U649 ( .A1(G902), .A2(n734), .ZN(n549) );
  NAND2_X1 U650 ( .A1(n588), .A2(n589), .ZN(n707) );
  NAND2_X1 U651 ( .A1(n550), .A2(G221), .ZN(n551) );
  XNOR2_X1 U652 ( .A(n551), .B(KEYINPUT21), .ZN(n689) );
  NAND2_X1 U653 ( .A1(G214), .A2(n553), .ZN(n704) );
  NAND2_X1 U654 ( .A1(n755), .A2(G952), .ZN(n603) );
  NAND2_X1 U655 ( .A1(G953), .A2(G902), .ZN(n604) );
  OR2_X1 U656 ( .A1(n604), .A2(G898), .ZN(n556) );
  NAND2_X1 U657 ( .A1(n603), .A2(n556), .ZN(n558) );
  XOR2_X1 U658 ( .A(KEYINPUT14), .B(n557), .Z(n608) );
  INV_X1 U659 ( .A(n608), .ZN(n717) );
  NAND2_X1 U660 ( .A1(n558), .A2(n717), .ZN(n560) );
  INV_X1 U661 ( .A(KEYINPUT91), .ZN(n559) );
  NAND2_X1 U662 ( .A1(n560), .A2(n559), .ZN(n564) );
  NOR2_X1 U663 ( .A1(G898), .A2(n755), .ZN(n742) );
  NAND2_X1 U664 ( .A1(n742), .A2(KEYINPUT91), .ZN(n561) );
  NOR2_X1 U665 ( .A1(n406), .A2(n561), .ZN(n562) );
  NAND2_X1 U666 ( .A1(n562), .A2(n717), .ZN(n563) );
  NAND2_X1 U667 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U668 ( .A(KEYINPUT85), .B(n568), .ZN(n577) );
  NAND2_X1 U669 ( .A1(G227), .A2(n755), .ZN(n570) );
  XNOR2_X1 U670 ( .A(n571), .B(n570), .ZN(n572) );
  NAND2_X1 U671 ( .A1(n577), .A2(n581), .ZN(n578) );
  INV_X1 U672 ( .A(n688), .ZN(n579) );
  AND2_X1 U673 ( .A1(n641), .A2(n688), .ZN(n582) );
  INV_X1 U674 ( .A(KEYINPUT65), .ZN(n584) );
  XNOR2_X1 U675 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n586) );
  NOR2_X1 U676 ( .A1(n588), .A2(n589), .ZN(n626) );
  NAND2_X1 U677 ( .A1(n590), .A2(n589), .ZN(n611) );
  INV_X1 U678 ( .A(n611), .ZN(n678) );
  NOR2_X1 U679 ( .A1(n590), .A2(n589), .ZN(n680) );
  NOR2_X1 U680 ( .A1(n678), .A2(n680), .ZN(n709) );
  XNOR2_X1 U681 ( .A(KEYINPUT94), .B(n591), .ZN(n630) );
  OR2_X1 U682 ( .A1(n592), .A2(n630), .ZN(n593) );
  NOR2_X1 U683 ( .A1(n698), .A2(n593), .ZN(n666) );
  NOR2_X1 U684 ( .A1(n620), .A2(n594), .ZN(n700) );
  XNOR2_X1 U685 ( .A(n595), .B(KEYINPUT31), .ZN(n681) );
  NOR2_X1 U686 ( .A1(n666), .A2(n681), .ZN(n596) );
  NOR2_X1 U687 ( .A1(n766), .A2(KEYINPUT44), .ZN(n598) );
  XNOR2_X1 U688 ( .A(KEYINPUT68), .B(n598), .ZN(n601) );
  INV_X1 U689 ( .A(n599), .ZN(n600) );
  NAND2_X1 U690 ( .A1(n601), .A2(n600), .ZN(n602) );
  INV_X1 U691 ( .A(n603), .ZN(n606) );
  NOR2_X1 U692 ( .A1(G900), .A2(n604), .ZN(n605) );
  NOR2_X1 U693 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U694 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U695 ( .A(n609), .B(KEYINPUT81), .ZN(n627) );
  NOR2_X1 U696 ( .A1(n689), .A2(n627), .ZN(n610) );
  NAND2_X1 U697 ( .A1(n610), .A2(n688), .ZN(n619) );
  NOR2_X1 U698 ( .A1(n611), .A2(n619), .ZN(n612) );
  NOR2_X1 U699 ( .A1(n692), .A2(n637), .ZN(n614) );
  NAND2_X1 U700 ( .A1(n614), .A2(n704), .ZN(n615) );
  XNOR2_X1 U701 ( .A(n615), .B(KEYINPUT43), .ZN(n617) );
  NAND2_X1 U702 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U703 ( .A(KEYINPUT101), .B(n618), .ZN(n764) );
  NOR2_X1 U704 ( .A1(n620), .A2(n619), .ZN(n621) );
  INV_X1 U705 ( .A(n644), .ZN(n676) );
  NAND2_X1 U706 ( .A1(KEYINPUT82), .A2(n709), .ZN(n624) );
  NAND2_X1 U707 ( .A1(n676), .A2(n624), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n625), .A2(KEYINPUT47), .ZN(n648) );
  INV_X1 U709 ( .A(n626), .ZN(n635) );
  INV_X1 U710 ( .A(n627), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n698), .A2(n704), .ZN(n628) );
  XNOR2_X1 U712 ( .A(KEYINPUT30), .B(n628), .ZN(n629) );
  NOR2_X1 U713 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U714 ( .A1(n616), .A2(n654), .ZN(n633) );
  XOR2_X1 U715 ( .A(KEYINPUT102), .B(n633), .Z(n634) );
  NOR2_X1 U716 ( .A1(n635), .A2(n634), .ZN(n674) );
  NOR2_X1 U717 ( .A1(KEYINPUT82), .A2(KEYINPUT47), .ZN(n636) );
  NOR2_X1 U718 ( .A1(n674), .A2(n636), .ZN(n643) );
  NOR2_X1 U719 ( .A1(n355), .A2(n638), .ZN(n640) );
  NAND2_X1 U720 ( .A1(n642), .A2(n641), .ZN(n683) );
  NOR2_X1 U721 ( .A1(n644), .A2(KEYINPUT47), .ZN(n646) );
  INV_X1 U722 ( .A(KEYINPUT82), .ZN(n645) );
  NOR2_X1 U723 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U724 ( .A(KEYINPUT46), .B(KEYINPUT84), .Z(n657) );
  XOR2_X1 U725 ( .A(KEYINPUT38), .B(n616), .Z(n655) );
  NAND2_X1 U726 ( .A1(n705), .A2(n704), .ZN(n708) );
  NOR2_X1 U727 ( .A1(n707), .A2(n708), .ZN(n650) );
  XOR2_X1 U728 ( .A(KEYINPUT41), .B(KEYINPUT105), .Z(n649) );
  XNOR2_X1 U729 ( .A(n650), .B(n649), .ZN(n721) );
  NOR2_X1 U730 ( .A1(n651), .A2(n721), .ZN(n653) );
  XNOR2_X1 U731 ( .A(KEYINPUT106), .B(KEYINPUT42), .ZN(n652) );
  XNOR2_X1 U732 ( .A(n653), .B(n652), .ZN(n763) );
  NAND2_X1 U733 ( .A1(n658), .A2(n680), .ZN(n686) );
  INV_X1 U734 ( .A(KEYINPUT2), .ZN(n659) );
  XOR2_X1 U735 ( .A(KEYINPUT62), .B(KEYINPUT108), .Z(n662) );
  XOR2_X1 U736 ( .A(G101), .B(n664), .Z(G3) );
  NAND2_X1 U737 ( .A1(n666), .A2(n678), .ZN(n665) );
  XNOR2_X1 U738 ( .A(n665), .B(G104), .ZN(G6) );
  XOR2_X1 U739 ( .A(KEYINPUT26), .B(KEYINPUT109), .Z(n668) );
  NAND2_X1 U740 ( .A1(n666), .A2(n680), .ZN(n667) );
  XNOR2_X1 U741 ( .A(n668), .B(n667), .ZN(n670) );
  XOR2_X1 U742 ( .A(G107), .B(KEYINPUT27), .Z(n669) );
  XNOR2_X1 U743 ( .A(n670), .B(n669), .ZN(G9) );
  XNOR2_X1 U744 ( .A(n354), .B(G110), .ZN(G12) );
  XOR2_X1 U745 ( .A(G128), .B(KEYINPUT29), .Z(n673) );
  NAND2_X1 U746 ( .A1(n680), .A2(n676), .ZN(n672) );
  XNOR2_X1 U747 ( .A(n673), .B(n672), .ZN(G30) );
  XOR2_X1 U748 ( .A(G143), .B(n674), .Z(n675) );
  XNOR2_X1 U749 ( .A(KEYINPUT110), .B(n675), .ZN(G45) );
  NAND2_X1 U750 ( .A1(n676), .A2(n678), .ZN(n677) );
  XNOR2_X1 U751 ( .A(n677), .B(G146), .ZN(G48) );
  NAND2_X1 U752 ( .A1(n681), .A2(n678), .ZN(n679) );
  XNOR2_X1 U753 ( .A(n679), .B(G113), .ZN(G15) );
  NAND2_X1 U754 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U755 ( .A(n682), .B(G116), .ZN(G18) );
  XNOR2_X1 U756 ( .A(KEYINPUT111), .B(KEYINPUT37), .ZN(n684) );
  XNOR2_X1 U757 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U758 ( .A(G125), .B(n685), .ZN(G27) );
  XNOR2_X1 U759 ( .A(G134), .B(KEYINPUT112), .ZN(n687) );
  XNOR2_X1 U760 ( .A(n687), .B(n686), .ZN(G36) );
  XOR2_X1 U761 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n691) );
  NAND2_X1 U762 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U763 ( .A(n691), .B(n690), .ZN(n696) );
  NOR2_X1 U764 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U765 ( .A(KEYINPUT50), .B(n694), .Z(n695) );
  NAND2_X1 U766 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U767 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U768 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U769 ( .A(n701), .B(KEYINPUT115), .ZN(n702) );
  XNOR2_X1 U770 ( .A(KEYINPUT51), .B(n702), .ZN(n703) );
  NOR2_X1 U771 ( .A1(n721), .A2(n703), .ZN(n715) );
  NOR2_X1 U772 ( .A1(n705), .A2(n704), .ZN(n706) );
  NOR2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n712) );
  NOR2_X1 U774 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U775 ( .A(n710), .B(KEYINPUT116), .ZN(n711) );
  NOR2_X1 U776 ( .A1(n712), .A2(n711), .ZN(n713) );
  NOR2_X1 U777 ( .A1(n722), .A2(n713), .ZN(n714) );
  NOR2_X1 U778 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U779 ( .A(KEYINPUT52), .B(n716), .Z(n719) );
  AND2_X1 U780 ( .A1(G952), .A2(n717), .ZN(n718) );
  NAND2_X1 U781 ( .A1(n719), .A2(n718), .ZN(n720) );
  NOR2_X1 U782 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U783 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n727) );
  XNOR2_X1 U784 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n726) );
  XNOR2_X1 U785 ( .A(n727), .B(n726), .ZN(n728) );
  XOR2_X1 U786 ( .A(n725), .B(n728), .Z(n730) );
  NAND2_X1 U787 ( .A1(n373), .A2(G469), .ZN(n729) );
  XNOR2_X1 U788 ( .A(n730), .B(n729), .ZN(n731) );
  NOR2_X1 U789 ( .A1(n738), .A2(n731), .ZN(G54) );
  NAND2_X1 U790 ( .A1(G478), .A2(n373), .ZN(n733) );
  XNOR2_X1 U791 ( .A(n734), .B(n733), .ZN(n735) );
  NOR2_X1 U792 ( .A1(n738), .A2(n735), .ZN(G63) );
  XOR2_X1 U793 ( .A(n739), .B(G110), .Z(n740) );
  XNOR2_X1 U794 ( .A(G101), .B(n740), .ZN(n741) );
  NOR2_X1 U795 ( .A1(n742), .A2(n741), .ZN(n751) );
  INV_X1 U796 ( .A(G898), .ZN(n745) );
  NAND2_X1 U797 ( .A1(G953), .A2(G224), .ZN(n743) );
  XOR2_X1 U798 ( .A(KEYINPUT61), .B(n743), .Z(n744) );
  NOR2_X1 U799 ( .A1(n745), .A2(n744), .ZN(n749) );
  NAND2_X1 U800 ( .A1(n746), .A2(n755), .ZN(n747) );
  XOR2_X1 U801 ( .A(KEYINPUT124), .B(n747), .Z(n748) );
  NOR2_X1 U802 ( .A1(n749), .A2(n748), .ZN(n750) );
  XOR2_X1 U803 ( .A(n753), .B(n752), .Z(n757) );
  XOR2_X1 U804 ( .A(n757), .B(n754), .Z(n756) );
  NAND2_X1 U805 ( .A1(n756), .A2(n755), .ZN(n762) );
  XNOR2_X1 U806 ( .A(G227), .B(n757), .ZN(n758) );
  NAND2_X1 U807 ( .A1(n758), .A2(G900), .ZN(n759) );
  XNOR2_X1 U808 ( .A(KEYINPUT126), .B(n759), .ZN(n760) );
  NAND2_X1 U809 ( .A1(n760), .A2(G953), .ZN(n761) );
  NAND2_X1 U810 ( .A1(n762), .A2(n761), .ZN(G72) );
  XOR2_X1 U811 ( .A(G137), .B(n763), .Z(G39) );
  XNOR2_X1 U812 ( .A(G140), .B(n764), .ZN(n765) );
  XNOR2_X1 U813 ( .A(n765), .B(KEYINPUT113), .ZN(G42) );
  XOR2_X1 U814 ( .A(G122), .B(n766), .Z(G24) );
  XOR2_X1 U815 ( .A(n767), .B(G131), .Z(G33) );
  XNOR2_X1 U816 ( .A(n768), .B(G119), .ZN(G21) );
endmodule

