//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1282, new_n1283;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  NOR2_X1   g0006(.A1(G97), .A2(G107), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(G50), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n211), .B1(new_n212), .B2(new_n213), .C1(new_n203), .C2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G232), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n202), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n210), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  OR2_X1    g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n204), .A2(new_n205), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n223), .A2(new_n212), .ZN(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n210), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT0), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n222), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n217), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n235), .B(new_n236), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n237), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n245), .B(new_n248), .Z(G351));
  NAND2_X1  g0049(.A1(G33), .A2(G41), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G1), .A3(G13), .ZN(new_n251));
  INV_X1    g0051(.A(G41), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT5), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n254), .B(G45), .C1(new_n252), .C2(KEYINPUT5), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT78), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n253), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G45), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G1), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT5), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(G41), .ZN(new_n261));
  AOI21_X1  g0061(.A(KEYINPUT78), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  OAI211_X1 g0062(.A(G270), .B(new_n251), .C1(new_n257), .C2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  OAI211_X1 g0065(.A(G264), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n219), .A2(G1698), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(new_n264), .B2(new_n265), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n271), .A2(G303), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n266), .A2(new_n268), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n255), .A2(new_n256), .ZN(new_n277));
  INV_X1    g0077(.A(G274), .ZN(new_n278));
  INV_X1    g0078(.A(new_n225), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n278), .B1(new_n279), .B2(new_n250), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n259), .A2(KEYINPUT78), .A3(new_n261), .ZN(new_n281));
  NAND4_X1  g0081(.A1(new_n277), .A2(new_n280), .A3(new_n281), .A4(new_n253), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n263), .A2(new_n276), .A3(G179), .A4(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g0084(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n225), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n254), .A2(G13), .A3(G20), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n254), .A2(G33), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n287), .A2(G116), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G116), .ZN(new_n291));
  AOI22_X1  g0091(.A1(new_n285), .A2(new_n225), .B1(G20), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(G33), .A2(G283), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n293), .B(new_n226), .C1(G33), .C2(new_n218), .ZN(new_n294));
  AND3_X1   g0094(.A1(new_n292), .A2(KEYINPUT20), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(KEYINPUT20), .B1(new_n292), .B2(new_n294), .ZN(new_n296));
  OAI221_X1 g0096(.A(new_n290), .B1(G116), .B2(new_n288), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n284), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n263), .A2(new_n276), .A3(new_n282), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n297), .B1(G200), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G190), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(new_n299), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n297), .A2(new_n299), .A3(G169), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT80), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n303), .A2(new_n304), .A3(KEYINPUT21), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT21), .B1(new_n303), .B2(new_n304), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n298), .B(new_n302), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n271), .A2(new_n272), .ZN(new_n309));
  INV_X1    g0109(.A(G1698), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n309), .A2(G222), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G77), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n309), .A2(G1698), .ZN(new_n313));
  INV_X1    g0113(.A(G223), .ZN(new_n314));
  OAI221_X1 g0114(.A(new_n311), .B1(new_n312), .B2(new_n309), .C1(new_n313), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n275), .ZN(new_n316));
  XNOR2_X1  g0116(.A(KEYINPUT66), .B(G45), .ZN(new_n317));
  OAI211_X1 g0117(.A(new_n254), .B(G274), .C1(new_n317), .C2(G41), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n251), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n319), .B1(G226), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n316), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(new_n301), .ZN(new_n324));
  OR2_X1    g0124(.A1(new_n324), .A2(KEYINPUT70), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(KEYINPUT70), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n325), .A2(new_n326), .B1(G200), .B2(new_n323), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n226), .B1(new_n223), .B2(new_n212), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n328), .B(KEYINPUT68), .ZN(new_n329));
  NOR2_X1   g0129(.A1(KEYINPUT8), .A2(G58), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT67), .B(G58), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n330), .B1(new_n332), .B2(KEYINPUT8), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n226), .A2(G33), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NOR2_X1   g0135(.A1(G20), .A2(G33), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n333), .A2(new_n335), .B1(G150), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n287), .B1(new_n329), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n288), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n212), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n286), .B1(new_n254), .B2(G20), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n340), .B1(new_n342), .B2(new_n212), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT9), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n344), .B(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n327), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n347), .B(KEYINPUT10), .ZN(new_n348));
  INV_X1    g0148(.A(G169), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n323), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(G179), .B2(new_n323), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(new_n344), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n333), .A2(new_n342), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(new_n339), .B2(new_n333), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n204), .B(new_n205), .C1(new_n331), .C2(new_n203), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n358), .A2(G20), .B1(G159), .B2(new_n336), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n264), .A2(new_n265), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT7), .B1(new_n360), .B2(new_n226), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n271), .A2(KEYINPUT7), .A3(new_n226), .A4(new_n272), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(G68), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n359), .A2(KEYINPUT16), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n286), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n271), .A2(new_n226), .A3(new_n272), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT7), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT73), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n369), .A2(new_n370), .A3(new_n362), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n363), .A2(KEYINPUT73), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(G68), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n359), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT16), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT74), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n366), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT16), .B1(new_n373), .B2(new_n359), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT74), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n357), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n321), .A2(G232), .ZN(new_n382));
  NOR2_X1   g0182(.A1(G223), .A2(G1698), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n383), .B1(new_n213), .B2(G1698), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n384), .A2(new_n309), .B1(G33), .B2(G87), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n382), .B(new_n318), .C1(new_n385), .C2(new_n251), .ZN(new_n386));
  INV_X1    g0186(.A(G179), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(G169), .B2(new_n386), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT18), .B1(new_n381), .B2(new_n389), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n286), .B(new_n365), .C1(new_n379), .C2(KEYINPUT74), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n376), .A2(new_n377), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n356), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT18), .ZN(new_n394));
  INV_X1    g0194(.A(new_n389), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n386), .A2(G190), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT75), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT75), .ZN(new_n399));
  INV_X1    g0199(.A(G200), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n399), .B1(new_n386), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n398), .B1(new_n401), .B2(new_n397), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n356), .B(new_n402), .C1(new_n391), .C2(new_n392), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT17), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n378), .A2(new_n380), .ZN(new_n406));
  NAND4_X1  g0206(.A1(new_n406), .A2(KEYINPUT17), .A3(new_n356), .A4(new_n402), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n390), .A2(new_n396), .A3(new_n405), .A4(new_n407), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n309), .A2(G232), .A3(G1698), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G97), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n309), .A2(new_n310), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n409), .B(new_n410), .C1(new_n411), .C2(new_n213), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n275), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT13), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n321), .A2(G238), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n415), .A2(new_n318), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n413), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n414), .B1(new_n413), .B2(new_n416), .ZN(new_n418));
  OAI21_X1  g0218(.A(G169), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT14), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n413), .A2(new_n416), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT13), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n413), .A2(new_n414), .A3(new_n416), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n425), .A2(KEYINPUT14), .A3(G169), .ZN(new_n426));
  XNOR2_X1  g0226(.A(new_n424), .B(KEYINPUT71), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n418), .A2(new_n387), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n421), .A2(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n341), .A2(G68), .ZN(new_n430));
  XOR2_X1   g0230(.A(new_n430), .B(KEYINPUT72), .Z(new_n431));
  INV_X1    g0231(.A(new_n336), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n432), .A2(new_n212), .ZN(new_n433));
  OAI22_X1  g0233(.A1(new_n334), .A2(new_n312), .B1(new_n226), .B2(G68), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n286), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT11), .ZN(new_n436));
  AND2_X1   g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n288), .A2(G68), .ZN(new_n438));
  XNOR2_X1  g0238(.A(new_n438), .B(KEYINPUT12), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n435), .A2(new_n436), .ZN(new_n440));
  NOR4_X1   g0240(.A1(new_n431), .A2(new_n437), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n429), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n427), .A2(G190), .A3(new_n423), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n425), .A2(G200), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n442), .A2(new_n446), .ZN(new_n447));
  XOR2_X1   g0247(.A(KEYINPUT8), .B(G58), .Z(new_n448));
  AOI22_X1  g0248(.A1(new_n448), .A2(new_n336), .B1(G20), .B2(G77), .ZN(new_n449));
  XNOR2_X1  g0249(.A(KEYINPUT15), .B(G87), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(KEYINPUT69), .A3(new_n335), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT69), .B1(new_n451), .B2(new_n335), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n286), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n288), .A2(G77), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n456), .B1(new_n341), .B2(G77), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n360), .A2(G107), .ZN(new_n459));
  OAI221_X1 g0259(.A(new_n459), .B1(new_n313), .B2(new_n214), .C1(new_n217), .C2(new_n411), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n275), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n319), .B1(G244), .B2(new_n321), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n458), .B1(new_n464), .B2(G190), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n463), .A2(G200), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n458), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n468), .B1(new_n349), .B2(new_n463), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n464), .A2(new_n387), .ZN(new_n470));
  AND2_X1   g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n447), .A2(new_n467), .A3(new_n472), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n354), .A2(new_n408), .A3(new_n473), .ZN(new_n474));
  AND2_X1   g0274(.A1(KEYINPUT4), .A2(G244), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n310), .B(new_n475), .C1(new_n264), .C2(new_n265), .ZN(new_n476));
  INV_X1    g0276(.A(G244), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n477), .B1(new_n271), .B2(new_n272), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n476), .B(new_n293), .C1(new_n478), .C2(KEYINPUT4), .ZN(new_n479));
  OAI21_X1  g0279(.A(G250), .B1(new_n264), .B2(new_n265), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n310), .B1(new_n480), .B2(KEYINPUT4), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n275), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  OAI211_X1 g0282(.A(G257), .B(new_n251), .C1(new_n257), .C2(new_n262), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n282), .A3(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G179), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n483), .A2(new_n282), .ZN(new_n486));
  AOI21_X1  g0286(.A(G169), .B1(new_n486), .B2(new_n482), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n287), .A2(KEYINPUT77), .A3(new_n288), .A4(new_n289), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT77), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n288), .A2(new_n289), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n490), .B1(new_n491), .B2(new_n286), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n489), .A2(new_n492), .A3(G97), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n339), .A2(new_n218), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n371), .A2(G107), .A3(new_n372), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n432), .A2(new_n312), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT6), .ZN(new_n499));
  AND2_X1   g0299(.A1(G97), .A2(G107), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(new_n207), .ZN(new_n501));
  INV_X1    g0301(.A(G107), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n502), .A2(KEYINPUT6), .A3(G97), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g0304(.A(KEYINPUT76), .B(new_n498), .C1(new_n504), .C2(new_n226), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT76), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n226), .B1(new_n501), .B2(new_n503), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n506), .B1(new_n507), .B2(new_n497), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n496), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n495), .B1(new_n509), .B2(new_n286), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n488), .A2(new_n511), .ZN(new_n512));
  AND3_X1   g0312(.A1(new_n482), .A2(new_n282), .A3(new_n483), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n513), .A2(G200), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n484), .A2(G190), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n510), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n288), .A2(G107), .ZN(new_n518));
  XNOR2_X1  g0318(.A(new_n518), .B(KEYINPUT25), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n489), .A2(new_n492), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n519), .B1(new_n520), .B2(new_n502), .ZN(new_n521));
  AOI21_X1  g0321(.A(G20), .B1(new_n271), .B2(new_n272), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT22), .ZN(new_n523));
  OAI21_X1  g0323(.A(KEYINPUT82), .B1(new_n523), .B2(KEYINPUT81), .ZN(new_n524));
  OR3_X1    g0324(.A1(new_n523), .A2(KEYINPUT81), .A3(KEYINPUT82), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n522), .A2(G87), .A3(new_n524), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G33), .A2(G116), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n527), .A2(G20), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT23), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n226), .B2(G107), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n502), .A2(KEYINPUT23), .A3(G20), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n526), .A2(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n522), .A2(G87), .B1(new_n525), .B2(new_n524), .ZN(new_n534));
  OAI21_X1  g0334(.A(KEYINPUT24), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n534), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT24), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n536), .A2(new_n537), .A3(new_n526), .A4(new_n532), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n521), .B1(new_n539), .B2(new_n286), .ZN(new_n540));
  OAI211_X1 g0340(.A(G257), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n541));
  OAI211_X1 g0341(.A(G250), .B(new_n310), .C1(new_n264), .C2(new_n265), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G294), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n275), .ZN(new_n545));
  OAI211_X1 g0345(.A(G264), .B(new_n251), .C1(new_n257), .C2(new_n262), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n546), .A3(new_n282), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n400), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(G190), .B2(new_n547), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n540), .A2(new_n549), .ZN(new_n550));
  OR2_X1    g0350(.A1(new_n547), .A2(G179), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n547), .A2(new_n349), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n287), .B1(new_n535), .B2(new_n538), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n551), .B(new_n552), .C1(new_n553), .C2(new_n521), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n550), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT19), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n226), .B1(new_n410), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(G87), .B2(new_n208), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n556), .B1(new_n334), .B2(new_n218), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n226), .B(G68), .C1(new_n264), .C2(new_n265), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n561), .A2(new_n286), .B1(new_n339), .B2(new_n450), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n520), .B2(new_n450), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n254), .A2(G45), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(G250), .ZN(new_n565));
  OAI21_X1  g0365(.A(KEYINPUT79), .B1(new_n275), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT79), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n251), .A2(new_n567), .A3(G250), .A4(new_n564), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n566), .A2(new_n568), .B1(new_n259), .B2(new_n280), .ZN(new_n569));
  OAI211_X1 g0369(.A(G244), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n570));
  OAI211_X1 g0370(.A(G238), .B(new_n310), .C1(new_n264), .C2(new_n265), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n570), .A2(new_n571), .A3(new_n527), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n275), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n349), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n563), .B(new_n575), .C1(G179), .C2(new_n574), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n574), .A2(G200), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n489), .A2(new_n492), .A3(G87), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n569), .A2(new_n573), .A3(G190), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n577), .A2(new_n578), .A3(new_n562), .A4(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n555), .A2(new_n581), .ZN(new_n582));
  AND4_X1   g0382(.A1(new_n308), .A2(new_n474), .A3(new_n517), .A4(new_n582), .ZN(G372));
  NOR2_X1   g0383(.A1(new_n446), .A2(new_n472), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n405), .B(new_n407), .C1(new_n584), .C2(new_n442), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n390), .A2(new_n396), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n352), .B1(new_n587), .B2(new_n348), .ZN(new_n588));
  INV_X1    g0388(.A(new_n474), .ZN(new_n589));
  INV_X1    g0389(.A(new_n576), .ZN(new_n590));
  AND3_X1   g0390(.A1(new_n562), .A2(KEYINPUT83), .A3(new_n578), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT83), .B1(new_n562), .B2(new_n578), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n577), .B(new_n579), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  AND4_X1   g0393(.A1(new_n512), .A2(new_n516), .A3(new_n550), .A4(new_n593), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n554), .B(new_n298), .C1(new_n305), .C2(new_n306), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n590), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n488), .A2(new_n511), .A3(new_n580), .A4(new_n576), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT26), .ZN(new_n598));
  OAI21_X1  g0398(.A(KEYINPUT84), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n581), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT84), .ZN(new_n601));
  NOR3_X1   g0401(.A1(new_n510), .A2(new_n485), .A3(new_n487), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n600), .A2(new_n601), .A3(new_n602), .A4(KEYINPUT26), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n593), .A2(new_n488), .A3(new_n511), .A4(new_n576), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n598), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n599), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n596), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n588), .B1(new_n589), .B2(new_n608), .ZN(G369));
  NOR2_X1   g0409(.A1(new_n305), .A2(new_n306), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n297), .B2(new_n284), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n254), .A2(new_n226), .A3(G13), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n612), .A2(KEYINPUT27), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(KEYINPUT27), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(G213), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(G343), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n555), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n617), .B(KEYINPUT85), .ZN(new_n621));
  INV_X1    g0421(.A(new_n621), .ZN(new_n622));
  OR2_X1    g0422(.A1(new_n554), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT86), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n620), .A2(KEYINPUT86), .A3(new_n623), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n297), .A2(new_n617), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n308), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n611), .B2(new_n629), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(G330), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n617), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n619), .B1(new_n540), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n554), .B2(new_n634), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n628), .A2(new_n637), .ZN(G399));
  INV_X1    g0438(.A(new_n229), .ZN(new_n639));
  OR3_X1    g0439(.A1(new_n639), .A2(KEYINPUT87), .A3(G41), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT87), .B1(new_n639), .B2(G41), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(G1), .A3(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n224), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n644), .B(KEYINPUT88), .C1(new_n645), .C2(new_n642), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(KEYINPUT88), .B2(new_n644), .ZN(new_n647));
  XOR2_X1   g0447(.A(new_n647), .B(KEYINPUT28), .Z(new_n648));
  AOI21_X1  g0448(.A(new_n622), .B1(new_n596), .B2(new_n606), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(KEYINPUT29), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT90), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n651), .B1(new_n604), .B2(new_n598), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n593), .A2(new_n576), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n653), .A2(KEYINPUT90), .A3(KEYINPUT26), .A4(new_n602), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n597), .A2(new_n598), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n652), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n617), .B1(new_n656), .B2(new_n596), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n650), .B1(KEYINPUT29), .B2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n582), .A2(new_n517), .A3(new_n308), .A4(new_n621), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n547), .A2(new_n299), .A3(new_n387), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT89), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n574), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n569), .A2(new_n573), .A3(KEYINPUT89), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n660), .A2(new_n484), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n569), .A2(new_n545), .A3(new_n573), .A4(new_n546), .ZN(new_n665));
  NOR4_X1   g0465(.A1(new_n484), .A2(new_n665), .A3(new_n283), .A4(KEYINPUT30), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT30), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n665), .A2(new_n283), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n667), .B1(new_n668), .B2(new_n513), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n664), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(new_n617), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT31), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n670), .A2(KEYINPUT31), .A3(new_n622), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n659), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n658), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n648), .B1(new_n677), .B2(G1), .ZN(G364));
  INV_X1    g0478(.A(new_n642), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n226), .A2(G13), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT91), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n254), .B1(new_n681), .B2(G45), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n349), .A2(KEYINPUT95), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n226), .B1(KEYINPUT95), .B2(new_n349), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n225), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n226), .A2(new_n387), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(G200), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(new_n301), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n691), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n695), .A2(new_n301), .A3(G200), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI221_X1 g0497(.A(new_n309), .B1(new_n694), .B2(new_n212), .C1(new_n331), .C2(new_n697), .ZN(new_n698));
  NOR3_X1   g0498(.A1(new_n695), .A2(G190), .A3(G200), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n699), .A2(KEYINPUT96), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n699), .A2(KEYINPUT96), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n698), .B1(new_n703), .B2(G77), .ZN(new_n704));
  NOR4_X1   g0504(.A1(new_n226), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT97), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(KEYINPUT97), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(G159), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT32), .ZN(new_n711));
  NOR4_X1   g0511(.A1(new_n226), .A2(new_n301), .A3(new_n400), .A4(G179), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(G87), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n387), .A2(new_n400), .A3(G190), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G20), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n715), .B1(G97), .B2(new_n717), .ZN(new_n718));
  NOR4_X1   g0518(.A1(new_n226), .A2(new_n400), .A3(G179), .A4(G190), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n502), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n692), .A2(G190), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(G68), .B2(new_n722), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n704), .A2(new_n711), .A3(new_n718), .A4(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n717), .ZN(new_n725));
  INV_X1    g0525(.A(G294), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n722), .ZN(new_n728));
  XOR2_X1   g0528(.A(KEYINPUT33), .B(G317), .Z(new_n729));
  INV_X1    g0529(.A(G303), .ZN(new_n730));
  OAI22_X1  g0530(.A1(new_n728), .A2(new_n729), .B1(new_n730), .B2(new_n713), .ZN(new_n731));
  AOI211_X1 g0531(.A(new_n727), .B(new_n731), .C1(G326), .C2(new_n693), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n703), .A2(G311), .ZN(new_n733));
  INV_X1    g0533(.A(new_n708), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G329), .ZN(new_n735));
  INV_X1    g0535(.A(G283), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n720), .A2(new_n736), .ZN(new_n737));
  AOI211_X1 g0537(.A(new_n309), .B(new_n737), .C1(G322), .C2(new_n696), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n732), .A2(new_n733), .A3(new_n735), .A4(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n690), .B1(new_n724), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G13), .A2(G33), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n689), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n639), .A2(new_n360), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT92), .ZN(new_n746));
  AOI22_X1  g0546(.A1(new_n746), .A2(G355), .B1(new_n291), .B2(new_n639), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(KEYINPUT93), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n360), .A2(new_n229), .ZN(new_n749));
  XOR2_X1   g0549(.A(new_n749), .B(KEYINPUT94), .Z(new_n750));
  NOR2_X1   g0550(.A1(new_n645), .A2(new_n317), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n751), .B1(G45), .B2(new_n245), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n748), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n747), .A2(KEYINPUT93), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI211_X1 g0555(.A(new_n685), .B(new_n740), .C1(new_n744), .C2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n743), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n756), .B1(new_n631), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n632), .A2(new_n685), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n631), .A2(G330), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(G396));
  NOR2_X1   g0561(.A1(new_n689), .A2(new_n741), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n736), .A2(new_n728), .B1(new_n694), .B2(new_n730), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n764), .B1(new_n703), .B2(G116), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT98), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n713), .A2(new_n502), .B1(new_n720), .B2(new_n714), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n360), .B1(new_n218), .B2(new_n725), .C1(new_n697), .C2(new_n726), .ZN(new_n768));
  AOI211_X1 g0568(.A(new_n767), .B(new_n768), .C1(G311), .C2(new_n734), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n696), .A2(G143), .B1(new_n693), .B2(G137), .ZN(new_n770));
  INV_X1    g0570(.A(G150), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n770), .B1(new_n771), .B2(new_n728), .C1(new_n702), .C2(new_n709), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT34), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n720), .A2(new_n203), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(G50), .B2(new_n712), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n360), .B1(new_n332), .B2(new_n717), .ZN(new_n777));
  INV_X1    g0577(.A(G132), .ZN(new_n778));
  OAI211_X1 g0578(.A(new_n776), .B(new_n777), .C1(new_n708), .C2(new_n778), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(new_n772), .B2(new_n773), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n766), .A2(new_n769), .B1(new_n774), .B2(new_n780), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n684), .B1(G77), .B2(new_n763), .C1(new_n781), .C2(new_n690), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n469), .A2(new_n470), .A3(new_n634), .ZN(new_n783));
  AOI22_X1  g0583(.A1(new_n465), .A2(new_n466), .B1(new_n458), .B2(new_n617), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n783), .B1(new_n784), .B2(new_n471), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n782), .B1(new_n741), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n607), .A2(new_n621), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n785), .ZN(new_n788));
  INV_X1    g0588(.A(new_n785), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n649), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n676), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n684), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n788), .A2(new_n676), .A3(new_n790), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n786), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(G384));
  NOR2_X1   g0596(.A1(new_n681), .A2(new_n254), .ZN(new_n797));
  INV_X1    g0597(.A(G330), .ZN(new_n798));
  OR2_X1    g0598(.A1(new_n441), .A2(new_n634), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n445), .B(new_n799), .C1(new_n429), .C2(new_n441), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n429), .A2(new_n799), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n785), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AND4_X1   g0602(.A1(new_n546), .A2(new_n569), .A3(new_n545), .A4(new_n573), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n513), .A2(new_n803), .A3(new_n284), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(KEYINPUT30), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n668), .A2(new_n667), .A3(new_n513), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n634), .B1(new_n807), .B2(new_n664), .ZN(new_n808));
  OAI21_X1  g0608(.A(KEYINPUT100), .B1(new_n808), .B2(KEYINPUT31), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT100), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n671), .A2(new_n810), .A3(new_n672), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n809), .A2(new_n659), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n670), .A2(KEYINPUT31), .A3(new_n617), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(KEYINPUT101), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT101), .ZN(new_n815));
  NAND4_X1  g0615(.A1(new_n670), .A2(new_n815), .A3(KEYINPUT31), .A4(new_n617), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n802), .B1(new_n812), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(KEYINPUT102), .ZN(new_n819));
  AOI21_X1  g0619(.A(KEYINPUT16), .B1(new_n359), .B2(new_n364), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n366), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n821), .A2(new_n357), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n822), .A2(new_n615), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n408), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n822), .B1(new_n389), .B2(new_n615), .ZN(new_n825));
  INV_X1    g0625(.A(new_n403), .ZN(new_n826));
  OAI21_X1  g0626(.A(KEYINPUT37), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n393), .A2(new_n395), .ZN(new_n828));
  INV_X1    g0628(.A(new_n615), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n393), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT37), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n828), .A2(new_n830), .A3(new_n831), .A4(new_n403), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n827), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n824), .A2(KEYINPUT38), .A3(new_n833), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n403), .B1(new_n381), .B2(new_n389), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n381), .A2(new_n615), .ZN(new_n836));
  OAI21_X1  g0636(.A(KEYINPUT37), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n832), .A2(new_n837), .B1(new_n408), .B2(new_n836), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n834), .B1(new_n838), .B2(KEYINPUT38), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n814), .A2(new_n816), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n840), .A2(new_n659), .A3(new_n811), .A4(new_n809), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT102), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n841), .A2(new_n842), .A3(new_n802), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n819), .A2(KEYINPUT40), .A3(new_n839), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT103), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT40), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n837), .A2(new_n832), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n408), .A2(new_n836), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT38), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n846), .B1(new_n851), .B2(new_n834), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT103), .ZN(new_n853));
  NAND4_X1  g0653(.A1(new_n852), .A2(new_n853), .A3(new_n819), .A4(new_n843), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n824), .A2(new_n833), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n850), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n834), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n857), .A2(new_n802), .A3(new_n841), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n845), .A2(new_n854), .B1(new_n846), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n841), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n589), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n798), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n859), .B2(new_n861), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n586), .A2(new_n829), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n800), .A2(new_n801), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n790), .B2(new_n783), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n864), .B1(new_n867), .B2(new_n857), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT39), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n824), .A2(KEYINPUT38), .A3(new_n833), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT38), .B1(new_n847), .B2(new_n848), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n856), .A2(KEYINPUT39), .A3(new_n834), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n429), .A2(new_n441), .A3(new_n617), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n868), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n658), .A2(new_n474), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n588), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n876), .B(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n797), .B1(new_n863), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n879), .B2(new_n863), .ZN(new_n881));
  INV_X1    g0681(.A(new_n504), .ZN(new_n882));
  OR2_X1    g0682(.A1(new_n882), .A2(KEYINPUT35), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(KEYINPUT35), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n883), .A2(G116), .A3(new_n227), .A4(new_n884), .ZN(new_n885));
  XOR2_X1   g0685(.A(new_n885), .B(KEYINPUT36), .Z(new_n886));
  AOI211_X1 g0686(.A(new_n312), .B(new_n645), .C1(G68), .C2(new_n332), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n888), .A2(KEYINPUT99), .B1(new_n212), .B2(G68), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(KEYINPUT99), .B2(new_n888), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n254), .A2(G13), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n886), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n881), .A2(new_n892), .ZN(G367));
  INV_X1    g0693(.A(new_n750), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n241), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n744), .B1(new_n229), .B2(new_n450), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n684), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n309), .B1(new_n697), .B2(new_n771), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(G77), .B2(new_n719), .ZN(new_n899));
  INV_X1    g0699(.A(G137), .ZN(new_n900));
  OAI221_X1 g0700(.A(new_n899), .B1(new_n900), .B2(new_n708), .C1(new_n212), .C2(new_n702), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n693), .A2(G143), .B1(new_n332), .B2(new_n712), .ZN(new_n902));
  OAI221_X1 g0702(.A(new_n902), .B1(new_n203), .B2(new_n725), .C1(new_n709), .C2(new_n728), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n360), .B1(new_n697), .B2(new_n730), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(G97), .B2(new_n719), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n734), .A2(G317), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n905), .B(new_n906), .C1(new_n736), .C2(new_n702), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n712), .A2(G116), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT46), .ZN(new_n909));
  XOR2_X1   g0709(.A(KEYINPUT107), .B(G311), .Z(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n693), .A2(new_n911), .B1(G107), .B2(new_n717), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n909), .B(new_n912), .C1(new_n726), .C2(new_n728), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n901), .A2(new_n903), .B1(new_n907), .B2(new_n913), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(KEYINPUT47), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n897), .B1(new_n915), .B2(new_n689), .ZN(new_n916));
  OR3_X1    g0716(.A1(new_n591), .A2(new_n592), .A3(new_n634), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n653), .A2(new_n917), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n917), .A2(new_n576), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n916), .B1(new_n757), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n637), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n517), .B1(new_n510), .B2(new_n621), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n512), .B2(new_n621), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT105), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n924), .A2(new_n925), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(new_n628), .ZN(new_n930));
  INV_X1    g0730(.A(KEYINPUT45), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n929), .A2(KEYINPUT45), .A3(new_n628), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT44), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(new_n628), .B2(new_n929), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n928), .A2(new_n626), .A3(KEYINPUT44), .A4(new_n627), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(KEYINPUT106), .B(new_n922), .C1(new_n934), .C2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT106), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n932), .A2(new_n933), .B1(new_n936), .B2(new_n937), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n940), .B1(new_n941), .B2(new_n637), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n620), .B1(new_n636), .B2(new_n618), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n633), .B(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n677), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n941), .B2(new_n637), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n939), .A2(new_n942), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n677), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n642), .B(KEYINPUT41), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n683), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n928), .A2(new_n620), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT42), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n512), .B1(new_n928), .B2(new_n554), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(new_n621), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n920), .ZN(new_n957));
  XOR2_X1   g0757(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n928), .A2(new_n637), .ZN(new_n962));
  INV_X1    g0762(.A(new_n956), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT43), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n959), .B1(new_n964), .B2(new_n957), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n961), .B(new_n962), .C1(new_n963), .C2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n963), .A2(new_n965), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n967), .A2(new_n960), .B1(new_n637), .B2(new_n928), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n921), .B1(new_n951), .B2(new_n969), .ZN(G387));
  NAND2_X1  g0770(.A1(new_n944), .A2(new_n683), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n696), .A2(G317), .B1(new_n693), .B2(G322), .ZN(new_n972));
  OAI221_X1 g0772(.A(new_n972), .B1(new_n728), .B2(new_n910), .C1(new_n702), .C2(new_n730), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT48), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n974), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n712), .A2(G294), .B1(new_n717), .B2(G283), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT49), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n979), .A2(KEYINPUT113), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(KEYINPUT113), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n734), .A2(G326), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n309), .B1(new_n719), .B2(G116), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n980), .A2(new_n981), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n703), .A2(G68), .B1(G150), .B2(new_n734), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n333), .A2(new_n722), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n693), .A2(G159), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT112), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n309), .B1(new_n218), .B2(new_n720), .C1(new_n697), .C2(new_n212), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n713), .A2(new_n312), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n725), .A2(new_n450), .ZN(new_n991));
  NOR3_X1   g0791(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n985), .A2(new_n986), .A3(new_n988), .A4(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n690), .B1(new_n984), .B2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(new_n237), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n995), .A2(new_n317), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(KEYINPUT108), .ZN(new_n997));
  INV_X1    g0797(.A(new_n643), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n258), .B1(new_n203), .B2(new_n312), .C1(new_n998), .C2(KEYINPUT109), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(KEYINPUT109), .B2(new_n998), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT110), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n448), .A2(new_n212), .ZN(new_n1002));
  XOR2_X1   g0802(.A(new_n1002), .B(KEYINPUT50), .Z(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n996), .A2(KEYINPUT108), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n997), .A2(new_n750), .A3(new_n1004), .A4(new_n1005), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n746), .A2(new_n998), .B1(new_n502), .B2(new_n639), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n685), .B1(new_n1008), .B2(new_n744), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT111), .Z(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n636), .B2(new_n757), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n945), .A2(new_n679), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n677), .A2(new_n944), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n971), .B1(new_n994), .B2(new_n1011), .C1(new_n1012), .C2(new_n1013), .ZN(G393));
  XNOR2_X1  g0814(.A(new_n941), .B(new_n922), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n945), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n947), .B(new_n679), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n744), .B1(new_n218), .B2(new_n229), .C1(new_n894), .C2(new_n248), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n309), .B(new_n721), .C1(new_n703), .C2(G294), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n696), .A2(G311), .B1(new_n693), .B2(G317), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT52), .Z(new_n1021));
  OAI22_X1  g0821(.A1(new_n713), .A2(new_n736), .B1(new_n291), .B2(new_n725), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G303), .B2(new_n722), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n734), .A2(G322), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1019), .A2(new_n1021), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(new_n696), .A2(G159), .B1(new_n693), .B2(G150), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT51), .Z(new_n1027));
  OAI22_X1  g0827(.A1(new_n728), .A2(new_n212), .B1(new_n312), .B2(new_n725), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G68), .B2(new_n712), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n703), .A2(new_n448), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n309), .B1(new_n720), .B2(new_n714), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(new_n734), .B2(G143), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1027), .A2(new_n1029), .A3(new_n1030), .A4(new_n1032), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1025), .A2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n684), .B(new_n1018), .C1(new_n1034), .C2(new_n690), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n928), .B2(new_n743), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n1015), .B2(new_n683), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1017), .A2(new_n1037), .ZN(G390));
  NAND2_X1  g0838(.A1(new_n872), .A2(new_n873), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n622), .B(new_n785), .C1(new_n596), .C2(new_n606), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n783), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n865), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n874), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n656), .A2(new_n596), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n784), .A2(new_n471), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1045), .A2(new_n634), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n866), .B1(new_n1048), .B2(new_n783), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n874), .B1(new_n851), .B2(new_n834), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n1039), .A2(new_n1044), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n675), .A2(new_n865), .A3(G330), .A4(new_n789), .ZN(new_n1053));
  AOI21_X1  g0853(.A(KEYINPUT114), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n872), .A2(new_n873), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1043), .B1(new_n870), .B2(new_n871), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1056), .A2(new_n1049), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT114), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1053), .ZN(new_n1059));
  NOR4_X1   g0859(.A1(new_n1055), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n860), .A2(new_n798), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n802), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1039), .A2(new_n1044), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  NOR3_X1   g0865(.A1(new_n1054), .A2(new_n1060), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n474), .A2(new_n1061), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n877), .A2(new_n1067), .A3(new_n588), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n676), .A2(new_n789), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n866), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1062), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n1041), .B2(new_n1040), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n1053), .A2(new_n783), .A3(new_n1048), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n841), .A2(G330), .A3(new_n789), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n866), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1074), .A2(KEYINPUT115), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(KEYINPUT115), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1073), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1066), .A2(new_n1069), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1063), .A2(new_n1064), .A3(new_n1053), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n1058), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1052), .A2(KEYINPUT114), .A3(new_n1053), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n802), .B(new_n1061), .C1(new_n1055), .C2(new_n1057), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1083), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1080), .A2(new_n1069), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n642), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1081), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1066), .A2(new_n683), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n684), .B1(new_n333), .B2(new_n763), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n502), .A2(new_n728), .B1(new_n694), .B2(new_n736), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n775), .B(new_n1092), .C1(G77), .C2(new_n717), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n734), .A2(G294), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n703), .A2(G97), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n309), .B(new_n715), .C1(G116), .C2(new_n696), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .A4(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(KEYINPUT54), .B(G143), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n702), .A2(new_n1098), .B1(new_n900), .B2(new_n728), .ZN(new_n1099));
  OR2_X1    g0899(.A1(new_n1099), .A2(KEYINPUT116), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(KEYINPUT116), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n712), .A2(G150), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1102), .A2(KEYINPUT53), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n734), .A2(G125), .B1(KEYINPUT53), .B2(new_n1102), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1100), .A2(new_n1101), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(G128), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n697), .A2(new_n778), .B1(new_n694), .B2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G159), .B2(new_n717), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n309), .B1(new_n720), .B2(new_n212), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT117), .ZN(new_n1110));
  OR2_X1    g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1108), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1097), .B1(new_n1105), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1091), .B1(new_n1114), .B2(new_n689), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1039), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n742), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1117), .B(KEYINPUT118), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1089), .A2(new_n1090), .A3(new_n1118), .ZN(G378));
  NOR2_X1   g0919(.A1(new_n344), .A2(new_n615), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(new_n1120), .B(KEYINPUT55), .ZN(new_n1121));
  OR2_X1    g0921(.A1(new_n354), .A2(new_n1121), .ZN(new_n1122));
  XOR2_X1   g0922(.A(KEYINPUT121), .B(KEYINPUT56), .Z(new_n1123));
  NAND2_X1  g0923(.A1(new_n354), .A2(new_n1121), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1122), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1123), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n845), .A2(new_n854), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n798), .B1(new_n858), .B2(new_n846), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n1129), .A2(new_n876), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n876), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1128), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n841), .A2(new_n842), .A3(new_n802), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n842), .B1(new_n841), .B2(new_n802), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n853), .B1(new_n1136), .B2(new_n852), .ZN(new_n1137));
  OAI21_X1  g0937(.A(KEYINPUT40), .B1(new_n870), .B2(new_n871), .ZN(new_n1138));
  NOR4_X1   g0938(.A1(new_n1138), .A2(new_n1134), .A3(new_n1135), .A4(KEYINPUT103), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1130), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n876), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1129), .A2(new_n876), .A3(new_n1130), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1142), .A2(new_n1143), .A3(new_n1127), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1133), .A2(new_n1144), .A3(new_n683), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n684), .B1(G50), .B2(new_n763), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n309), .A2(G41), .ZN(new_n1147));
  AOI211_X1 g0947(.A(G50), .B(new_n1147), .C1(new_n270), .C2(new_n252), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n1147), .B1(new_n203), .B2(new_n725), .C1(new_n697), .C2(new_n502), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(G283), .B2(new_n734), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n218), .A2(new_n728), .B1(new_n694), .B2(new_n291), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n720), .A2(new_n331), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1151), .A2(new_n990), .A3(new_n1152), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1150), .B(new_n1153), .C1(new_n450), .C2(new_n702), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT58), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1148), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  AOI211_X1 g0956(.A(G33), .B(G41), .C1(new_n719), .C2(G159), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT120), .B(G124), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n722), .A2(G132), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1159), .B1(new_n713), .B2(new_n1098), .C1(new_n697), .C2(new_n1106), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n693), .A2(G125), .B1(G150), .B2(new_n717), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n1161), .B(KEYINPUT119), .Z(new_n1162));
  AOI211_X1 g0962(.A(new_n1160), .B(new_n1162), .C1(G137), .C2(new_n703), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT59), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1157), .B1(new_n708), .B2(new_n1158), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1163), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1156), .B1(new_n1155), .B2(new_n1154), .C1(new_n1165), .C2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1146), .B1(new_n1168), .B2(new_n689), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n1127), .B2(new_n742), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1145), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NOR3_X1   g0972(.A1(new_n1131), .A2(new_n1132), .A3(new_n1128), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1127), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1080), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1069), .B1(new_n1086), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(KEYINPUT57), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1133), .A2(new_n1144), .A3(KEYINPUT57), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1068), .B1(new_n1066), .B2(new_n1080), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n679), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1172), .B1(new_n1178), .B2(new_n1181), .ZN(G375));
  OAI21_X1  g0982(.A(new_n684), .B1(G68), .B2(new_n763), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n865), .A2(new_n742), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n708), .A2(new_n730), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n697), .A2(new_n736), .B1(new_n450), .B2(new_n725), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1185), .B(new_n1186), .C1(new_n703), .C2(G107), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n693), .A2(G294), .B1(G97), .B2(new_n712), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1187), .B(new_n1188), .C1(new_n291), .C2(new_n728), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n309), .B1(new_n719), .B2(G77), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT122), .Z(new_n1191));
  NOR2_X1   g0991(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  OR2_X1    g0992(.A1(new_n1192), .A2(KEYINPUT123), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(KEYINPUT123), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n703), .A2(G150), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n694), .A2(new_n778), .B1(new_n709), .B2(new_n713), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n728), .A2(new_n1098), .B1(new_n212), .B2(new_n725), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n734), .A2(G128), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n360), .B(new_n1152), .C1(G137), .C2(new_n696), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1195), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1193), .A2(new_n1194), .A3(new_n1201), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1183), .B(new_n1184), .C1(new_n689), .C2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(new_n1080), .B2(new_n683), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1087), .A2(new_n950), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1079), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n1077), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1207), .A2(new_n1068), .A3(new_n1073), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1204), .B1(new_n1205), .B2(new_n1209), .ZN(G381));
  INV_X1    g1010(.A(G390), .ZN(new_n1211));
  INV_X1    g1011(.A(G381), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  OR4_X1    g1014(.A1(G387), .A2(new_n1214), .A3(G378), .A4(G375), .ZN(G407));
  OAI21_X1  g1015(.A(new_n1118), .B1(new_n1086), .B2(new_n682), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n1081), .B2(new_n1088), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n616), .A2(G213), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  OAI211_X1 g1020(.A(G407), .B(G213), .C1(G375), .C2(new_n1220), .ZN(G409));
  NAND2_X1  g1021(.A1(G387), .A2(new_n1211), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n949), .B1(new_n947), .B2(new_n677), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n968), .B(new_n966), .C1(new_n1223), .C2(new_n683), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1224), .A2(new_n921), .A3(G390), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1222), .A2(KEYINPUT125), .A3(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(G393), .B(G396), .ZN(new_n1227));
  AOI21_X1  g1027(.A(G390), .B1(new_n1224), .B2(new_n921), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT125), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1227), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1226), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1222), .A2(new_n1227), .A3(new_n1225), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT126), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1222), .A2(KEYINPUT126), .A3(new_n1227), .A4(new_n1225), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1231), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G378), .B(new_n1172), .C1(new_n1178), .C2(new_n1181), .ZN(new_n1237));
  AND4_X1   g1037(.A1(new_n950), .A2(new_n1177), .A3(new_n1144), .A4(new_n1133), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1217), .B1(new_n1238), .B2(new_n1171), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1176), .A2(KEYINPUT60), .A3(new_n1068), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT60), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1208), .A2(new_n1242), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1241), .A2(new_n679), .A3(new_n1087), .A4(new_n1243), .ZN(new_n1244));
  OR2_X1    g1044(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1204), .A2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1244), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1244), .A2(new_n1246), .A3(new_n1248), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1240), .A2(new_n1218), .A3(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT63), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1219), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(KEYINPUT63), .A3(new_n1252), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1240), .A2(new_n1218), .ZN(new_n1258));
  AND3_X1   g1058(.A1(new_n1244), .A2(new_n1246), .A3(new_n1248), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1248), .B1(new_n1244), .B2(new_n1246), .ZN(new_n1260));
  INV_X1    g1060(.A(G2897), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n1259), .A2(new_n1260), .B1(new_n1261), .B2(new_n1218), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1218), .A2(new_n1261), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1250), .A2(new_n1251), .A3(new_n1263), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT61), .B1(new_n1258), .B2(new_n1265), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1236), .A2(new_n1255), .A3(new_n1257), .A4(new_n1266), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1231), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT61), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1269), .B1(new_n1256), .B2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT62), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1253), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1256), .A2(KEYINPUT62), .A3(new_n1252), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1271), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1268), .B1(new_n1275), .B2(KEYINPUT127), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1274), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT62), .B1(new_n1256), .B2(new_n1252), .ZN(new_n1278));
  OAI211_X1 g1078(.A(KEYINPUT127), .B(new_n1266), .C1(new_n1277), .C2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1267), .B1(new_n1276), .B2(new_n1280), .ZN(G405));
  XNOR2_X1  g1081(.A(G375), .B(G378), .ZN(new_n1282));
  XNOR2_X1  g1082(.A(new_n1282), .B(new_n1252), .ZN(new_n1283));
  XNOR2_X1  g1083(.A(new_n1283), .B(new_n1236), .ZN(G402));
endmodule


