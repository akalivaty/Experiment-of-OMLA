

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U550 ( .A(n717), .B(KEYINPUT29), .Z(n514) );
  OR2_X1 U551 ( .A1(n790), .A2(G1966), .ZN(n679) );
  XNOR2_X1 U552 ( .A(n679), .B(KEYINPUT96), .ZN(n737) );
  NAND2_X1 U553 ( .A1(n754), .A2(n753), .ZN(n719) );
  AND2_X1 U554 ( .A1(n793), .A2(n742), .ZN(n748) );
  NOR2_X1 U555 ( .A1(n752), .A2(n751), .ZN(n786) );
  XNOR2_X1 U556 ( .A(n678), .B(n677), .ZN(n753) );
  INV_X1 U557 ( .A(KEYINPUT103), .ZN(n810) );
  NOR2_X1 U558 ( .A1(G543), .A2(G651), .ZN(n629) );
  XNOR2_X1 U559 ( .A(n811), .B(n810), .ZN(n825) );
  XOR2_X1 U560 ( .A(KEYINPUT1), .B(n525), .Z(n628) );
  NAND2_X1 U561 ( .A1(n825), .A2(n824), .ZN(n826) );
  NOR2_X1 U562 ( .A1(n524), .A2(n523), .ZN(n676) );
  BUF_X1 U563 ( .A(n676), .Z(G160) );
  NOR2_X1 U564 ( .A1(G2104), .A2(G2105), .ZN(n515) );
  XOR2_X2 U565 ( .A(KEYINPUT17), .B(n515), .Z(n879) );
  NAND2_X1 U566 ( .A1(n879), .A2(G137), .ZN(n517) );
  AND2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n876) );
  NAND2_X1 U568 ( .A1(n876), .A2(G113), .ZN(n516) );
  NAND2_X1 U569 ( .A1(n517), .A2(n516), .ZN(n524) );
  AND2_X1 U570 ( .A1(G2104), .A2(G101), .ZN(n518) );
  INV_X1 U571 ( .A(G2105), .ZN(n540) );
  NAND2_X1 U572 ( .A1(n518), .A2(n540), .ZN(n519) );
  XOR2_X1 U573 ( .A(KEYINPUT23), .B(n519), .Z(n521) );
  NOR2_X2 U574 ( .A1(G2104), .A2(n540), .ZN(n875) );
  NAND2_X1 U575 ( .A1(n875), .A2(G125), .ZN(n520) );
  NAND2_X1 U576 ( .A1(n521), .A2(n520), .ZN(n522) );
  XOR2_X1 U577 ( .A(KEYINPUT65), .B(n522), .Z(n523) );
  XOR2_X1 U578 ( .A(G651), .B(KEYINPUT66), .Z(n529) );
  NOR2_X1 U579 ( .A1(G543), .A2(n529), .ZN(n525) );
  NAND2_X1 U580 ( .A1(G64), .A2(n628), .ZN(n528) );
  XOR2_X1 U581 ( .A(G543), .B(KEYINPUT0), .Z(n622) );
  NOR2_X1 U582 ( .A1(G651), .A2(n622), .ZN(n526) );
  XNOR2_X1 U583 ( .A(KEYINPUT64), .B(n526), .ZN(n630) );
  NAND2_X1 U584 ( .A1(G52), .A2(n630), .ZN(n527) );
  NAND2_X1 U585 ( .A1(n528), .A2(n527), .ZN(n534) );
  NOR2_X1 U586 ( .A1(n622), .A2(n529), .ZN(n633) );
  NAND2_X1 U587 ( .A1(G77), .A2(n633), .ZN(n531) );
  NAND2_X1 U588 ( .A1(G90), .A2(n629), .ZN(n530) );
  NAND2_X1 U589 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U590 ( .A(KEYINPUT9), .B(n532), .Z(n533) );
  NOR2_X1 U591 ( .A1(n534), .A2(n533), .ZN(G171) );
  INV_X1 U592 ( .A(G171), .ZN(G301) );
  AND2_X1 U593 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U594 ( .A1(G111), .A2(n876), .ZN(n535) );
  XNOR2_X1 U595 ( .A(n535), .B(KEYINPUT76), .ZN(n539) );
  XOR2_X1 U596 ( .A(KEYINPUT75), .B(KEYINPUT18), .Z(n537) );
  NAND2_X1 U597 ( .A1(G123), .A2(n875), .ZN(n536) );
  XNOR2_X1 U598 ( .A(n537), .B(n536), .ZN(n538) );
  NAND2_X1 U599 ( .A1(n539), .A2(n538), .ZN(n544) );
  AND2_X1 U600 ( .A1(n540), .A2(G2104), .ZN(n881) );
  NAND2_X1 U601 ( .A1(G99), .A2(n881), .ZN(n542) );
  NAND2_X1 U602 ( .A1(G135), .A2(n879), .ZN(n541) );
  NAND2_X1 U603 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U604 ( .A1(n544), .A2(n543), .ZN(n975) );
  XNOR2_X1 U605 ( .A(n975), .B(G2096), .ZN(n545) );
  XNOR2_X1 U606 ( .A(n545), .B(KEYINPUT77), .ZN(n546) );
  OR2_X1 U607 ( .A1(G2100), .A2(n546), .ZN(G156) );
  INV_X1 U608 ( .A(G57), .ZN(G237) );
  NAND2_X1 U609 ( .A1(n629), .A2(G89), .ZN(n547) );
  XNOR2_X1 U610 ( .A(n547), .B(KEYINPUT4), .ZN(n549) );
  NAND2_X1 U611 ( .A1(G76), .A2(n633), .ZN(n548) );
  NAND2_X1 U612 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U613 ( .A(KEYINPUT5), .B(n550), .ZN(n557) );
  XNOR2_X1 U614 ( .A(KEYINPUT74), .B(KEYINPUT6), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n628), .A2(G63), .ZN(n553) );
  NAND2_X1 U616 ( .A1(G51), .A2(n630), .ZN(n551) );
  XOR2_X1 U617 ( .A(KEYINPUT73), .B(n551), .Z(n552) );
  NAND2_X1 U618 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U619 ( .A(n555), .B(n554), .Z(n556) );
  NAND2_X1 U620 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U621 ( .A(KEYINPUT7), .B(n558), .ZN(G168) );
  XOR2_X1 U622 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U623 ( .A1(G7), .A2(G661), .ZN(n559) );
  XOR2_X1 U624 ( .A(n559), .B(KEYINPUT10), .Z(n838) );
  NAND2_X1 U625 ( .A1(n838), .A2(G567), .ZN(n560) );
  XOR2_X1 U626 ( .A(KEYINPUT11), .B(n560), .Z(G234) );
  NAND2_X1 U627 ( .A1(n628), .A2(G56), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(KEYINPUT14), .ZN(n563) );
  NAND2_X1 U629 ( .A1(G43), .A2(n630), .ZN(n562) );
  NAND2_X1 U630 ( .A1(n563), .A2(n562), .ZN(n569) );
  NAND2_X1 U631 ( .A1(n629), .A2(G81), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(KEYINPUT12), .ZN(n566) );
  NAND2_X1 U633 ( .A1(G68), .A2(n633), .ZN(n565) );
  NAND2_X1 U634 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U635 ( .A(KEYINPUT13), .B(n567), .Z(n568) );
  NOR2_X1 U636 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U637 ( .A(KEYINPUT71), .B(n570), .Z(n924) );
  INV_X1 U638 ( .A(n924), .ZN(n700) );
  INV_X1 U639 ( .A(n700), .ZN(n647) );
  NAND2_X1 U640 ( .A1(n647), .A2(G860), .ZN(n571) );
  XNOR2_X1 U641 ( .A(KEYINPUT72), .B(n571), .ZN(G153) );
  NAND2_X1 U642 ( .A1(G868), .A2(G301), .ZN(n580) );
  NAND2_X1 U643 ( .A1(G66), .A2(n628), .ZN(n573) );
  NAND2_X1 U644 ( .A1(G54), .A2(n630), .ZN(n572) );
  NAND2_X1 U645 ( .A1(n573), .A2(n572), .ZN(n577) );
  NAND2_X1 U646 ( .A1(G79), .A2(n633), .ZN(n575) );
  NAND2_X1 U647 ( .A1(G92), .A2(n629), .ZN(n574) );
  NAND2_X1 U648 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U649 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U650 ( .A(KEYINPUT15), .B(n578), .ZN(n923) );
  INV_X1 U651 ( .A(G868), .ZN(n651) );
  NAND2_X1 U652 ( .A1(n923), .A2(n651), .ZN(n579) );
  NAND2_X1 U653 ( .A1(n580), .A2(n579), .ZN(G284) );
  NAND2_X1 U654 ( .A1(G53), .A2(n630), .ZN(n581) );
  XOR2_X1 U655 ( .A(KEYINPUT69), .B(n581), .Z(n583) );
  NAND2_X1 U656 ( .A1(n628), .A2(G65), .ZN(n582) );
  NAND2_X1 U657 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U658 ( .A(KEYINPUT70), .B(n584), .Z(n588) );
  NAND2_X1 U659 ( .A1(n633), .A2(G78), .ZN(n586) );
  NAND2_X1 U660 ( .A1(G91), .A2(n629), .ZN(n585) );
  AND2_X1 U661 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U662 ( .A1(n588), .A2(n587), .ZN(G299) );
  NOR2_X1 U663 ( .A1(G286), .A2(n651), .ZN(n590) );
  NOR2_X1 U664 ( .A1(G868), .A2(G299), .ZN(n589) );
  NOR2_X1 U665 ( .A1(n590), .A2(n589), .ZN(G297) );
  INV_X1 U666 ( .A(G559), .ZN(n593) );
  NOR2_X1 U667 ( .A1(G860), .A2(n593), .ZN(n591) );
  NOR2_X1 U668 ( .A1(n923), .A2(n591), .ZN(n592) );
  XOR2_X1 U669 ( .A(KEYINPUT16), .B(n592), .Z(G148) );
  INV_X1 U670 ( .A(n923), .ZN(n708) );
  NAND2_X1 U671 ( .A1(n593), .A2(n708), .ZN(n594) );
  NAND2_X1 U672 ( .A1(n594), .A2(G868), .ZN(n596) );
  NAND2_X1 U673 ( .A1(n700), .A2(n651), .ZN(n595) );
  NAND2_X1 U674 ( .A1(n596), .A2(n595), .ZN(G282) );
  NAND2_X1 U675 ( .A1(n708), .A2(G559), .ZN(n649) );
  XOR2_X1 U676 ( .A(n647), .B(n649), .Z(n597) );
  NOR2_X1 U677 ( .A1(n597), .A2(G860), .ZN(n604) );
  NAND2_X1 U678 ( .A1(G67), .A2(n628), .ZN(n599) );
  NAND2_X1 U679 ( .A1(G55), .A2(n630), .ZN(n598) );
  NAND2_X1 U680 ( .A1(n599), .A2(n598), .ZN(n603) );
  NAND2_X1 U681 ( .A1(G80), .A2(n633), .ZN(n601) );
  NAND2_X1 U682 ( .A1(G93), .A2(n629), .ZN(n600) );
  NAND2_X1 U683 ( .A1(n601), .A2(n600), .ZN(n602) );
  OR2_X1 U684 ( .A1(n603), .A2(n602), .ZN(n652) );
  XOR2_X1 U685 ( .A(n604), .B(n652), .Z(G145) );
  NAND2_X1 U686 ( .A1(G73), .A2(n633), .ZN(n605) );
  XNOR2_X1 U687 ( .A(n605), .B(KEYINPUT2), .ZN(n612) );
  NAND2_X1 U688 ( .A1(G61), .A2(n628), .ZN(n607) );
  NAND2_X1 U689 ( .A1(G86), .A2(n629), .ZN(n606) );
  NAND2_X1 U690 ( .A1(n607), .A2(n606), .ZN(n610) );
  NAND2_X1 U691 ( .A1(G48), .A2(n630), .ZN(n608) );
  XNOR2_X1 U692 ( .A(KEYINPUT79), .B(n608), .ZN(n609) );
  NOR2_X1 U693 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U694 ( .A1(n612), .A2(n611), .ZN(G305) );
  NAND2_X1 U695 ( .A1(G75), .A2(n633), .ZN(n614) );
  NAND2_X1 U696 ( .A1(G88), .A2(n629), .ZN(n613) );
  NAND2_X1 U697 ( .A1(n614), .A2(n613), .ZN(n620) );
  NAND2_X1 U698 ( .A1(G62), .A2(n628), .ZN(n615) );
  XNOR2_X1 U699 ( .A(n615), .B(KEYINPUT80), .ZN(n618) );
  NAND2_X1 U700 ( .A1(n630), .A2(G50), .ZN(n616) );
  XOR2_X1 U701 ( .A(KEYINPUT81), .B(n616), .Z(n617) );
  NAND2_X1 U702 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U703 ( .A1(n620), .A2(n619), .ZN(G166) );
  NAND2_X1 U704 ( .A1(G74), .A2(G651), .ZN(n621) );
  XNOR2_X1 U705 ( .A(n621), .B(KEYINPUT78), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n622), .A2(G87), .ZN(n624) );
  NAND2_X1 U707 ( .A1(G49), .A2(n630), .ZN(n623) );
  NAND2_X1 U708 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U709 ( .A1(n628), .A2(n625), .ZN(n626) );
  NAND2_X1 U710 ( .A1(n627), .A2(n626), .ZN(G288) );
  NAND2_X1 U711 ( .A1(n628), .A2(G60), .ZN(n638) );
  NAND2_X1 U712 ( .A1(n629), .A2(G85), .ZN(n632) );
  NAND2_X1 U713 ( .A1(G47), .A2(n630), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U715 ( .A1(G72), .A2(n633), .ZN(n634) );
  XNOR2_X1 U716 ( .A(KEYINPUT67), .B(n634), .ZN(n635) );
  NOR2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U719 ( .A(n639), .B(KEYINPUT68), .ZN(G290) );
  XNOR2_X1 U720 ( .A(KEYINPUT19), .B(KEYINPUT82), .ZN(n641) );
  XNOR2_X1 U721 ( .A(G288), .B(KEYINPUT83), .ZN(n640) );
  XNOR2_X1 U722 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U723 ( .A(n642), .B(n652), .ZN(n644) );
  XOR2_X1 U724 ( .A(G290), .B(G299), .Z(n643) );
  XNOR2_X1 U725 ( .A(n644), .B(n643), .ZN(n645) );
  XOR2_X1 U726 ( .A(G166), .B(n645), .Z(n646) );
  XNOR2_X1 U727 ( .A(G305), .B(n646), .ZN(n648) );
  XOR2_X1 U728 ( .A(n648), .B(n647), .Z(n910) );
  XOR2_X1 U729 ( .A(n910), .B(n649), .Z(n650) );
  NAND2_X1 U730 ( .A1(G868), .A2(n650), .ZN(n654) );
  NAND2_X1 U731 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U732 ( .A1(n654), .A2(n653), .ZN(G295) );
  NAND2_X1 U733 ( .A1(G2078), .A2(G2084), .ZN(n655) );
  XOR2_X1 U734 ( .A(KEYINPUT20), .B(n655), .Z(n656) );
  NAND2_X1 U735 ( .A1(G2090), .A2(n656), .ZN(n657) );
  XNOR2_X1 U736 ( .A(KEYINPUT21), .B(n657), .ZN(n658) );
  NAND2_X1 U737 ( .A1(n658), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U738 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U739 ( .A1(G120), .A2(G69), .ZN(n659) );
  NOR2_X1 U740 ( .A1(G237), .A2(n659), .ZN(n660) );
  NAND2_X1 U741 ( .A1(G108), .A2(n660), .ZN(n843) );
  NAND2_X1 U742 ( .A1(G567), .A2(n843), .ZN(n667) );
  NAND2_X1 U743 ( .A1(G132), .A2(G82), .ZN(n661) );
  XNOR2_X1 U744 ( .A(n661), .B(KEYINPUT22), .ZN(n662) );
  XNOR2_X1 U745 ( .A(n662), .B(KEYINPUT84), .ZN(n663) );
  NOR2_X1 U746 ( .A1(G218), .A2(n663), .ZN(n664) );
  XOR2_X1 U747 ( .A(KEYINPUT85), .B(n664), .Z(n665) );
  NAND2_X1 U748 ( .A1(G96), .A2(n665), .ZN(n842) );
  NAND2_X1 U749 ( .A1(G2106), .A2(n842), .ZN(n666) );
  NAND2_X1 U750 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U751 ( .A(KEYINPUT86), .B(n668), .ZN(n922) );
  NAND2_X1 U752 ( .A1(G661), .A2(G483), .ZN(n669) );
  NOR2_X1 U753 ( .A1(n922), .A2(n669), .ZN(n841) );
  NAND2_X1 U754 ( .A1(n841), .A2(G36), .ZN(G176) );
  NAND2_X1 U755 ( .A1(G102), .A2(n881), .ZN(n671) );
  NAND2_X1 U756 ( .A1(G138), .A2(n879), .ZN(n670) );
  NAND2_X1 U757 ( .A1(n671), .A2(n670), .ZN(n675) );
  NAND2_X1 U758 ( .A1(G126), .A2(n875), .ZN(n673) );
  NAND2_X1 U759 ( .A1(G114), .A2(n876), .ZN(n672) );
  NAND2_X1 U760 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U761 ( .A1(n675), .A2(n674), .ZN(G164) );
  XNOR2_X1 U762 ( .A(KEYINPUT87), .B(G166), .ZN(G303) );
  NOR2_X1 U763 ( .A1(G164), .A2(G1384), .ZN(n754) );
  NAND2_X1 U764 ( .A1(G40), .A2(n676), .ZN(n678) );
  INV_X1 U765 ( .A(KEYINPUT88), .ZN(n677) );
  NAND2_X1 U766 ( .A1(G8), .A2(n719), .ZN(n790) );
  INV_X1 U767 ( .A(G8), .ZN(n680) );
  NOR2_X1 U768 ( .A1(G2084), .A2(n719), .ZN(n735) );
  NOR2_X1 U769 ( .A1(n680), .A2(n735), .ZN(n681) );
  AND2_X1 U770 ( .A1(n737), .A2(n681), .ZN(n682) );
  XOR2_X1 U771 ( .A(KEYINPUT30), .B(n682), .Z(n683) );
  NOR2_X1 U772 ( .A1(G168), .A2(n683), .ZN(n687) );
  XNOR2_X1 U773 ( .A(KEYINPUT25), .B(G2078), .ZN(n1000) );
  NOR2_X1 U774 ( .A1(n719), .A2(n1000), .ZN(n685) );
  INV_X1 U775 ( .A(n719), .ZN(n701) );
  INV_X1 U776 ( .A(G1961), .ZN(n929) );
  NOR2_X1 U777 ( .A1(n701), .A2(n929), .ZN(n684) );
  NOR2_X1 U778 ( .A1(n685), .A2(n684), .ZN(n690) );
  NOR2_X1 U779 ( .A1(G171), .A2(n690), .ZN(n686) );
  NOR2_X1 U780 ( .A1(n687), .A2(n686), .ZN(n688) );
  XNOR2_X1 U781 ( .A(n688), .B(KEYINPUT99), .ZN(n689) );
  XNOR2_X1 U782 ( .A(n689), .B(KEYINPUT31), .ZN(n733) );
  NAND2_X1 U783 ( .A1(G171), .A2(n690), .ZN(n718) );
  INV_X1 U784 ( .A(G299), .ZN(n712) );
  NAND2_X1 U785 ( .A1(n719), .A2(G1956), .ZN(n693) );
  NAND2_X1 U786 ( .A1(n701), .A2(G2072), .ZN(n691) );
  XOR2_X1 U787 ( .A(KEYINPUT27), .B(n691), .Z(n692) );
  NAND2_X1 U788 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U789 ( .A(n694), .B(KEYINPUT97), .ZN(n711) );
  NOR2_X1 U790 ( .A1(n712), .A2(n711), .ZN(n695) );
  XOR2_X1 U791 ( .A(n695), .B(KEYINPUT28), .Z(n716) );
  INV_X1 U792 ( .A(G1996), .ZN(n899) );
  NOR2_X1 U793 ( .A1(n719), .A2(n899), .ZN(n696) );
  XOR2_X1 U794 ( .A(n696), .B(KEYINPUT26), .Z(n698) );
  NAND2_X1 U795 ( .A1(n719), .A2(G1341), .ZN(n697) );
  NAND2_X1 U796 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U797 ( .A1(n700), .A2(n699), .ZN(n707) );
  NAND2_X1 U798 ( .A1(n708), .A2(n707), .ZN(n706) );
  AND2_X1 U799 ( .A1(n701), .A2(G2067), .ZN(n702) );
  XOR2_X1 U800 ( .A(n702), .B(KEYINPUT98), .Z(n704) );
  NAND2_X1 U801 ( .A1(n719), .A2(G1348), .ZN(n703) );
  NAND2_X1 U802 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U803 ( .A1(n706), .A2(n705), .ZN(n710) );
  OR2_X1 U804 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U805 ( .A1(n710), .A2(n709), .ZN(n714) );
  NAND2_X1 U806 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U807 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U808 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U809 ( .A1(n718), .A2(n514), .ZN(n734) );
  NOR2_X1 U810 ( .A1(G2090), .A2(n719), .ZN(n720) );
  XOR2_X1 U811 ( .A(KEYINPUT101), .B(n720), .Z(n723) );
  NOR2_X1 U812 ( .A1(G1971), .A2(n790), .ZN(n721) );
  XNOR2_X1 U813 ( .A(KEYINPUT100), .B(n721), .ZN(n722) );
  NOR2_X1 U814 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U815 ( .A1(n724), .A2(G303), .ZN(n725) );
  OR2_X1 U816 ( .A1(n680), .A2(n725), .ZN(n727) );
  AND2_X1 U817 ( .A1(n734), .A2(n727), .ZN(n726) );
  NAND2_X1 U818 ( .A1(n733), .A2(n726), .ZN(n731) );
  INV_X1 U819 ( .A(n727), .ZN(n729) );
  AND2_X1 U820 ( .A1(G286), .A2(G8), .ZN(n728) );
  OR2_X1 U821 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U822 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U823 ( .A(n732), .B(KEYINPUT32), .ZN(n793) );
  NAND2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n739) );
  NAND2_X1 U825 ( .A1(G8), .A2(n735), .ZN(n736) );
  AND2_X1 U826 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U827 ( .A1(n739), .A2(n738), .ZN(n791) );
  NAND2_X1 U828 ( .A1(G1976), .A2(G288), .ZN(n927) );
  INV_X1 U829 ( .A(n927), .ZN(n740) );
  OR2_X1 U830 ( .A1(n790), .A2(n740), .ZN(n744) );
  INV_X1 U831 ( .A(n744), .ZN(n741) );
  AND2_X1 U832 ( .A1(n791), .A2(n741), .ZN(n742) );
  NOR2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n749) );
  NOR2_X1 U834 ( .A1(G1971), .A2(G303), .ZN(n743) );
  NOR2_X1 U835 ( .A1(n749), .A2(n743), .ZN(n933) );
  OR2_X1 U836 ( .A1(n744), .A2(n933), .ZN(n746) );
  INV_X1 U837 ( .A(KEYINPUT33), .ZN(n745) );
  NAND2_X1 U838 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U839 ( .A1(n748), .A2(n747), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n749), .A2(KEYINPUT33), .ZN(n750) );
  NOR2_X1 U841 ( .A1(n790), .A2(n750), .ZN(n751) );
  XOR2_X1 U842 ( .A(G1981), .B(G305), .Z(n938) );
  INV_X1 U843 ( .A(n753), .ZN(n755) );
  NOR2_X1 U844 ( .A1(n755), .A2(n754), .ZN(n822) );
  XNOR2_X1 U845 ( .A(G2067), .B(KEYINPUT37), .ZN(n820) );
  NAND2_X1 U846 ( .A1(n881), .A2(G104), .ZN(n756) );
  XNOR2_X1 U847 ( .A(KEYINPUT89), .B(n756), .ZN(n759) );
  NAND2_X1 U848 ( .A1(n879), .A2(G140), .ZN(n757) );
  XOR2_X1 U849 ( .A(KEYINPUT90), .B(n757), .Z(n758) );
  NOR2_X1 U850 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U851 ( .A(KEYINPUT34), .B(n760), .ZN(n766) );
  NAND2_X1 U852 ( .A1(n875), .A2(G128), .ZN(n761) );
  XOR2_X1 U853 ( .A(KEYINPUT91), .B(n761), .Z(n763) );
  NAND2_X1 U854 ( .A1(n876), .A2(G116), .ZN(n762) );
  NAND2_X1 U855 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U856 ( .A(KEYINPUT35), .B(n764), .ZN(n765) );
  NAND2_X1 U857 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U858 ( .A(n767), .B(KEYINPUT36), .ZN(n768) );
  XOR2_X1 U859 ( .A(KEYINPUT92), .B(n768), .Z(n868) );
  OR2_X1 U860 ( .A1(n820), .A2(n868), .ZN(n769) );
  XNOR2_X1 U861 ( .A(KEYINPUT93), .B(n769), .ZN(n994) );
  NAND2_X1 U862 ( .A1(n822), .A2(n994), .ZN(n818) );
  NAND2_X1 U863 ( .A1(G119), .A2(n875), .ZN(n771) );
  NAND2_X1 U864 ( .A1(G107), .A2(n876), .ZN(n770) );
  NAND2_X1 U865 ( .A1(n771), .A2(n770), .ZN(n775) );
  NAND2_X1 U866 ( .A1(G95), .A2(n881), .ZN(n773) );
  NAND2_X1 U867 ( .A1(G131), .A2(n879), .ZN(n772) );
  NAND2_X1 U868 ( .A1(n773), .A2(n772), .ZN(n774) );
  NOR2_X1 U869 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U870 ( .A(KEYINPUT94), .B(n776), .Z(n867) );
  AND2_X1 U871 ( .A1(G1991), .A2(n867), .ZN(n978) );
  NAND2_X1 U872 ( .A1(G129), .A2(n875), .ZN(n778) );
  NAND2_X1 U873 ( .A1(G117), .A2(n876), .ZN(n777) );
  NAND2_X1 U874 ( .A1(n778), .A2(n777), .ZN(n781) );
  NAND2_X1 U875 ( .A1(n881), .A2(G105), .ZN(n779) );
  XOR2_X1 U876 ( .A(KEYINPUT38), .B(n779), .Z(n780) );
  NOR2_X1 U877 ( .A1(n781), .A2(n780), .ZN(n783) );
  NAND2_X1 U878 ( .A1(n879), .A2(G141), .ZN(n782) );
  NAND2_X1 U879 ( .A1(n783), .A2(n782), .ZN(n872) );
  AND2_X1 U880 ( .A1(n872), .A2(G1996), .ZN(n976) );
  OR2_X1 U881 ( .A1(n978), .A2(n976), .ZN(n784) );
  NAND2_X1 U882 ( .A1(n822), .A2(n784), .ZN(n812) );
  AND2_X1 U883 ( .A1(n818), .A2(n812), .ZN(n804) );
  AND2_X1 U884 ( .A1(n938), .A2(n804), .ZN(n785) );
  NAND2_X1 U885 ( .A1(n786), .A2(n785), .ZN(n806) );
  NOR2_X1 U886 ( .A1(G1981), .A2(G305), .ZN(n787) );
  XNOR2_X1 U887 ( .A(n787), .B(KEYINPUT95), .ZN(n788) );
  XNOR2_X1 U888 ( .A(KEYINPUT24), .B(n788), .ZN(n789) );
  NOR2_X1 U889 ( .A1(n790), .A2(n789), .ZN(n796) );
  OR2_X1 U890 ( .A1(n796), .A2(n790), .ZN(n794) );
  AND2_X1 U891 ( .A1(n791), .A2(n794), .ZN(n792) );
  NAND2_X1 U892 ( .A1(n793), .A2(n792), .ZN(n802) );
  INV_X1 U893 ( .A(n794), .ZN(n800) );
  NOR2_X1 U894 ( .A1(G2090), .A2(G303), .ZN(n795) );
  NAND2_X1 U895 ( .A1(G8), .A2(n795), .ZN(n798) );
  INV_X1 U896 ( .A(n796), .ZN(n797) );
  AND2_X1 U897 ( .A1(n798), .A2(n797), .ZN(n799) );
  OR2_X1 U898 ( .A1(n800), .A2(n799), .ZN(n801) );
  NAND2_X1 U899 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U900 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U901 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U902 ( .A(n807), .B(KEYINPUT102), .ZN(n809) );
  XNOR2_X1 U903 ( .A(G290), .B(G1986), .ZN(n935) );
  NAND2_X1 U904 ( .A1(n822), .A2(n935), .ZN(n808) );
  NAND2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n811) );
  NOR2_X1 U906 ( .A1(G1996), .A2(n872), .ZN(n973) );
  INV_X1 U907 ( .A(n812), .ZN(n815) );
  NOR2_X1 U908 ( .A1(G290), .A2(G1986), .ZN(n813) );
  NOR2_X1 U909 ( .A1(G1991), .A2(n867), .ZN(n977) );
  NOR2_X1 U910 ( .A1(n813), .A2(n977), .ZN(n814) );
  NOR2_X1 U911 ( .A1(n815), .A2(n814), .ZN(n816) );
  NOR2_X1 U912 ( .A1(n973), .A2(n816), .ZN(n817) );
  XNOR2_X1 U913 ( .A(KEYINPUT39), .B(n817), .ZN(n819) );
  NAND2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n868), .A2(n820), .ZN(n991) );
  NAND2_X1 U916 ( .A1(n821), .A2(n991), .ZN(n823) );
  NAND2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U918 ( .A(n826), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U919 ( .A(G2446), .B(G2451), .ZN(n836) );
  XOR2_X1 U920 ( .A(G2430), .B(G2443), .Z(n828) );
  XNOR2_X1 U921 ( .A(G2454), .B(G2435), .ZN(n827) );
  XNOR2_X1 U922 ( .A(n828), .B(n827), .ZN(n832) );
  XOR2_X1 U923 ( .A(G2438), .B(KEYINPUT104), .Z(n830) );
  XNOR2_X1 U924 ( .A(G1348), .B(G1341), .ZN(n829) );
  XNOR2_X1 U925 ( .A(n830), .B(n829), .ZN(n831) );
  XOR2_X1 U926 ( .A(n832), .B(n831), .Z(n834) );
  XNOR2_X1 U927 ( .A(G2427), .B(KEYINPUT105), .ZN(n833) );
  XNOR2_X1 U928 ( .A(n834), .B(n833), .ZN(n835) );
  XNOR2_X1 U929 ( .A(n836), .B(n835), .ZN(n837) );
  NAND2_X1 U930 ( .A1(n837), .A2(G14), .ZN(n918) );
  XOR2_X1 U931 ( .A(KEYINPUT106), .B(n918), .Z(G401) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n838), .ZN(G217) );
  INV_X1 U933 ( .A(n838), .ZN(G223) );
  AND2_X1 U934 ( .A1(G15), .A2(G2), .ZN(n839) );
  NAND2_X1 U935 ( .A1(G661), .A2(n839), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U937 ( .A1(n841), .A2(n840), .ZN(G188) );
  XNOR2_X1 U938 ( .A(G96), .B(KEYINPUT107), .ZN(G221) );
  XOR2_X1 U939 ( .A(G69), .B(KEYINPUT108), .Z(G235) );
  NOR2_X1 U941 ( .A1(n843), .A2(n842), .ZN(n844) );
  XOR2_X1 U942 ( .A(KEYINPUT109), .B(n844), .Z(G325) );
  XOR2_X1 U943 ( .A(KEYINPUT110), .B(G325), .Z(G261) );
  INV_X1 U944 ( .A(G132), .ZN(G219) );
  INV_X1 U945 ( .A(G120), .ZN(G236) );
  INV_X1 U946 ( .A(G82), .ZN(G220) );
  XOR2_X1 U947 ( .A(KEYINPUT44), .B(KEYINPUT114), .Z(n846) );
  NAND2_X1 U948 ( .A1(G124), .A2(n875), .ZN(n845) );
  XNOR2_X1 U949 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U950 ( .A(n847), .B(KEYINPUT113), .ZN(n850) );
  NAND2_X1 U951 ( .A1(G100), .A2(n881), .ZN(n848) );
  XOR2_X1 U952 ( .A(KEYINPUT115), .B(n848), .Z(n849) );
  NAND2_X1 U953 ( .A1(n850), .A2(n849), .ZN(n854) );
  NAND2_X1 U954 ( .A1(G112), .A2(n876), .ZN(n852) );
  NAND2_X1 U955 ( .A1(G136), .A2(n879), .ZN(n851) );
  NAND2_X1 U956 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U957 ( .A1(n854), .A2(n853), .ZN(G162) );
  XOR2_X1 U958 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n856) );
  XNOR2_X1 U959 ( .A(G164), .B(G162), .ZN(n855) );
  XNOR2_X1 U960 ( .A(n856), .B(n855), .ZN(n866) );
  NAND2_X1 U961 ( .A1(G103), .A2(n881), .ZN(n858) );
  NAND2_X1 U962 ( .A1(G139), .A2(n879), .ZN(n857) );
  NAND2_X1 U963 ( .A1(n858), .A2(n857), .ZN(n864) );
  NAND2_X1 U964 ( .A1(G127), .A2(n875), .ZN(n860) );
  NAND2_X1 U965 ( .A1(G115), .A2(n876), .ZN(n859) );
  NAND2_X1 U966 ( .A1(n860), .A2(n859), .ZN(n861) );
  XNOR2_X1 U967 ( .A(KEYINPUT117), .B(n861), .ZN(n862) );
  XNOR2_X1 U968 ( .A(KEYINPUT47), .B(n862), .ZN(n863) );
  NOR2_X1 U969 ( .A1(n864), .A2(n863), .ZN(n865) );
  XOR2_X1 U970 ( .A(KEYINPUT118), .B(n865), .Z(n985) );
  XOR2_X1 U971 ( .A(n866), .B(n985), .Z(n870) );
  XNOR2_X1 U972 ( .A(n868), .B(n867), .ZN(n869) );
  XNOR2_X1 U973 ( .A(n870), .B(n869), .ZN(n871) );
  XOR2_X1 U974 ( .A(n871), .B(n975), .Z(n874) );
  XOR2_X1 U975 ( .A(G160), .B(n872), .Z(n873) );
  XNOR2_X1 U976 ( .A(n874), .B(n873), .ZN(n888) );
  NAND2_X1 U977 ( .A1(G130), .A2(n875), .ZN(n878) );
  NAND2_X1 U978 ( .A1(G118), .A2(n876), .ZN(n877) );
  NAND2_X1 U979 ( .A1(n878), .A2(n877), .ZN(n886) );
  NAND2_X1 U980 ( .A1(n879), .A2(G142), .ZN(n880) );
  XNOR2_X1 U981 ( .A(n880), .B(KEYINPUT116), .ZN(n883) );
  NAND2_X1 U982 ( .A1(G106), .A2(n881), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U984 ( .A(n884), .B(KEYINPUT45), .Z(n885) );
  NOR2_X1 U985 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U986 ( .A(n888), .B(n887), .Z(n889) );
  NOR2_X1 U987 ( .A1(G37), .A2(n889), .ZN(G395) );
  XOR2_X1 U988 ( .A(KEYINPUT42), .B(G2090), .Z(n891) );
  XNOR2_X1 U989 ( .A(G2067), .B(G2084), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U991 ( .A(n892), .B(G2100), .Z(n894) );
  XNOR2_X1 U992 ( .A(G2078), .B(G2072), .ZN(n893) );
  XNOR2_X1 U993 ( .A(n894), .B(n893), .ZN(n898) );
  XOR2_X1 U994 ( .A(G2096), .B(KEYINPUT43), .Z(n896) );
  XNOR2_X1 U995 ( .A(G2678), .B(KEYINPUT111), .ZN(n895) );
  XNOR2_X1 U996 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U997 ( .A(n898), .B(n897), .Z(G227) );
  XNOR2_X1 U998 ( .A(G1991), .B(G2474), .ZN(n909) );
  XOR2_X1 U999 ( .A(G1981), .B(G1956), .Z(n901) );
  XOR2_X1 U1000 ( .A(n899), .B(G1966), .Z(n900) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n905) );
  XOR2_X1 U1002 ( .A(G1976), .B(G1971), .Z(n903) );
  XOR2_X1 U1003 ( .A(G1986), .B(n929), .Z(n902) );
  XNOR2_X1 U1004 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1005 ( .A(n905), .B(n904), .Z(n907) );
  XNOR2_X1 U1006 ( .A(KEYINPUT112), .B(KEYINPUT41), .ZN(n906) );
  XNOR2_X1 U1007 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1008 ( .A(n909), .B(n908), .ZN(G229) );
  XOR2_X1 U1009 ( .A(KEYINPUT119), .B(n910), .Z(n912) );
  XOR2_X1 U1010 ( .A(G301), .B(G286), .Z(n911) );
  XNOR2_X1 U1011 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1012 ( .A(n913), .B(n923), .Z(n914) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n914), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(KEYINPUT120), .B(n915), .ZN(G397) );
  NOR2_X1 U1015 ( .A1(G227), .A2(G229), .ZN(n916) );
  XOR2_X1 U1016 ( .A(KEYINPUT49), .B(n916), .Z(n917) );
  NAND2_X1 U1017 ( .A1(n918), .A2(n917), .ZN(n919) );
  NOR2_X1 U1018 ( .A1(G395), .A2(n919), .ZN(n921) );
  NOR2_X1 U1019 ( .A1(n922), .A2(G397), .ZN(n920) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1021 ( .A(G225), .ZN(G308) );
  INV_X1 U1022 ( .A(n922), .ZN(G319) );
  INV_X1 U1023 ( .A(G108), .ZN(G238) );
  INV_X1 U1024 ( .A(G16), .ZN(n969) );
  XOR2_X1 U1025 ( .A(KEYINPUT56), .B(n969), .Z(n947) );
  XNOR2_X1 U1026 ( .A(G1348), .B(n923), .ZN(n926) );
  XOR2_X1 U1027 ( .A(n924), .B(G1341), .Z(n925) );
  NOR2_X1 U1028 ( .A1(n926), .A2(n925), .ZN(n928) );
  NAND2_X1 U1029 ( .A1(n928), .A2(n927), .ZN(n931) );
  XOR2_X1 U1030 ( .A(n929), .B(G301), .Z(n930) );
  NOR2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n937) );
  NAND2_X1 U1032 ( .A1(G1971), .A2(G303), .ZN(n932) );
  NAND2_X1 U1033 ( .A1(n933), .A2(n932), .ZN(n934) );
  NOR2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n944) );
  XOR2_X1 U1036 ( .A(G299), .B(G1956), .Z(n942) );
  XNOR2_X1 U1037 ( .A(G1966), .B(G168), .ZN(n939) );
  NAND2_X1 U1038 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1039 ( .A(n940), .B(KEYINPUT57), .ZN(n941) );
  NAND2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1042 ( .A(KEYINPUT125), .B(n945), .ZN(n946) );
  NAND2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n1026) );
  XOR2_X1 U1044 ( .A(G5), .B(G1961), .Z(n960) );
  XNOR2_X1 U1045 ( .A(G1966), .B(G21), .ZN(n958) );
  XOR2_X1 U1046 ( .A(G1348), .B(KEYINPUT59), .Z(n948) );
  XNOR2_X1 U1047 ( .A(G4), .B(n948), .ZN(n950) );
  XNOR2_X1 U1048 ( .A(G6), .B(G1981), .ZN(n949) );
  NOR2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(G1341), .B(G19), .ZN(n952) );
  XNOR2_X1 U1051 ( .A(G1956), .B(G20), .ZN(n951) );
  NOR2_X1 U1052 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1054 ( .A(n955), .B(KEYINPUT126), .ZN(n956) );
  XNOR2_X1 U1055 ( .A(KEYINPUT60), .B(n956), .ZN(n957) );
  NOR2_X1 U1056 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n967) );
  XNOR2_X1 U1058 ( .A(G1986), .B(G24), .ZN(n962) );
  XNOR2_X1 U1059 ( .A(G1971), .B(G22), .ZN(n961) );
  NOR2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n964) );
  XOR2_X1 U1061 ( .A(G1976), .B(G23), .Z(n963) );
  NAND2_X1 U1062 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1063 ( .A(KEYINPUT58), .B(n965), .ZN(n966) );
  NOR2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1065 ( .A(KEYINPUT61), .B(n968), .ZN(n970) );
  NAND2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1067 ( .A1(n971), .A2(G11), .ZN(n1024) );
  INV_X1 U1068 ( .A(G29), .ZN(n1020) );
  XOR2_X1 U1069 ( .A(G2090), .B(G162), .Z(n972) );
  NOR2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n974) );
  XOR2_X1 U1071 ( .A(KEYINPUT51), .B(n974), .Z(n984) );
  NOR2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n982) );
  XOR2_X1 U1075 ( .A(G160), .B(G2084), .Z(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n990) );
  XOR2_X1 U1078 ( .A(G164), .B(G2078), .Z(n987) );
  XNOR2_X1 U1079 ( .A(G2072), .B(n985), .ZN(n986) );
  NOR2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1081 ( .A(KEYINPUT50), .B(n988), .Z(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n992) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1084 ( .A1(n994), .A2(n993), .ZN(n995) );
  XOR2_X1 U1085 ( .A(KEYINPUT52), .B(n995), .Z(n996) );
  NOR2_X1 U1086 ( .A1(KEYINPUT55), .A2(n996), .ZN(n997) );
  NOR2_X1 U1087 ( .A1(n1020), .A2(n997), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(n998), .B(KEYINPUT121), .ZN(n1022) );
  XOR2_X1 U1089 ( .A(KEYINPUT55), .B(KEYINPUT124), .Z(n1018) );
  XNOR2_X1 U1090 ( .A(G2090), .B(G35), .ZN(n1013) );
  XOR2_X1 U1091 ( .A(G25), .B(G1991), .Z(n999) );
  NAND2_X1 U1092 ( .A1(n999), .A2(G28), .ZN(n1010) );
  XNOR2_X1 U1093 ( .A(G27), .B(n1000), .ZN(n1004) );
  XNOR2_X1 U1094 ( .A(G2067), .B(G26), .ZN(n1002) );
  XNOR2_X1 U1095 ( .A(G33), .B(G2072), .ZN(n1001) );
  NOR2_X1 U1096 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1097 ( .A1(n1004), .A2(n1003), .ZN(n1007) );
  XNOR2_X1 U1098 ( .A(G32), .B(G1996), .ZN(n1005) );
  XNOR2_X1 U1099 ( .A(KEYINPUT122), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1100 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1101 ( .A(n1008), .B(KEYINPUT123), .ZN(n1009) );
  NOR2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XNOR2_X1 U1103 ( .A(KEYINPUT53), .B(n1011), .ZN(n1012) );
  NOR2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1016) );
  XOR2_X1 U1105 ( .A(G2084), .B(G34), .Z(n1014) );
  XNOR2_X1 U1106 ( .A(KEYINPUT54), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1107 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1108 ( .A(n1018), .B(n1017), .ZN(n1019) );
  NAND2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1112 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1113 ( .A(n1027), .B(KEYINPUT62), .ZN(n1028) );
  XOR2_X1 U1114 ( .A(KEYINPUT127), .B(n1028), .Z(G150) );
  INV_X1 U1115 ( .A(G150), .ZN(G311) );
endmodule

