

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764;

  NOR2_X1 U383 ( .A1(n698), .A2(n697), .ZN(n374) );
  NAND2_X1 U384 ( .A1(n692), .A2(n369), .ZN(n639) );
  XNOR2_X1 U385 ( .A(n430), .B(n429), .ZN(n744) );
  INV_X1 U386 ( .A(G953), .ZN(n753) );
  NOR2_X2 U387 ( .A1(n554), .A2(n553), .ZN(n601) );
  NOR2_X2 U388 ( .A1(n631), .A2(n764), .ZN(n596) );
  XNOR2_X2 U389 ( .A(n587), .B(n586), .ZN(n631) );
  AND2_X1 U390 ( .A1(n579), .A2(n578), .ZN(n598) );
  AND2_X1 U391 ( .A1(n397), .A2(n564), .ZN(n396) );
  XNOR2_X1 U392 ( .A(n504), .B(n503), .ZN(n571) );
  NOR2_X1 U393 ( .A1(n659), .A2(G902), .ZN(n504) );
  INV_X2 U394 ( .A(G116), .ZN(n424) );
  NAND2_X1 U395 ( .A1(n688), .A2(n620), .ZN(n373) );
  XNOR2_X2 U396 ( .A(n556), .B(KEYINPUT19), .ZN(n565) );
  NAND2_X2 U397 ( .A1(n574), .A2(n711), .ZN(n556) );
  XNOR2_X1 U398 ( .A(n440), .B(KEYINPUT66), .ZN(n529) );
  AND2_X1 U399 ( .A1(n386), .A2(n760), .ZN(n524) );
  XNOR2_X2 U400 ( .A(n546), .B(n545), .ZN(n688) );
  XNOR2_X2 U401 ( .A(G143), .B(G128), .ZN(n447) );
  XNOR2_X1 U402 ( .A(n439), .B(KEYINPUT0), .ZN(n440) );
  XNOR2_X1 U403 ( .A(n393), .B(KEYINPUT81), .ZN(n582) );
  NAND2_X1 U404 ( .A1(n396), .A2(n394), .ZN(n393) );
  XNOR2_X1 U405 ( .A(n572), .B(n395), .ZN(n394) );
  AND2_X1 U406 ( .A1(n695), .A2(n694), .ZN(n531) );
  NOR2_X1 U407 ( .A1(n677), .A2(n570), .ZN(n406) );
  INV_X1 U408 ( .A(KEYINPUT86), .ZN(n405) );
  XNOR2_X1 U409 ( .A(n628), .B(n403), .ZN(n402) );
  INV_X1 U410 ( .A(KEYINPUT88), .ZN(n403) );
  XNOR2_X1 U411 ( .A(n577), .B(n401), .ZN(n400) );
  INV_X1 U412 ( .A(KEYINPUT87), .ZN(n401) );
  NOR2_X1 U413 ( .A1(n715), .A2(n535), .ZN(n536) );
  XOR2_X1 U414 ( .A(KEYINPUT5), .B(G116), .Z(n492) );
  XNOR2_X1 U415 ( .A(G137), .B(G113), .ZN(n494) );
  NAND2_X1 U416 ( .A1(n391), .A2(n390), .ZN(n459) );
  NAND2_X1 U417 ( .A1(n415), .A2(G146), .ZN(n390) );
  NOR2_X1 U418 ( .A1(G953), .A2(G237), .ZN(n490) );
  XNOR2_X1 U419 ( .A(n498), .B(n497), .ZN(n506) );
  INV_X1 U420 ( .A(G472), .ZN(n503) );
  XNOR2_X1 U421 ( .A(G119), .B(KEYINPUT3), .ZN(n427) );
  XNOR2_X1 U422 ( .A(G113), .B(G104), .ZN(n428) );
  AND2_X1 U423 ( .A1(n370), .A2(n433), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n420), .B(n419), .ZN(n422) );
  XNOR2_X1 U425 ( .A(n474), .B(n473), .ZN(n475) );
  INV_X1 U426 ( .A(KEYINPUT65), .ZN(n473) );
  OR2_X1 U427 ( .A1(n621), .A2(G902), .ZN(n368) );
  AND2_X1 U428 ( .A1(n521), .A2(n384), .ZN(n383) );
  XNOR2_X1 U429 ( .A(n398), .B(KEYINPUT85), .ZN(n578) );
  NAND2_X1 U430 ( .A1(n404), .A2(n399), .ZN(n398) );
  AND2_X1 U431 ( .A1(n402), .A2(n400), .ZN(n399) );
  XNOR2_X1 U432 ( .A(G119), .B(G110), .ZN(n483) );
  XNOR2_X1 U433 ( .A(n418), .B(n417), .ZN(n419) );
  NAND2_X1 U434 ( .A1(G234), .A2(G237), .ZN(n408) );
  AND2_X1 U435 ( .A1(n695), .A2(n363), .ZN(n397) );
  INV_X1 U436 ( .A(KEYINPUT30), .ZN(n395) );
  XNOR2_X1 U437 ( .A(n392), .B(n502), .ZN(n659) );
  XNOR2_X1 U438 ( .A(n506), .B(n499), .ZN(n392) );
  BUF_X1 U439 ( .A(n616), .Z(n752) );
  XNOR2_X1 U440 ( .A(n447), .B(n629), .ZN(n498) );
  XNOR2_X1 U441 ( .A(n459), .B(n389), .ZN(n749) );
  XNOR2_X1 U442 ( .A(KEYINPUT10), .B(KEYINPUT68), .ZN(n389) );
  XNOR2_X1 U443 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U444 ( .A(G107), .B(G104), .ZN(n508) );
  XNOR2_X1 U445 ( .A(n506), .B(n505), .ZN(n751) );
  XNOR2_X1 U446 ( .A(n518), .B(n407), .ZN(n725) );
  XNOR2_X1 U447 ( .A(n619), .B(n618), .ZN(n620) );
  INV_X1 U448 ( .A(KEYINPUT35), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(KEYINPUT32), .ZN(n760) );
  AND2_X1 U450 ( .A1(n582), .A2(n576), .ZN(n628) );
  NOR2_X1 U451 ( .A1(n704), .A2(n534), .ZN(n670) );
  NAND2_X1 U452 ( .A1(n376), .A2(n375), .ZN(n761) );
  INV_X1 U453 ( .A(n383), .ZN(n376) );
  INV_X1 U454 ( .A(n387), .ZN(n673) );
  AND2_X1 U455 ( .A1(n573), .A2(n694), .ZN(n363) );
  XOR2_X1 U456 ( .A(n489), .B(KEYINPUT25), .Z(n364) );
  AND2_X1 U457 ( .A1(n564), .A2(n531), .ZN(n365) );
  INV_X1 U458 ( .A(n522), .ZN(n704) );
  NAND2_X1 U459 ( .A1(n575), .A2(n384), .ZN(n366) );
  XOR2_X1 U460 ( .A(n595), .B(KEYINPUT64), .Z(n367) );
  INV_X2 U461 ( .A(KEYINPUT78), .ZN(n423) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n596), .B(n367), .ZN(n597) );
  XNOR2_X2 U464 ( .A(n368), .B(n364), .ZN(n695) );
  XNOR2_X1 U465 ( .A(n487), .B(n486), .ZN(n621) );
  NAND2_X1 U466 ( .A1(n372), .A2(n371), .ZN(n370) );
  INV_X1 U467 ( .A(KEYINPUT2), .ZN(n371) );
  NAND2_X1 U468 ( .A1(n688), .A2(n614), .ZN(n372) );
  XNOR2_X2 U469 ( .A(n373), .B(KEYINPUT80), .ZN(n692) );
  NAND2_X1 U470 ( .A1(n374), .A2(n547), .ZN(n518) );
  AND2_X1 U471 ( .A1(n374), .A2(n704), .ZN(n707) );
  INV_X1 U472 ( .A(n378), .ZN(n375) );
  NAND2_X1 U473 ( .A1(n380), .A2(n377), .ZN(n386) );
  NAND2_X1 U474 ( .A1(n378), .A2(n387), .ZN(n377) );
  NAND2_X1 U475 ( .A1(n379), .A2(n366), .ZN(n378) );
  NAND2_X1 U476 ( .A1(n382), .A2(n381), .ZN(n379) );
  NAND2_X1 U477 ( .A1(n383), .A2(n387), .ZN(n380) );
  NOR2_X1 U478 ( .A1(n575), .A2(n384), .ZN(n381) );
  INV_X1 U479 ( .A(n521), .ZN(n382) );
  NAND2_X1 U480 ( .A1(n523), .A2(n517), .ZN(n385) );
  NAND2_X1 U481 ( .A1(n523), .A2(n388), .ZN(n387) );
  AND2_X1 U482 ( .A1(n697), .A2(n522), .ZN(n388) );
  NAND2_X1 U483 ( .A1(n416), .A2(G125), .ZN(n391) );
  BUF_X1 U484 ( .A(n688), .Z(n739) );
  OR2_X2 U485 ( .A1(n652), .A2(G902), .ZN(n516) );
  XNOR2_X1 U486 ( .A(KEYINPUT33), .B(KEYINPUT73), .ZN(n407) );
  INV_X1 U487 ( .A(n459), .ZN(n417) );
  INV_X1 U488 ( .A(KEYINPUT77), .ZN(n493) );
  INV_X1 U489 ( .A(KEYINPUT92), .ZN(n618) );
  XNOR2_X1 U490 ( .A(n494), .B(n493), .ZN(n495) );
  INV_X1 U491 ( .A(KEYINPUT99), .ZN(n455) );
  XNOR2_X1 U492 ( .A(n496), .B(n495), .ZN(n499) );
  XNOR2_X1 U493 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U494 ( .A(n422), .B(n421), .ZN(n431) );
  XNOR2_X1 U495 ( .A(n458), .B(n457), .ZN(n462) );
  INV_X1 U496 ( .A(KEYINPUT36), .ZN(n557) );
  XNOR2_X1 U497 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U498 ( .A(n463), .B(n632), .ZN(n464) );
  XNOR2_X1 U499 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U500 ( .A(n465), .B(n464), .ZN(n527) );
  INV_X1 U501 ( .A(KEYINPUT125), .ZN(n626) );
  XNOR2_X1 U502 ( .A(n408), .B(KEYINPUT14), .ZN(n410) );
  NAND2_X1 U503 ( .A1(G952), .A2(n410), .ZN(n724) );
  NOR2_X1 U504 ( .A1(n724), .A2(G953), .ZN(n409) );
  XNOR2_X1 U505 ( .A(n409), .B(KEYINPUT97), .ZN(n551) );
  NOR2_X1 U506 ( .A1(G898), .A2(n753), .ZN(n746) );
  NAND2_X1 U507 ( .A1(G902), .A2(n410), .ZN(n548) );
  INV_X1 U508 ( .A(n548), .ZN(n411) );
  NAND2_X1 U509 ( .A1(n746), .A2(n411), .ZN(n412) );
  NAND2_X1 U510 ( .A1(n551), .A2(n412), .ZN(n438) );
  XOR2_X1 U511 ( .A(KEYINPUT18), .B(KEYINPUT83), .Z(n414) );
  XNOR2_X1 U512 ( .A(KEYINPUT84), .B(KEYINPUT17), .ZN(n413) );
  XNOR2_X1 U513 ( .A(n414), .B(n413), .ZN(n420) );
  NAND2_X1 U514 ( .A1(G224), .A2(n753), .ZN(n418) );
  INV_X1 U515 ( .A(G125), .ZN(n415) );
  INV_X1 U516 ( .A(G146), .ZN(n416) );
  XNOR2_X1 U517 ( .A(KEYINPUT4), .B(G101), .ZN(n500) );
  XNOR2_X1 U518 ( .A(n500), .B(n447), .ZN(n421) );
  XOR2_X1 U519 ( .A(KEYINPUT75), .B(KEYINPUT16), .Z(n426) );
  XNOR2_X2 U520 ( .A(n423), .B(G110), .ZN(n509) );
  XNOR2_X2 U521 ( .A(n424), .B(G107), .ZN(n442) );
  XNOR2_X1 U522 ( .A(n509), .B(n442), .ZN(n425) );
  XNOR2_X1 U523 ( .A(n426), .B(n425), .ZN(n430) );
  XNOR2_X1 U524 ( .A(n427), .B(KEYINPUT71), .ZN(n501) );
  XNOR2_X1 U525 ( .A(n428), .B(G122), .ZN(n454) );
  XNOR2_X1 U526 ( .A(n501), .B(n454), .ZN(n429) );
  XNOR2_X1 U527 ( .A(n431), .B(n744), .ZN(n640) );
  INV_X1 U528 ( .A(KEYINPUT15), .ZN(n432) );
  XNOR2_X1 U529 ( .A(n432), .B(G902), .ZN(n433) );
  INV_X1 U530 ( .A(n433), .ZN(n615) );
  NAND2_X1 U531 ( .A1(n640), .A2(n615), .ZN(n436) );
  OR2_X1 U532 ( .A1(G237), .A2(G902), .ZN(n437) );
  INV_X1 U533 ( .A(n437), .ZN(n434) );
  INV_X1 U534 ( .A(G210), .ZN(n638) );
  NOR2_X1 U535 ( .A1(n434), .A2(n638), .ZN(n435) );
  XNOR2_X2 U536 ( .A(n436), .B(n435), .ZN(n574) );
  NAND2_X1 U537 ( .A1(G214), .A2(n437), .ZN(n711) );
  NAND2_X1 U538 ( .A1(n438), .A2(n565), .ZN(n439) );
  INV_X1 U539 ( .A(n529), .ZN(n472) );
  NAND2_X1 U540 ( .A1(G234), .A2(n753), .ZN(n441) );
  XOR2_X1 U541 ( .A(KEYINPUT8), .B(n441), .Z(n482) );
  NAND2_X1 U542 ( .A1(n482), .A2(G217), .ZN(n446) );
  XOR2_X1 U543 ( .A(KEYINPUT7), .B(n442), .Z(n444) );
  XNOR2_X1 U544 ( .A(G122), .B(KEYINPUT9), .ZN(n443) );
  XNOR2_X1 U545 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U546 ( .A(n446), .B(n445), .ZN(n448) );
  INV_X1 U547 ( .A(G134), .ZN(n629) );
  XNOR2_X1 U548 ( .A(n448), .B(n498), .ZN(n734) );
  INV_X1 U549 ( .A(G902), .ZN(n449) );
  NAND2_X1 U550 ( .A1(n734), .A2(n449), .ZN(n450) );
  XNOR2_X1 U551 ( .A(n450), .B(G478), .ZN(n525) );
  XOR2_X1 U552 ( .A(KEYINPUT12), .B(KEYINPUT100), .Z(n452) );
  XNOR2_X1 U553 ( .A(G140), .B(KEYINPUT11), .ZN(n451) );
  XNOR2_X1 U554 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U555 ( .A(n454), .B(n453), .Z(n458) );
  NAND2_X1 U556 ( .A1(G214), .A2(n490), .ZN(n456) );
  XNOR2_X1 U557 ( .A(KEYINPUT69), .B(G131), .ZN(n497) );
  XOR2_X1 U558 ( .A(G143), .B(n497), .Z(n460) );
  XNOR2_X1 U559 ( .A(n749), .B(n460), .ZN(n461) );
  XNOR2_X1 U560 ( .A(n462), .B(n461), .ZN(n633) );
  NOR2_X1 U561 ( .A1(G902), .A2(n633), .ZN(n465) );
  XNOR2_X1 U562 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n463) );
  INV_X1 U563 ( .A(G475), .ZN(n632) );
  NOR2_X1 U564 ( .A1(n525), .A2(n527), .ZN(n466) );
  XNOR2_X1 U565 ( .A(KEYINPUT103), .B(n466), .ZN(n713) );
  NAND2_X1 U566 ( .A1(G234), .A2(n615), .ZN(n467) );
  XNOR2_X1 U567 ( .A(KEYINPUT20), .B(n467), .ZN(n488) );
  NAND2_X1 U568 ( .A1(n488), .A2(G221), .ZN(n469) );
  INV_X1 U569 ( .A(KEYINPUT21), .ZN(n468) );
  XNOR2_X1 U570 ( .A(n469), .B(n468), .ZN(n694) );
  INV_X1 U571 ( .A(n694), .ZN(n470) );
  NOR2_X1 U572 ( .A1(n713), .A2(n470), .ZN(n471) );
  NAND2_X1 U573 ( .A1(n472), .A2(n471), .ZN(n476) );
  XNOR2_X1 U574 ( .A(KEYINPUT22), .B(KEYINPUT74), .ZN(n474) );
  XNOR2_X1 U575 ( .A(n476), .B(n475), .ZN(n537) );
  XOR2_X1 U576 ( .A(KEYINPUT89), .B(KEYINPUT24), .Z(n478) );
  XNOR2_X1 U577 ( .A(G128), .B(KEYINPUT23), .ZN(n477) );
  XNOR2_X1 U578 ( .A(n478), .B(n477), .ZN(n480) );
  XOR2_X1 U579 ( .A(KEYINPUT82), .B(KEYINPUT72), .Z(n479) );
  XNOR2_X1 U580 ( .A(n749), .B(n481), .ZN(n487) );
  NAND2_X1 U581 ( .A1(n482), .A2(G221), .ZN(n485) );
  XNOR2_X1 U582 ( .A(G140), .B(G137), .ZN(n505) );
  XNOR2_X1 U583 ( .A(n483), .B(n505), .ZN(n484) );
  XNOR2_X1 U584 ( .A(n485), .B(n484), .ZN(n486) );
  NAND2_X1 U585 ( .A1(n488), .A2(G217), .ZN(n489) );
  NOR2_X1 U586 ( .A1(n537), .A2(n695), .ZN(n523) );
  NAND2_X1 U587 ( .A1(n490), .A2(G210), .ZN(n491) );
  XNOR2_X1 U588 ( .A(n492), .B(n491), .ZN(n496) );
  XNOR2_X1 U589 ( .A(n500), .B(G146), .ZN(n512) );
  XNOR2_X1 U590 ( .A(n501), .B(n512), .ZN(n502) );
  XOR2_X1 U591 ( .A(n571), .B(KEYINPUT6), .Z(n547) );
  NAND2_X1 U592 ( .A1(n753), .A2(G227), .ZN(n507) );
  XNOR2_X1 U593 ( .A(n508), .B(n507), .ZN(n510) );
  XNOR2_X1 U594 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U595 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U596 ( .A(n751), .B(n513), .ZN(n652) );
  INV_X1 U597 ( .A(KEYINPUT70), .ZN(n514) );
  XNOR2_X1 U598 ( .A(n514), .B(G469), .ZN(n515) );
  XNOR2_X2 U599 ( .A(n516), .B(n515), .ZN(n589) );
  XNOR2_X2 U600 ( .A(n589), .B(KEYINPUT1), .ZN(n697) );
  NOR2_X1 U601 ( .A1(n547), .A2(n697), .ZN(n517) );
  INV_X1 U602 ( .A(n531), .ZN(n698) );
  OR2_X1 U603 ( .A1(n529), .A2(n725), .ZN(n519) );
  XNOR2_X1 U604 ( .A(KEYINPUT34), .B(n519), .ZN(n521) );
  NAND2_X1 U605 ( .A1(n527), .A2(n525), .ZN(n520) );
  XNOR2_X1 U606 ( .A(n520), .B(KEYINPUT104), .ZN(n575) );
  INV_X1 U607 ( .A(n571), .ZN(n522) );
  XNOR2_X1 U608 ( .A(n524), .B(KEYINPUT44), .ZN(n544) );
  INV_X1 U609 ( .A(n525), .ZN(n526) );
  AND2_X1 U610 ( .A1(n527), .A2(n526), .ZN(n679) );
  INV_X1 U611 ( .A(n679), .ZN(n528) );
  OR2_X1 U612 ( .A1(n527), .A2(n526), .ZN(n611) );
  AND2_X1 U613 ( .A1(n528), .A2(n611), .ZN(n715) );
  INV_X1 U614 ( .A(n529), .ZN(n532) );
  NAND2_X1 U615 ( .A1(n532), .A2(n707), .ZN(n530) );
  XNOR2_X1 U616 ( .A(KEYINPUT31), .B(n530), .ZN(n683) );
  INV_X1 U617 ( .A(n589), .ZN(n564) );
  NAND2_X1 U618 ( .A1(n532), .A2(n365), .ZN(n533) );
  XNOR2_X1 U619 ( .A(n533), .B(KEYINPUT98), .ZN(n534) );
  NOR2_X1 U620 ( .A1(n683), .A2(n670), .ZN(n535) );
  XNOR2_X1 U621 ( .A(KEYINPUT102), .B(n536), .ZN(n542) );
  INV_X1 U622 ( .A(n695), .ZN(n539) );
  OR2_X1 U623 ( .A1(n537), .A2(n547), .ZN(n538) );
  NOR2_X1 U624 ( .A1(n539), .A2(n538), .ZN(n540) );
  NAND2_X1 U625 ( .A1(n540), .A2(n697), .ZN(n665) );
  INV_X1 U626 ( .A(n665), .ZN(n541) );
  NOR2_X1 U627 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U628 ( .A1(n544), .A2(n543), .ZN(n546) );
  XOR2_X1 U629 ( .A(KEYINPUT91), .B(KEYINPUT45), .Z(n545) );
  INV_X1 U630 ( .A(n547), .ZN(n554) );
  NOR2_X1 U631 ( .A1(G900), .A2(n548), .ZN(n549) );
  NAND2_X1 U632 ( .A1(n549), .A2(G953), .ZN(n550) );
  NAND2_X1 U633 ( .A1(n551), .A2(n550), .ZN(n573) );
  NAND2_X1 U634 ( .A1(n694), .A2(n573), .ZN(n552) );
  NOR2_X1 U635 ( .A1(n695), .A2(n552), .ZN(n562) );
  NAND2_X1 U636 ( .A1(n679), .A2(n562), .ZN(n553) );
  XNOR2_X1 U637 ( .A(n601), .B(KEYINPUT107), .ZN(n555) );
  NOR2_X1 U638 ( .A1(n556), .A2(n555), .ZN(n560) );
  XNOR2_X1 U639 ( .A(KEYINPUT94), .B(KEYINPUT108), .ZN(n558) );
  NOR2_X1 U640 ( .A1(n561), .A2(n697), .ZN(n686) );
  AND2_X1 U641 ( .A1(n704), .A2(n562), .ZN(n563) );
  XOR2_X1 U642 ( .A(KEYINPUT28), .B(n563), .Z(n590) );
  NAND2_X1 U643 ( .A1(n565), .A2(n564), .ZN(n566) );
  NOR2_X1 U644 ( .A1(n590), .A2(n566), .ZN(n677) );
  XOR2_X1 U645 ( .A(KEYINPUT67), .B(KEYINPUT47), .Z(n567) );
  NOR2_X1 U646 ( .A1(n715), .A2(n567), .ZN(n568) );
  AND2_X1 U647 ( .A1(n677), .A2(n568), .ZN(n569) );
  NOR2_X1 U648 ( .A1(n686), .A2(n569), .ZN(n579) );
  INV_X1 U649 ( .A(KEYINPUT47), .ZN(n570) );
  NAND2_X1 U650 ( .A1(n571), .A2(n711), .ZN(n572) );
  INV_X1 U651 ( .A(n574), .ZN(n606) );
  NOR2_X1 U652 ( .A1(n575), .A2(n606), .ZN(n576) );
  NAND2_X1 U653 ( .A1(n715), .A2(KEYINPUT47), .ZN(n577) );
  INV_X1 U654 ( .A(KEYINPUT76), .ZN(n580) );
  XNOR2_X1 U655 ( .A(n580), .B(KEYINPUT38), .ZN(n581) );
  XNOR2_X1 U656 ( .A(n574), .B(n581), .ZN(n710) );
  NAND2_X1 U657 ( .A1(n582), .A2(n710), .ZN(n584) );
  INV_X1 U658 ( .A(KEYINPUT39), .ZN(n583) );
  XNOR2_X1 U659 ( .A(n584), .B(n583), .ZN(n610) );
  INV_X1 U660 ( .A(n610), .ZN(n585) );
  NAND2_X1 U661 ( .A1(n585), .A2(n679), .ZN(n587) );
  INV_X1 U662 ( .A(KEYINPUT40), .ZN(n586) );
  NAND2_X1 U663 ( .A1(n711), .A2(n710), .ZN(n714) );
  NOR2_X1 U664 ( .A1(n714), .A2(n713), .ZN(n588) );
  XNOR2_X1 U665 ( .A(n588), .B(KEYINPUT41), .ZN(n726) );
  INV_X1 U666 ( .A(n726), .ZN(n592) );
  NOR2_X1 U667 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U668 ( .A1(n592), .A2(n591), .ZN(n594) );
  INV_X1 U669 ( .A(KEYINPUT42), .ZN(n593) );
  XNOR2_X1 U670 ( .A(n594), .B(n593), .ZN(n764) );
  XNOR2_X1 U671 ( .A(KEYINPUT93), .B(KEYINPUT46), .ZN(n595) );
  NAND2_X1 U672 ( .A1(n598), .A2(n597), .ZN(n600) );
  INV_X1 U673 ( .A(KEYINPUT48), .ZN(n599) );
  XNOR2_X1 U674 ( .A(n600), .B(n599), .ZN(n613) );
  NAND2_X1 U675 ( .A1(n601), .A2(n711), .ZN(n603) );
  INV_X1 U676 ( .A(n697), .ZN(n602) );
  NOR2_X1 U677 ( .A1(n603), .A2(n602), .ZN(n605) );
  XNOR2_X1 U678 ( .A(KEYINPUT43), .B(KEYINPUT105), .ZN(n604) );
  XNOR2_X1 U679 ( .A(n605), .B(n604), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n607), .A2(n606), .ZN(n609) );
  INV_X1 U681 ( .A(KEYINPUT106), .ZN(n608) );
  XNOR2_X1 U682 ( .A(n609), .B(n608), .ZN(n763) );
  INV_X1 U683 ( .A(n611), .ZN(n682) );
  AND2_X1 U684 ( .A1(n585), .A2(n682), .ZN(n630) );
  NOR2_X1 U685 ( .A1(n763), .A2(n630), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n616) );
  XNOR2_X1 U687 ( .A(n752), .B(KEYINPUT79), .ZN(n614) );
  INV_X1 U688 ( .A(n616), .ZN(n617) );
  NAND2_X1 U689 ( .A1(n617), .A2(KEYINPUT2), .ZN(n619) );
  INV_X2 U690 ( .A(n639), .ZN(n733) );
  NAND2_X1 U691 ( .A1(n733), .A2(G217), .ZN(n623) );
  XNOR2_X1 U692 ( .A(n621), .B(KEYINPUT124), .ZN(n622) );
  XNOR2_X1 U693 ( .A(n623), .B(n622), .ZN(n625) );
  INV_X1 U694 ( .A(G952), .ZN(n624) );
  AND2_X1 U695 ( .A1(n624), .A2(G953), .ZN(n738) );
  NOR2_X2 U696 ( .A1(n625), .A2(n738), .ZN(n627) );
  XNOR2_X1 U697 ( .A(n627), .B(n626), .ZN(G66) );
  XOR2_X1 U698 ( .A(G143), .B(n628), .Z(G45) );
  XNOR2_X1 U699 ( .A(n630), .B(n629), .ZN(G36) );
  XOR2_X1 U700 ( .A(G131), .B(n631), .Z(G33) );
  NOR2_X1 U701 ( .A1(n639), .A2(n632), .ZN(n635) );
  XNOR2_X1 U702 ( .A(n633), .B(KEYINPUT59), .ZN(n634) );
  XNOR2_X1 U703 ( .A(n635), .B(n634), .ZN(n636) );
  NOR2_X1 U704 ( .A1(n636), .A2(n738), .ZN(n637) );
  XNOR2_X1 U705 ( .A(n637), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X1 U706 ( .A1(n639), .A2(n638), .ZN(n645) );
  BUF_X1 U707 ( .A(n640), .Z(n643) );
  XNOR2_X1 U708 ( .A(KEYINPUT96), .B(KEYINPUT54), .ZN(n641) );
  XOR2_X1 U709 ( .A(n641), .B(KEYINPUT55), .Z(n642) );
  XNOR2_X1 U710 ( .A(n643), .B(n642), .ZN(n644) );
  XNOR2_X1 U711 ( .A(n645), .B(n644), .ZN(n646) );
  NOR2_X1 U712 ( .A1(n646), .A2(n738), .ZN(n648) );
  XOR2_X1 U713 ( .A(KEYINPUT119), .B(KEYINPUT56), .Z(n647) );
  XNOR2_X1 U714 ( .A(n648), .B(n647), .ZN(G51) );
  NAND2_X1 U715 ( .A1(n733), .A2(G469), .ZN(n654) );
  XNOR2_X1 U716 ( .A(KEYINPUT121), .B(KEYINPUT57), .ZN(n650) );
  XNOR2_X1 U717 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n649) );
  XNOR2_X1 U718 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U719 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U720 ( .A(n654), .B(n653), .ZN(n655) );
  NOR2_X2 U721 ( .A1(n655), .A2(n738), .ZN(n656) );
  XNOR2_X1 U722 ( .A(n656), .B(KEYINPUT122), .ZN(G54) );
  NAND2_X1 U723 ( .A1(n733), .A2(G472), .ZN(n661) );
  XOR2_X1 U724 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n657) );
  XNOR2_X1 U725 ( .A(n657), .B(KEYINPUT62), .ZN(n658) );
  XNOR2_X1 U726 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U727 ( .A(n661), .B(n660), .ZN(n662) );
  NOR2_X2 U728 ( .A1(n662), .A2(n738), .ZN(n664) );
  XNOR2_X1 U729 ( .A(KEYINPUT95), .B(KEYINPUT63), .ZN(n663) );
  XNOR2_X1 U730 ( .A(n664), .B(n663), .ZN(G57) );
  XNOR2_X1 U731 ( .A(G101), .B(n665), .ZN(G3) );
  NAND2_X1 U732 ( .A1(n670), .A2(n679), .ZN(n666) );
  XNOR2_X1 U733 ( .A(n666), .B(G104), .ZN(G6) );
  XOR2_X1 U734 ( .A(KEYINPUT27), .B(KEYINPUT112), .Z(n668) );
  XNOR2_X1 U735 ( .A(G107), .B(KEYINPUT26), .ZN(n667) );
  XNOR2_X1 U736 ( .A(n668), .B(n667), .ZN(n669) );
  XOR2_X1 U737 ( .A(KEYINPUT111), .B(n669), .Z(n672) );
  NAND2_X1 U738 ( .A1(n670), .A2(n682), .ZN(n671) );
  XNOR2_X1 U739 ( .A(n672), .B(n671), .ZN(G9) );
  XNOR2_X1 U740 ( .A(G110), .B(n673), .ZN(n674) );
  XNOR2_X1 U741 ( .A(n674), .B(KEYINPUT113), .ZN(G12) );
  XOR2_X1 U742 ( .A(G128), .B(KEYINPUT29), .Z(n676) );
  NAND2_X1 U743 ( .A1(n677), .A2(n682), .ZN(n675) );
  XNOR2_X1 U744 ( .A(n676), .B(n675), .ZN(G30) );
  NAND2_X1 U745 ( .A1(n677), .A2(n679), .ZN(n678) );
  XNOR2_X1 U746 ( .A(n678), .B(G146), .ZN(G48) );
  NAND2_X1 U747 ( .A1(n683), .A2(n679), .ZN(n680) );
  XNOR2_X1 U748 ( .A(n680), .B(KEYINPUT114), .ZN(n681) );
  XNOR2_X1 U749 ( .A(G113), .B(n681), .ZN(G15) );
  XOR2_X1 U750 ( .A(G116), .B(KEYINPUT115), .Z(n685) );
  NAND2_X1 U751 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U752 ( .A(n685), .B(n684), .ZN(G18) );
  XNOR2_X1 U753 ( .A(G125), .B(n686), .ZN(n687) );
  XNOR2_X1 U754 ( .A(n687), .B(KEYINPUT37), .ZN(G27) );
  INV_X1 U755 ( .A(n752), .ZN(n689) );
  NAND2_X1 U756 ( .A1(n739), .A2(n689), .ZN(n690) );
  NAND2_X1 U757 ( .A1(n690), .A2(n371), .ZN(n691) );
  NAND2_X1 U758 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U759 ( .A(n693), .B(KEYINPUT90), .ZN(n730) );
  NOR2_X1 U760 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U761 ( .A(KEYINPUT49), .B(n696), .ZN(n702) );
  NAND2_X1 U762 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U763 ( .A(n699), .B(KEYINPUT116), .ZN(n700) );
  XNOR2_X1 U764 ( .A(KEYINPUT50), .B(n700), .ZN(n701) );
  NAND2_X1 U765 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U766 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U767 ( .A(KEYINPUT117), .B(n705), .Z(n706) );
  NOR2_X1 U768 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U769 ( .A(KEYINPUT51), .B(n708), .Z(n709) );
  NOR2_X1 U770 ( .A1(n726), .A2(n709), .ZN(n721) );
  NOR2_X1 U771 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U772 ( .A1(n713), .A2(n712), .ZN(n717) );
  NOR2_X1 U773 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U774 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U775 ( .A1(n718), .A2(n725), .ZN(n719) );
  XNOR2_X1 U776 ( .A(n719), .B(KEYINPUT118), .ZN(n720) );
  NOR2_X1 U777 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U778 ( .A(n722), .B(KEYINPUT52), .ZN(n723) );
  NOR2_X1 U779 ( .A1(n724), .A2(n723), .ZN(n728) );
  NOR2_X1 U780 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U781 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U782 ( .A1(n730), .A2(n729), .ZN(n731) );
  NOR2_X1 U783 ( .A1(n731), .A2(G953), .ZN(n732) );
  XNOR2_X1 U784 ( .A(n732), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U785 ( .A1(n733), .A2(G478), .ZN(n736) );
  XNOR2_X1 U786 ( .A(n734), .B(KEYINPUT123), .ZN(n735) );
  XNOR2_X1 U787 ( .A(n736), .B(n735), .ZN(n737) );
  NOR2_X1 U788 ( .A1(n738), .A2(n737), .ZN(G63) );
  NAND2_X1 U789 ( .A1(n753), .A2(n739), .ZN(n743) );
  NAND2_X1 U790 ( .A1(G953), .A2(G224), .ZN(n740) );
  XNOR2_X1 U791 ( .A(KEYINPUT61), .B(n740), .ZN(n741) );
  NAND2_X1 U792 ( .A1(n741), .A2(G898), .ZN(n742) );
  NAND2_X1 U793 ( .A1(n743), .A2(n742), .ZN(n748) );
  XOR2_X1 U794 ( .A(G101), .B(n744), .Z(n745) );
  NOR2_X1 U795 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U796 ( .A(n748), .B(n747), .ZN(G69) );
  XNOR2_X1 U797 ( .A(n749), .B(KEYINPUT4), .ZN(n750) );
  XNOR2_X1 U798 ( .A(n751), .B(n750), .ZN(n755) );
  XNOR2_X1 U799 ( .A(n752), .B(n755), .ZN(n754) );
  NAND2_X1 U800 ( .A1(n754), .A2(n753), .ZN(n759) );
  XNOR2_X1 U801 ( .A(n755), .B(G227), .ZN(n756) );
  NAND2_X1 U802 ( .A1(n756), .A2(G900), .ZN(n757) );
  NAND2_X1 U803 ( .A1(G953), .A2(n757), .ZN(n758) );
  NAND2_X1 U804 ( .A1(n759), .A2(n758), .ZN(G72) );
  XNOR2_X1 U805 ( .A(n760), .B(G119), .ZN(G21) );
  XNOR2_X1 U806 ( .A(G122), .B(KEYINPUT126), .ZN(n762) );
  XNOR2_X1 U807 ( .A(n762), .B(n761), .ZN(G24) );
  XOR2_X1 U808 ( .A(G140), .B(n763), .Z(G42) );
  XOR2_X1 U809 ( .A(G137), .B(n764), .Z(G39) );
endmodule

