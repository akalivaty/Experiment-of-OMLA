//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n817, new_n818, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1022, new_n1023;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT22), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n202), .A3(new_n206), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G226gat), .A2(G233gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n216));
  INV_X1    g015(.A(G183gat), .ZN(new_n217));
  INV_X1    g016(.A(G190gat), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(KEYINPUT23), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT64), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(KEYINPUT23), .A3(new_n228), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n221), .A2(KEYINPUT25), .A3(new_n225), .A4(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT65), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n223), .A2(KEYINPUT23), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n221), .A2(new_n225), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT25), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n224), .B1(new_n219), .B2(new_n220), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n236), .A2(new_n237), .A3(KEYINPUT25), .A4(new_n229), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n231), .A2(new_n235), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(KEYINPUT27), .B(G183gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(KEYINPUT28), .A3(new_n218), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(KEYINPUT66), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n240), .A2(new_n243), .A3(KEYINPUT28), .A4(new_n218), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n240), .A2(new_n218), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n242), .B(new_n244), .C1(KEYINPUT28), .C2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT26), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n227), .A2(new_n247), .A3(new_n228), .ZN(new_n248));
  INV_X1    g047(.A(new_n222), .ZN(new_n249));
  INV_X1    g048(.A(new_n223), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n249), .B1(new_n250), .B2(KEYINPUT26), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n248), .A2(new_n251), .B1(G183gat), .B2(G190gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n239), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT29), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n215), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n214), .B1(new_n239), .B2(new_n253), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n213), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT88), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n254), .A2(new_n215), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT29), .B1(new_n239), .B2(new_n253), .ZN(new_n261));
  OAI211_X1 g060(.A(new_n260), .B(new_n212), .C1(new_n215), .C2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n258), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT37), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT38), .ZN(new_n265));
  XNOR2_X1  g064(.A(G8gat), .B(G36gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(new_n266), .B(KEYINPUT73), .ZN(new_n267));
  XNOR2_X1  g066(.A(G64gat), .B(G92gat), .ZN(new_n268));
  XOR2_X1   g067(.A(new_n267), .B(new_n268), .Z(new_n269));
  INV_X1    g068(.A(KEYINPUT37), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n258), .A2(new_n259), .A3(new_n262), .A4(new_n270), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n264), .A2(new_n265), .A3(new_n269), .A4(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(new_n269), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n258), .A2(new_n273), .A3(new_n262), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n276));
  INV_X1    g075(.A(G134gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(new_n277), .A3(G127gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(G127gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT67), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n277), .A2(G127gat), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n278), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G113gat), .ZN(new_n283));
  INV_X1    g082(.A(G120gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G113gat), .A2(G120gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT68), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT1), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n285), .A2(KEYINPUT68), .A3(new_n286), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n282), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n287), .ZN(new_n292));
  INV_X1    g091(.A(new_n281), .ZN(new_n293));
  XNOR2_X1  g092(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n294));
  AND4_X1   g093(.A1(new_n292), .A2(new_n293), .A3(new_n279), .A4(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(G141gat), .B(G148gat), .Z(new_n297));
  NAND2_X1  g096(.A1(G155gat), .A2(G162gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT2), .ZN(new_n299));
  XNOR2_X1  g098(.A(G155gat), .B(G162gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n297), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(KEYINPUT75), .ZN(new_n303));
  INV_X1    g102(.A(G155gat), .ZN(new_n304));
  INV_X1    g103(.A(G162gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT75), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(new_n307), .A3(new_n298), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n299), .A2(KEYINPUT76), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT76), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n298), .A2(new_n312), .A3(KEYINPUT2), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n302), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(KEYINPUT78), .B(KEYINPUT4), .Z(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n296), .A2(new_n315), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n286), .ZN(new_n319));
  NOR2_X1   g118(.A1(G113gat), .A2(G120gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n288), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT1), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n321), .A2(new_n322), .A3(new_n290), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n276), .B1(G127gat), .B2(new_n277), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n293), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n323), .A2(new_n325), .A3(new_n278), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n314), .A2(new_n303), .A3(new_n308), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n292), .A2(new_n293), .A3(new_n279), .A4(new_n294), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n326), .A2(new_n327), .A3(new_n328), .A4(new_n301), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n318), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT5), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n297), .A2(new_n313), .A3(new_n311), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n301), .B1(new_n334), .B2(new_n309), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(KEYINPUT3), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT77), .B1(new_n291), .B2(new_n295), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT77), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n326), .A2(new_n338), .A3(new_n328), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT3), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n340), .B(new_n301), .C1(new_n334), .C2(new_n309), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n336), .A2(new_n337), .A3(new_n339), .A4(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G225gat), .A2(G233gat), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n332), .A2(new_n333), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT79), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n337), .A2(new_n339), .A3(new_n335), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(new_n329), .ZN(new_n347));
  INV_X1    g146(.A(new_n343), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n348), .B1(new_n329), .B2(new_n316), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n296), .A2(KEYINPUT4), .A3(new_n315), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n342), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  AND4_X1   g151(.A1(new_n345), .A2(new_n349), .A3(new_n352), .A4(KEYINPUT5), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n333), .B1(new_n347), .B2(new_n348), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n345), .B1(new_n354), .B2(new_n352), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n344), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  XOR2_X1   g155(.A(G1gat), .B(G29gat), .Z(new_n357));
  XNOR2_X1  g156(.A(G57gat), .B(G85gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT6), .ZN(new_n363));
  INV_X1    g162(.A(new_n361), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n364), .B(new_n344), .C1(new_n353), .C2(new_n355), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n356), .A2(KEYINPUT6), .A3(new_n361), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n264), .A2(new_n269), .A3(new_n271), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(KEYINPUT38), .ZN(new_n369));
  NAND4_X1  g168(.A1(new_n275), .A2(new_n366), .A3(new_n367), .A4(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT3), .B1(new_n212), .B2(new_n255), .ZN(new_n371));
  OR3_X1    g170(.A1(new_n371), .A2(new_n315), .A3(KEYINPUT85), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n212), .B1(new_n341), .B2(new_n255), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT85), .B1(new_n371), .B2(new_n315), .ZN(new_n375));
  INV_X1    g174(.A(G228gat), .ZN(new_n376));
  INV_X1    g175(.A(G233gat), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n372), .A2(new_n374), .A3(new_n375), .A4(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT84), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT83), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n374), .A2(new_n381), .ZN(new_n382));
  AOI211_X1 g181(.A(new_n381), .B(new_n212), .C1(new_n341), .C2(new_n255), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n210), .A2(KEYINPUT82), .A3(new_n211), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT82), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n208), .A2(new_n202), .A3(new_n386), .A4(new_n206), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n387), .A2(new_n255), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT3), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  OR2_X1    g188(.A1(new_n389), .A2(new_n315), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n382), .A2(new_n384), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n378), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n380), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI22_X1  g192(.A1(new_n373), .A2(KEYINPUT83), .B1(new_n389), .B2(new_n315), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n380), .B(new_n392), .C1(new_n394), .C2(new_n383), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n379), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  XOR2_X1   g196(.A(KEYINPUT31), .B(G50gat), .Z(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G78gat), .B(G106gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(G22gat), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n392), .B1(new_n394), .B2(new_n383), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT84), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n395), .ZN(new_n404));
  INV_X1    g203(.A(new_n398), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n405), .A3(new_n379), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n399), .A2(new_n401), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n401), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n405), .B1(new_n404), .B2(new_n379), .ZN(new_n409));
  INV_X1    g208(.A(new_n379), .ZN(new_n410));
  AOI211_X1 g209(.A(new_n398), .B(new_n410), .C1(new_n403), .C2(new_n395), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n408), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n342), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n318), .A2(new_n331), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n348), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n364), .B1(new_n417), .B2(KEYINPUT39), .ZN(new_n418));
  OAI211_X1 g217(.A(KEYINPUT86), .B(KEYINPUT39), .C1(new_n347), .C2(new_n348), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n417), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT39), .B1(new_n347), .B2(new_n348), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT86), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n418), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n425), .A2(KEYINPUT40), .B1(new_n356), .B2(new_n361), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT87), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT30), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n274), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n258), .A2(new_n262), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n269), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n258), .A2(KEYINPUT30), .A3(new_n262), .A4(new_n273), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n343), .B1(new_n332), .B2(new_n342), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT39), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n361), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n424), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n436), .B1(new_n437), .B2(new_n420), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT40), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n426), .A2(new_n427), .A3(new_n433), .A4(new_n440), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n436), .B(KEYINPUT40), .C1(new_n437), .C2(new_n420), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n440), .A2(new_n362), .A3(new_n433), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT87), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n370), .A2(new_n414), .A3(new_n441), .A4(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT36), .ZN(new_n446));
  NAND2_X1  g245(.A1(G227gat), .A2(G233gat), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT34), .B1(new_n448), .B2(KEYINPUT71), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n254), .A2(new_n296), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n326), .A2(new_n328), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n239), .A2(new_n253), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n449), .B1(new_n453), .B2(new_n447), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n239), .A2(new_n253), .A3(new_n451), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n451), .B1(new_n239), .B2(new_n253), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n447), .B(new_n449), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n450), .A2(new_n448), .A3(new_n452), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT32), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT33), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  XOR2_X1   g262(.A(G71gat), .B(G99gat), .Z(new_n464));
  XNOR2_X1  g263(.A(G15gat), .B(G43gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n461), .A2(new_n463), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT70), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n462), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n469), .B1(new_n468), .B2(new_n466), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n460), .A2(KEYINPUT32), .A3(new_n470), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n459), .A2(new_n467), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n454), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n467), .A2(new_n471), .B1(new_n473), .B2(new_n457), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n472), .A2(new_n474), .A3(KEYINPUT72), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n467), .A2(new_n471), .ZN(new_n476));
  INV_X1    g275(.A(new_n459), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT72), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n446), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT36), .B1(new_n472), .B2(new_n474), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n431), .A2(new_n432), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT74), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n431), .A2(KEYINPUT74), .A3(new_n432), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(new_n485), .A3(new_n429), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT81), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(new_n366), .B2(new_n367), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n365), .A2(new_n363), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n349), .A2(new_n352), .A3(KEYINPUT5), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT79), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n354), .A2(new_n345), .A3(new_n352), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n364), .B1(new_n494), .B2(new_n344), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n496), .A2(KEYINPUT81), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n487), .B1(new_n489), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n481), .B1(new_n498), .B2(new_n413), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n472), .A2(new_n474), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n500), .A2(new_n407), .A3(new_n412), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n501), .B(new_n487), .C1(new_n489), .C2(new_n497), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT35), .ZN(new_n503));
  INV_X1    g302(.A(new_n478), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n476), .A2(new_n477), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT72), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n459), .A2(new_n467), .A3(new_n471), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n413), .B1(new_n504), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n367), .B1(new_n490), .B2(new_n495), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n433), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT89), .B(KEYINPUT35), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n509), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n445), .A2(new_n499), .B1(new_n503), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(G229gat), .A2(G233gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(G43gat), .B(G50gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT15), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(KEYINPUT91), .B(G29gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT92), .B(G36gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OR3_X1    g323(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT93), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(new_n519), .B2(KEYINPUT15), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n521), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n519), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT15), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT93), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n522), .A2(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(new_n535), .A3(new_n520), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G15gat), .B(G22gat), .ZN(new_n538));
  INV_X1    g337(.A(G1gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT16), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(G8gat), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n541), .B(new_n542), .C1(G1gat), .C2(new_n538), .ZN(new_n543));
  INV_X1    g342(.A(G15gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(G22gat), .ZN(new_n545));
  INV_X1    g344(.A(G22gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(G15gat), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n540), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(G1gat), .B1(new_n545), .B2(new_n547), .ZN(new_n549));
  OAI21_X1  g348(.A(G8gat), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n537), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n531), .A2(new_n536), .A3(KEYINPUT17), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n543), .A2(new_n550), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(KEYINPUT17), .B1(new_n531), .B2(new_n536), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n518), .B(new_n552), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT18), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  XOR2_X1   g358(.A(new_n518), .B(KEYINPUT13), .Z(new_n560));
  INV_X1    g359(.A(KEYINPUT94), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n554), .A2(new_n561), .A3(new_n531), .A4(new_n536), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(new_n552), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n531), .A2(new_n536), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n561), .B1(new_n564), .B2(new_n554), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n560), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT17), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n537), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(new_n554), .A3(new_n553), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n569), .A2(KEYINPUT18), .A3(new_n518), .A4(new_n552), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n559), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(KEYINPUT90), .ZN(new_n572));
  XNOR2_X1  g371(.A(G113gat), .B(G141gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(G197gat), .ZN(new_n574));
  XOR2_X1   g373(.A(KEYINPUT11), .B(G169gat), .Z(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(KEYINPUT12), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n572), .B(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n517), .A2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(new_n304), .ZN(new_n582));
  XNOR2_X1  g381(.A(G183gat), .B(G211gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n582), .B(new_n583), .Z(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G71gat), .B(G78gat), .Z(new_n586));
  OR2_X1    g385(.A1(G57gat), .A2(G64gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(G57gat), .A2(G64gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT9), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n586), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n587), .A2(KEYINPUT95), .A3(new_n588), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT95), .ZN(new_n593));
  AND2_X1   g392(.A1(G57gat), .A2(G64gat), .ZN(new_n594));
  NOR2_X1   g393(.A1(G57gat), .A2(G64gat), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(G71gat), .B(G78gat), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n592), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g397(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT96), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n591), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT21), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G231gat), .A2(G233gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(G127gat), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n594), .A2(new_n595), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n597), .B1(KEYINPUT9), .B2(new_n609), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n592), .A2(new_n596), .A3(new_n597), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n599), .B(KEYINPUT96), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT21), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n554), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n606), .A2(new_n607), .ZN(new_n616));
  AND3_X1   g415(.A1(new_n608), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n615), .B1(new_n608), .B2(new_n616), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n585), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n608), .A2(new_n616), .ZN(new_n620));
  INV_X1    g419(.A(new_n615), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n608), .A2(new_n615), .A3(new_n616), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n622), .A2(new_n623), .A3(new_n584), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(G232gat), .A2(G233gat), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT41), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(new_n628), .B(KEYINPUT97), .Z(new_n629));
  XNOR2_X1  g428(.A(G134gat), .B(G162gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n626), .A2(new_n627), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(KEYINPUT98), .A2(G85gat), .A3(G92gat), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT7), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(KEYINPUT98), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G99gat), .B(G106gat), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(KEYINPUT99), .ZN(new_n642));
  OR2_X1    g441(.A1(G99gat), .A2(G106gat), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n644));
  NAND2_X1  g443(.A1(G99gat), .A2(G106gat), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(G85gat), .ZN(new_n647));
  INV_X1    g446(.A(G92gat), .ZN(new_n648));
  AOI22_X1  g447(.A1(KEYINPUT8), .A2(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n640), .A2(new_n642), .A3(new_n646), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n638), .A2(new_n639), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n645), .A2(KEYINPUT8), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n647), .A2(new_n648), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g453(.A(KEYINPUT99), .B(new_n641), .C1(new_n651), .C2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n633), .B(new_n635), .C1(new_n564), .C2(new_n657), .ZN(new_n658));
  AOI22_X1  g457(.A1(new_n531), .A2(new_n536), .B1(new_n655), .B2(new_n650), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT100), .B1(new_n659), .B2(new_n634), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(G190gat), .B(G218gat), .Z(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n568), .A2(new_n553), .A3(new_n657), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n661), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n663), .B1(new_n661), .B2(new_n664), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n632), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n667), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n669), .A2(new_n631), .A3(new_n665), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n625), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT101), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n625), .A2(new_n671), .A3(KEYINPUT101), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT103), .ZN(new_n677));
  NAND2_X1  g476(.A1(G230gat), .A2(G233gat), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n613), .A2(new_n656), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n602), .A2(new_n655), .A3(new_n650), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n678), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(G120gat), .B(G148gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(G176gat), .B(G204gat), .ZN(new_n683));
  XOR2_X1   g482(.A(new_n682), .B(new_n683), .Z(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT10), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n679), .A2(new_n686), .A3(new_n680), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT102), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n679), .A2(new_n689), .A3(new_n680), .A4(new_n686), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n613), .A2(new_n656), .A3(KEYINPUT10), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n688), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  AOI211_X1 g491(.A(new_n681), .B(new_n685), .C1(new_n692), .C2(new_n678), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n687), .A2(KEYINPUT102), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n690), .A2(new_n691), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n678), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n681), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n684), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n677), .B1(new_n693), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n678), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n690), .A2(new_n691), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n700), .B1(new_n701), .B2(new_n688), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n685), .B1(new_n702), .B2(new_n681), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n696), .A2(new_n697), .A3(new_n684), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(KEYINPUT103), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n676), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n580), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n489), .A2(new_n497), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(new_n539), .ZN(G1324gat));
  AND2_X1   g511(.A1(new_n580), .A2(new_n707), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n542), .B1(new_n713), .B2(new_n433), .ZN(new_n714));
  XNOR2_X1  g513(.A(KEYINPUT16), .B(G8gat), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n708), .A2(new_n512), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(KEYINPUT42), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(KEYINPUT42), .B2(new_n716), .ZN(G1325gat));
  NAND2_X1  g517(.A1(new_n504), .A2(new_n508), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n713), .A2(new_n544), .A3(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n480), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n721), .B1(new_n719), .B2(new_n446), .ZN(new_n722));
  OAI21_X1  g521(.A(G15gat), .B1(new_n708), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n720), .A2(new_n723), .ZN(G1326gat));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n713), .A2(new_n725), .A3(new_n413), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT104), .B1(new_n708), .B2(new_n414), .ZN(new_n727));
  XNOR2_X1  g526(.A(KEYINPUT43), .B(G22gat), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n726), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n728), .B1(new_n726), .B2(new_n727), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(G1327gat));
  NAND2_X1  g530(.A1(new_n510), .A2(KEYINPUT81), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n366), .A2(new_n488), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n486), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n445), .B(new_n722), .C1(new_n414), .C2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT35), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n736), .B1(new_n734), .B2(new_n501), .ZN(new_n737));
  INV_X1    g536(.A(new_n516), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n735), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n578), .ZN(new_n740));
  INV_X1    g539(.A(new_n706), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(new_n625), .ZN(new_n742));
  INV_X1    g541(.A(new_n671), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XOR2_X1   g543(.A(new_n744), .B(KEYINPUT105), .Z(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n740), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n710), .A2(new_n522), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT45), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n742), .A2(new_n578), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT106), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(KEYINPUT44), .B1(new_n517), .B2(new_n671), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n671), .B(KEYINPUT107), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n739), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n753), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n709), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n522), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n750), .A2(new_n760), .ZN(G1328gat));
  NOR2_X1   g560(.A1(new_n512), .A2(new_n523), .ZN(new_n762));
  AND2_X1   g561(.A1(new_n747), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT46), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n758), .A2(new_n433), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n523), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(G1329gat));
  INV_X1    g566(.A(KEYINPUT108), .ZN(new_n768));
  XNOR2_X1  g567(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n769));
  INV_X1    g568(.A(G43gat), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n758), .B2(new_n481), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n719), .A2(new_n770), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n740), .A2(new_n746), .A3(new_n772), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n768), .B(new_n769), .C1(new_n771), .C2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n769), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n755), .B1(new_n739), .B2(new_n743), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n756), .A2(new_n755), .ZN(new_n777));
  AOI22_X1  g576(.A1(new_n502), .A2(KEYINPUT35), .B1(new_n509), .B2(new_n515), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n777), .B1(new_n779), .B2(new_n735), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n481), .B(new_n752), .C1(new_n776), .C2(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n773), .B1(new_n781), .B2(G43gat), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n775), .B1(new_n782), .B2(KEYINPUT108), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n774), .A2(new_n783), .ZN(G1330gat));
  NAND2_X1  g583(.A1(new_n754), .A2(new_n757), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n785), .A2(G50gat), .A3(new_n413), .A4(new_n752), .ZN(new_n786));
  OR2_X1    g585(.A1(KEYINPUT110), .A2(KEYINPUT48), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n739), .A2(new_n745), .A3(new_n413), .A4(new_n578), .ZN(new_n788));
  INV_X1    g587(.A(G50gat), .ZN(new_n789));
  AOI22_X1  g588(.A1(new_n788), .A2(new_n789), .B1(KEYINPUT110), .B2(KEYINPUT48), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n786), .A2(new_n787), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n787), .B1(new_n786), .B2(new_n790), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(G1331gat));
  NAND2_X1  g592(.A1(new_n676), .A2(new_n579), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(new_n706), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n739), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n709), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT112), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n797), .B(new_n798), .ZN(new_n799));
  XNOR2_X1  g598(.A(KEYINPUT111), .B(G57gat), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n797), .B(KEYINPUT112), .ZN(new_n802));
  INV_X1    g601(.A(new_n800), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(G1332gat));
  NAND2_X1  g604(.A1(new_n739), .A2(new_n795), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(new_n512), .ZN(new_n807));
  NOR2_X1   g606(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n808));
  AND2_X1   g607(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n810), .B1(new_n807), .B2(new_n808), .ZN(G1333gat));
  INV_X1    g610(.A(G71gat), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n796), .A2(new_n812), .A3(new_n719), .ZN(new_n813));
  OAI21_X1  g612(.A(G71gat), .B1(new_n806), .B2(new_n722), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XOR2_X1   g614(.A(new_n815), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g615(.A1(new_n806), .A2(new_n414), .ZN(new_n817));
  XNOR2_X1  g616(.A(KEYINPUT113), .B(G78gat), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n817), .B(new_n818), .ZN(G1335gat));
  NOR3_X1   g618(.A1(new_n578), .A2(new_n706), .A3(new_n625), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n785), .A2(new_n709), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n578), .A2(new_n625), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n722), .B1(new_n734), .B2(new_n414), .ZN(new_n823));
  INV_X1    g622(.A(new_n445), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n743), .B(new_n822), .C1(new_n825), .C2(new_n778), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT51), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n739), .A2(KEYINPUT51), .A3(new_n743), .A4(new_n822), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n709), .A2(new_n647), .A3(new_n741), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT114), .ZN(new_n833));
  OAI22_X1  g632(.A1(new_n821), .A2(new_n647), .B1(new_n831), .B2(new_n833), .ZN(G1336gat));
  OAI211_X1 g633(.A(new_n433), .B(new_n820), .C1(new_n776), .C2(new_n780), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(G92gat), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n741), .A2(new_n648), .A3(new_n433), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT115), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n836), .B(new_n837), .C1(new_n831), .C2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n826), .A2(new_n841), .A3(KEYINPUT51), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT51), .B1(new_n826), .B2(new_n841), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n839), .ZN(new_n845));
  AOI22_X1  g644(.A1(new_n844), .A2(new_n845), .B1(G92gat), .B2(new_n835), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n840), .B1(new_n846), .B2(new_n837), .ZN(G1337gat));
  AND3_X1   g646(.A1(new_n785), .A2(new_n481), .A3(new_n820), .ZN(new_n848));
  INV_X1    g647(.A(G99gat), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n719), .A2(new_n849), .A3(new_n741), .ZN(new_n850));
  OAI22_X1  g649(.A1(new_n848), .A2(new_n849), .B1(new_n831), .B2(new_n850), .ZN(G1338gat));
  OAI211_X1 g650(.A(new_n413), .B(new_n820), .C1(new_n776), .C2(new_n780), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n852), .A2(G106gat), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n414), .A2(G106gat), .A3(new_n706), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n842), .A2(new_n843), .A3(new_n855), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT53), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT53), .B1(new_n852), .B2(G106gat), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n859), .B1(new_n830), .B2(new_n854), .ZN(new_n860));
  AOI211_X1 g659(.A(KEYINPUT117), .B(new_n855), .C1(new_n828), .C2(new_n829), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n858), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n857), .A2(new_n862), .ZN(G1339gat));
  INV_X1    g662(.A(new_n625), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n559), .A2(new_n570), .A3(new_n566), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n562), .A2(new_n552), .ZN(new_n866));
  INV_X1    g665(.A(new_n560), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT94), .B1(new_n537), .B2(new_n551), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n866), .A2(KEYINPUT119), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n552), .B1(new_n555), .B2(new_n556), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n870), .A2(G229gat), .A3(G233gat), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n868), .A2(new_n552), .A3(new_n867), .A4(new_n562), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n869), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  AOI22_X1  g674(.A1(new_n865), .A2(new_n577), .B1(new_n875), .B2(new_n576), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n699), .A2(new_n705), .A3(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT120), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n699), .A2(new_n705), .A3(new_n876), .A4(KEYINPUT120), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT55), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n688), .A2(new_n700), .A3(new_n690), .A4(new_n691), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n696), .A2(KEYINPUT54), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n685), .B1(new_n696), .B2(KEYINPUT54), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n882), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n684), .B1(new_n702), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n696), .A2(KEYINPUT54), .A3(new_n883), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(KEYINPUT55), .A3(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n886), .A2(new_n704), .A3(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT118), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n886), .A2(KEYINPUT118), .A3(new_n890), .A4(new_n704), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n893), .A2(new_n578), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n756), .B1(new_n881), .B2(new_n895), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n756), .A2(new_n893), .A3(new_n894), .A4(new_n876), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n864), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n674), .A2(new_n579), .A3(new_n706), .A4(new_n675), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n710), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n901), .A2(KEYINPUT122), .A3(new_n501), .ZN(new_n902));
  AOI21_X1  g701(.A(KEYINPUT122), .B1(new_n901), .B2(new_n501), .ZN(new_n903));
  OR2_X1    g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n904), .A2(new_n283), .A3(new_n512), .A4(new_n578), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n901), .A2(new_n512), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n907), .A2(new_n509), .A3(new_n578), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n906), .B1(new_n908), .B2(G113gat), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n908), .A2(new_n906), .A3(G113gat), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n905), .B1(new_n909), .B2(new_n910), .ZN(G1340gat));
  NAND2_X1  g710(.A1(new_n907), .A2(new_n509), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n912), .A2(new_n284), .A3(new_n706), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n904), .A2(new_n512), .A3(new_n741), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n913), .B1(new_n914), .B2(new_n284), .ZN(G1341gat));
  NAND4_X1  g714(.A1(new_n904), .A2(new_n607), .A3(new_n512), .A4(new_n625), .ZN(new_n916));
  OAI21_X1  g715(.A(G127gat), .B1(new_n912), .B2(new_n864), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1342gat));
  NOR2_X1   g717(.A1(new_n671), .A2(G134gat), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n512), .B(new_n919), .C1(new_n902), .C2(new_n903), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n920), .A2(KEYINPUT56), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(KEYINPUT56), .ZN(new_n922));
  OAI21_X1  g721(.A(G134gat), .B1(new_n912), .B2(new_n671), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(G1343gat));
  NOR2_X1   g723(.A1(new_n481), .A2(new_n414), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT123), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n901), .A2(new_n926), .A3(new_n512), .A4(new_n578), .ZN(new_n927));
  INV_X1    g726(.A(G141gat), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n414), .B1(new_n899), .B2(new_n900), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT57), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n709), .A2(new_n722), .A3(new_n512), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n877), .B1(new_n579), .B2(new_n891), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n671), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n625), .B1(new_n935), .B2(new_n897), .ZN(new_n936));
  INV_X1    g735(.A(new_n900), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n413), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n933), .B1(new_n938), .B2(KEYINPUT57), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n932), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n578), .A2(G141gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n929), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT58), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n942), .B(new_n943), .ZN(G1344gat));
  NOR2_X1   g743(.A1(new_n940), .A2(new_n706), .ZN(new_n945));
  INV_X1    g744(.A(G148gat), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n945), .A2(KEYINPUT59), .A3(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT59), .ZN(new_n948));
  INV_X1    g747(.A(new_n930), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT57), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n900), .B(KEYINPUT124), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n743), .A2(new_n876), .ZN(new_n952));
  OR2_X1    g751(.A1(new_n952), .A2(new_n891), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n625), .B1(new_n935), .B2(new_n953), .ZN(new_n954));
  OAI211_X1 g753(.A(new_n931), .B(new_n413), .C1(new_n951), .C2(new_n954), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n933), .A2(new_n706), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n950), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n948), .B1(new_n957), .B2(G148gat), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n907), .A2(new_n926), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n741), .A2(new_n946), .ZN(new_n960));
  OAI22_X1  g759(.A1(new_n947), .A2(new_n958), .B1(new_n959), .B2(new_n960), .ZN(G1345gat));
  OAI21_X1  g760(.A(G155gat), .B1(new_n940), .B2(new_n864), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n625), .A2(new_n304), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n962), .B1(new_n959), .B2(new_n963), .ZN(G1346gat));
  INV_X1    g763(.A(new_n756), .ZN(new_n965));
  OAI21_X1  g764(.A(KEYINPUT125), .B1(new_n940), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G162gat), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n940), .A2(KEYINPUT125), .A3(new_n965), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n743), .A2(new_n305), .ZN(new_n969));
  OAI22_X1  g768(.A1(new_n967), .A2(new_n968), .B1(new_n959), .B2(new_n969), .ZN(G1347gat));
  NAND2_X1  g769(.A1(new_n899), .A2(new_n900), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n709), .A2(new_n512), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(new_n501), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g774(.A(G169gat), .B1(new_n975), .B2(new_n578), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n971), .A2(new_n509), .A3(new_n972), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n578), .A2(G169gat), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(G1348gat));
  INV_X1    g778(.A(G176gat), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n975), .A2(new_n980), .A3(new_n741), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n977), .A2(new_n741), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n981), .B1(new_n982), .B2(new_n980), .ZN(G1349gat));
  NAND2_X1  g782(.A1(new_n977), .A2(new_n625), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(G183gat), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n975), .A2(new_n240), .A3(new_n625), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g786(.A(new_n987), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g787(.A1(new_n975), .A2(new_n218), .A3(new_n756), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT61), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n977), .A2(new_n743), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n990), .B1(new_n991), .B2(G190gat), .ZN(new_n992));
  AOI211_X1 g791(.A(KEYINPUT61), .B(new_n218), .C1(new_n977), .C2(new_n743), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n989), .B1(new_n992), .B2(new_n993), .ZN(G1351gat));
  NAND2_X1  g793(.A1(new_n972), .A2(new_n722), .ZN(new_n995));
  XNOR2_X1  g794(.A(new_n995), .B(KEYINPUT126), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n950), .A2(new_n955), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n578), .A2(G197gat), .ZN(new_n998));
  NOR3_X1   g797(.A1(new_n949), .A2(new_n579), .A3(new_n995), .ZN(new_n999));
  OAI22_X1  g798(.A1(new_n997), .A2(new_n998), .B1(G197gat), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g799(.A(new_n1000), .ZN(G1352gat));
  NOR2_X1   g800(.A1(new_n949), .A2(new_n995), .ZN(new_n1002));
  INV_X1    g801(.A(G204gat), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n1002), .A2(new_n1003), .A3(new_n741), .ZN(new_n1004));
  OR2_X1    g803(.A1(new_n1004), .A2(KEYINPUT62), .ZN(new_n1005));
  OAI21_X1  g804(.A(G204gat), .B1(new_n997), .B2(new_n706), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1004), .A2(KEYINPUT62), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(G1353gat));
  INV_X1    g807(.A(KEYINPUT63), .ZN(new_n1009));
  NOR2_X1   g808(.A1(new_n995), .A2(new_n864), .ZN(new_n1010));
  OAI211_X1 g809(.A(new_n955), .B(new_n1010), .C1(new_n930), .C2(new_n931), .ZN(new_n1011));
  AND2_X1   g810(.A1(new_n1011), .A2(KEYINPUT127), .ZN(new_n1012));
  OAI21_X1  g811(.A(G211gat), .B1(new_n1011), .B2(KEYINPUT127), .ZN(new_n1013));
  OAI21_X1  g812(.A(new_n1009), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g813(.A(KEYINPUT127), .ZN(new_n1015));
  NAND4_X1  g814(.A1(new_n950), .A2(new_n1015), .A3(new_n955), .A4(new_n1010), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1011), .A2(KEYINPUT127), .ZN(new_n1017));
  NAND4_X1  g816(.A1(new_n1016), .A2(new_n1017), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g818(.A1(new_n930), .A2(new_n204), .A3(new_n1010), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1019), .A2(new_n1020), .ZN(G1354gat));
  OAI21_X1  g820(.A(G218gat), .B1(new_n997), .B2(new_n671), .ZN(new_n1022));
  NAND3_X1  g821(.A1(new_n1002), .A2(new_n205), .A3(new_n756), .ZN(new_n1023));
  NAND2_X1  g822(.A1(new_n1022), .A2(new_n1023), .ZN(G1355gat));
endmodule


