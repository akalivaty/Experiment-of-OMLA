//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1120, new_n1121, new_n1122;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g019(.A(KEYINPUT66), .B(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT67), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT68), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT69), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n465), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n473), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(new_n462), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n472), .A2(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n470), .A2(G136), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n469), .A2(new_n462), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NOR2_X1   g054(.A1(G100), .A2(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(G2104), .B1(new_n462), .B2(G112), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n477), .B(new_n479), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G162));
  OAI21_X1  g058(.A(G2104), .B1(new_n462), .B2(G114), .ZN(new_n484));
  NOR2_X1   g059(.A1(G102), .A2(G2105), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AND2_X1   g061(.A1(G126), .A2(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n487), .B1(new_n467), .B2(new_n468), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT70), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(new_n487), .C1(new_n467), .C2(new_n468), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n486), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n462), .C1(new_n467), .C2(new_n468), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT72), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n493), .B(new_n494), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT4), .B1(new_n495), .B2(new_n493), .ZN(new_n500));
  OAI211_X1 g075(.A(new_n492), .B(new_n497), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT5), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G62), .ZN(new_n510));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  XOR2_X1   g086(.A(new_n511), .B(KEYINPUT73), .Z(new_n512));
  AOI21_X1  g087(.A(new_n503), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(G50), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G88), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n514), .B1(new_n508), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n513), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n521), .B(new_n522), .ZN(G166));
  NAND2_X1  g098(.A1(new_n520), .A2(KEYINPUT75), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n517), .A2(new_n519), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT75), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n524), .A2(G543), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n520), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n530), .A2(new_n508), .ZN(new_n531));
  NAND3_X1  g106(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n532), .B(KEYINPUT7), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n529), .A2(new_n531), .A3(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  NOR2_X1   g110(.A1(new_n508), .A2(new_n525), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G90), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n524), .A2(G543), .A3(new_n527), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  OAI221_X1 g115(.A(new_n537), .B1(new_n538), .B2(new_n503), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT76), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(new_n528), .A2(G43), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n503), .ZN(new_n546));
  XNOR2_X1  g121(.A(KEYINPUT77), .B(G81), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n536), .A2(new_n547), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(new_n528), .A2(G53), .ZN(new_n556));
  NAND2_X1  g131(.A1(KEYINPUT78), .A2(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n508), .B2(new_n559), .ZN(new_n560));
  AOI22_X1  g135(.A1(new_n556), .A2(new_n557), .B1(G651), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n536), .A2(G91), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n561), .B(new_n562), .C1(new_n556), .C2(new_n557), .ZN(G299));
  XNOR2_X1  g138(.A(new_n521), .B(KEYINPUT74), .ZN(G303));
  OAI21_X1  g139(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n565));
  INV_X1    g140(.A(new_n536), .ZN(new_n566));
  INV_X1    g141(.A(G87), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n568), .B1(G49), .B2(new_n528), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G288));
  INV_X1    g145(.A(G48), .ZN(new_n571));
  NOR3_X1   g146(.A1(new_n525), .A2(new_n571), .A3(new_n504), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G61), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n508), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n572), .B1(G651), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n536), .A2(G86), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(G305));
  AOI22_X1  g153(.A1(new_n528), .A2(G47), .B1(G85), .B2(new_n536), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n580), .B(KEYINPUT79), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n579), .B1(new_n581), .B2(new_n503), .ZN(G290));
  NAND2_X1  g157(.A1(G301), .A2(G868), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n536), .A2(G92), .ZN(new_n584));
  XOR2_X1   g159(.A(new_n584), .B(KEYINPUT10), .Z(new_n585));
  AND2_X1   g160(.A1(new_n509), .A2(G66), .ZN(new_n586));
  NAND2_X1  g161(.A1(G79), .A2(G543), .ZN(new_n587));
  XOR2_X1   g162(.A(new_n587), .B(KEYINPUT80), .Z(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n528), .A2(G54), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n585), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  XOR2_X1   g166(.A(new_n591), .B(KEYINPUT81), .Z(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n583), .B1(new_n593), .B2(G868), .ZN(G284));
  OAI21_X1  g169(.A(new_n583), .B1(new_n593), .B2(G868), .ZN(G321));
  INV_X1    g170(.A(G868), .ZN(new_n596));
  NAND2_X1  g171(.A1(G299), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n597), .B1(new_n596), .B2(G168), .ZN(G297));
  OAI21_X1  g173(.A(new_n597), .B1(new_n596), .B2(G168), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n593), .B1(new_n600), .B2(G860), .ZN(G148));
  INV_X1    g176(.A(new_n549), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(new_n596), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n592), .A2(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(new_n596), .ZN(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g181(.A1(new_n464), .A2(new_n473), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT12), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT13), .ZN(new_n609));
  INV_X1    g184(.A(G2100), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n470), .A2(G135), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n478), .A2(G123), .ZN(new_n613));
  NOR2_X1   g188(.A1(G99), .A2(G2105), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n615));
  OAI211_X1 g190(.A(new_n612), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(G2096), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n611), .A2(new_n618), .ZN(G156));
  XNOR2_X1  g194(.A(KEYINPUT15), .B(G2435), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT82), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2438), .ZN(new_n622));
  XNOR2_X1  g197(.A(G2427), .B(G2430), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(KEYINPUT14), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2443), .ZN(new_n626));
  XNOR2_X1  g201(.A(G1341), .B(G1348), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2446), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT16), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n626), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G2451), .B(G2454), .Z(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT83), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n630), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n633), .A2(G14), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT84), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(G401));
  XOR2_X1   g212(.A(G2084), .B(G2090), .Z(new_n638));
  XNOR2_X1  g213(.A(G2072), .B(G2078), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT17), .ZN(new_n640));
  XOR2_X1   g215(.A(G2067), .B(G2678), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n638), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n639), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT86), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n642), .A2(new_n638), .A3(new_n639), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT85), .B(KEYINPUT18), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n640), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n649), .A2(new_n638), .A3(new_n641), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n645), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(new_n617), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(new_n610), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G227));
  XNOR2_X1  g229(.A(G1971), .B(G1976), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT19), .ZN(new_n656));
  XOR2_X1   g231(.A(G1956), .B(G2474), .Z(new_n657));
  XOR2_X1   g232(.A(G1961), .B(G1966), .Z(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n656), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n657), .A2(new_n658), .ZN(new_n662));
  AOI22_X1  g237(.A1(new_n660), .A2(KEYINPUT20), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  INV_X1    g238(.A(new_n662), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n664), .A2(new_n656), .A3(new_n659), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n663), .B(new_n665), .C1(KEYINPUT20), .C2(new_n660), .ZN(new_n666));
  XOR2_X1   g241(.A(G1991), .B(G1996), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G229));
  INV_X1    g247(.A(G29), .ZN(new_n673));
  AND2_X1   g248(.A1(new_n673), .A2(G25), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n478), .A2(G119), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT87), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(G131), .B2(new_n470), .ZN(new_n677));
  OR2_X1    g252(.A1(G95), .A2(G2105), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n678), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n674), .B1(new_n680), .B2(G29), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT88), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT35), .B(G1991), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  AND2_X1   g261(.A1(new_n686), .A2(G24), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(G290), .B2(G16), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G1986), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(G16), .A2(G22), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(G166), .B2(G16), .ZN(new_n693));
  INV_X1    g268(.A(G1971), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  MUX2_X1   g270(.A(G6), .B(G305), .S(G16), .Z(new_n696));
  XOR2_X1   g271(.A(KEYINPUT32), .B(G1981), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n686), .A2(G23), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(new_n569), .B2(new_n686), .ZN(new_n700));
  XNOR2_X1  g275(.A(KEYINPUT89), .B(KEYINPUT33), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(G1976), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n700), .B(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n695), .A2(new_n698), .A3(new_n703), .ZN(new_n704));
  AOI211_X1 g279(.A(new_n684), .B(new_n691), .C1(KEYINPUT34), .C2(new_n704), .ZN(new_n705));
  OAI221_X1 g280(.A(new_n705), .B1(KEYINPUT34), .B2(new_n704), .C1(G1986), .C2(new_n689), .ZN(new_n706));
  AND2_X1   g281(.A1(KEYINPUT90), .A2(KEYINPUT36), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G27), .ZN(new_n709));
  OAI21_X1  g284(.A(KEYINPUT98), .B1(new_n709), .B2(G29), .ZN(new_n710));
  OR3_X1    g285(.A1(new_n709), .A2(KEYINPUT98), .A3(G29), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n710), .B(new_n711), .C1(G164), .C2(new_n673), .ZN(new_n712));
  INV_X1    g287(.A(G2078), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NOR2_X1   g289(.A1(G4), .A2(G16), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n593), .B2(G16), .ZN(new_n716));
  INV_X1    g291(.A(G1348), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n470), .A2(G140), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n478), .A2(G128), .ZN(new_n720));
  NOR2_X1   g295(.A1(G104), .A2(G2105), .ZN(new_n721));
  OAI21_X1  g296(.A(G2104), .B1(new_n462), .B2(G116), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n719), .B(new_n720), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n673), .A2(G26), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT92), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT28), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(G2067), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n686), .A2(G19), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(new_n549), .B2(new_n686), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT91), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1341), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n718), .A2(new_n730), .A3(new_n734), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT93), .Z(new_n736));
  INV_X1    g311(.A(KEYINPUT100), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n673), .A2(G35), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G162), .B2(new_n673), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT99), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT29), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(G2090), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(G2090), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n737), .A2(new_n742), .B1(new_n743), .B2(KEYINPUT101), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(KEYINPUT101), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT25), .Z(new_n747));
  NAND2_X1  g322(.A1(new_n470), .A2(G139), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n747), .B(new_n748), .C1(new_n462), .C2(new_n749), .ZN(new_n750));
  MUX2_X1   g325(.A(G33), .B(new_n750), .S(G29), .Z(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(G2072), .Z(new_n752));
  XOR2_X1   g327(.A(KEYINPUT96), .B(KEYINPUT30), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G28), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(new_n673), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT31), .B(G11), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n755), .B(new_n756), .C1(new_n616), .C2(new_n673), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT97), .ZN(new_n758));
  NOR2_X1   g333(.A1(G168), .A2(new_n686), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n686), .B2(G21), .ZN(new_n760));
  INV_X1    g335(.A(G1966), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n744), .A2(new_n745), .A3(new_n752), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(G299), .A2(G16), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(KEYINPUT23), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n686), .A2(G20), .ZN(new_n766));
  MUX2_X1   g341(.A(KEYINPUT23), .B(new_n765), .S(new_n766), .Z(new_n767));
  OR2_X1    g342(.A1(new_n767), .A2(G1956), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(G1956), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n768), .B(new_n769), .C1(new_n737), .C2(new_n742), .ZN(new_n770));
  OR2_X1    g345(.A1(KEYINPUT24), .A2(G34), .ZN(new_n771));
  NAND2_X1  g346(.A1(KEYINPUT24), .A2(G34), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n771), .A2(new_n673), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G160), .B2(new_n673), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n774), .A2(G2084), .ZN(new_n775));
  OAI22_X1  g350(.A1(new_n760), .A2(new_n761), .B1(G2084), .B2(new_n774), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n673), .A2(G32), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n464), .A2(G105), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n470), .A2(G141), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n478), .A2(G129), .ZN(new_n780));
  NAND3_X1  g355(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT26), .Z(new_n782));
  NAND4_X1  g357(.A1(new_n778), .A2(new_n779), .A3(new_n780), .A4(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT94), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n777), .B1(new_n784), .B2(G29), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT27), .B(G1996), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT95), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n776), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(G5), .A2(G16), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G171), .B2(G16), .ZN(new_n790));
  INV_X1    g365(.A(G1961), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n788), .B(new_n792), .C1(new_n787), .C2(new_n785), .ZN(new_n793));
  NOR4_X1   g368(.A1(new_n763), .A2(new_n770), .A3(new_n775), .A4(new_n793), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n708), .A2(new_n714), .A3(new_n736), .A4(new_n794), .ZN(G150));
  INV_X1    g370(.A(G150), .ZN(G311));
  NAND2_X1  g371(.A1(new_n536), .A2(G93), .ZN(new_n797));
  INV_X1    g372(.A(G55), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n539), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n799), .A2(KEYINPUT102), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n799), .A2(KEYINPUT102), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n802));
  OAI22_X1  g377(.A1(new_n800), .A2(new_n801), .B1(new_n503), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n803), .A2(G860), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT37), .Z(new_n805));
  NOR2_X1   g380(.A1(new_n592), .A2(new_n600), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT103), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n803), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n549), .B1(new_n803), .B2(new_n809), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n808), .B(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n805), .B1(new_n813), .B2(G860), .ZN(G145));
  NAND2_X1  g389(.A1(new_n470), .A2(G142), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n478), .A2(G130), .ZN(new_n816));
  NOR2_X1   g391(.A1(G106), .A2(G2105), .ZN(new_n817));
  OAI21_X1  g392(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n815), .B(new_n816), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n680), .B(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT105), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n821), .A2(new_n608), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT105), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n820), .B(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(new_n608), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n828));
  INV_X1    g403(.A(new_n486), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n490), .B1(new_n473), .B2(new_n487), .ZN(new_n830));
  INV_X1    g405(.A(new_n491), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(KEYINPUT104), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT104), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n492), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n828), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(new_n723), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n783), .A2(new_n750), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(new_n784), .B2(new_n750), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n837), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n827), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n822), .A2(new_n826), .A3(new_n840), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n842), .A2(KEYINPUT106), .A3(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(G160), .B(new_n616), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(G162), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n844), .B(new_n846), .C1(KEYINPUT106), .C2(new_n843), .ZN(new_n847));
  INV_X1    g422(.A(G37), .ZN(new_n848));
  INV_X1    g423(.A(new_n846), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n842), .A2(new_n843), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n847), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g427(.A(new_n812), .B(KEYINPUT107), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(G559), .B2(new_n592), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n812), .A2(KEYINPUT107), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n812), .A2(KEYINPUT107), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n855), .A2(new_n604), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n591), .ZN(new_n859));
  XNOR2_X1  g434(.A(G299), .B(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(G290), .B(G305), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(G166), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n569), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT108), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n864), .B1(new_n865), .B2(KEYINPUT42), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n860), .B(KEYINPUT41), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n861), .B(new_n867), .C1(new_n868), .C2(new_n858), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n865), .A2(KEYINPUT42), .ZN(new_n870));
  INV_X1    g445(.A(new_n868), .ZN(new_n871));
  AND3_X1   g446(.A1(new_n854), .A2(new_n871), .A3(new_n857), .ZN(new_n872));
  INV_X1    g447(.A(new_n860), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(new_n854), .B2(new_n857), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n866), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  AND3_X1   g450(.A1(new_n869), .A2(new_n870), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n870), .B1(new_n869), .B2(new_n875), .ZN(new_n877));
  OAI21_X1  g452(.A(G868), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n803), .A2(new_n596), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(G295));
  NAND2_X1  g455(.A1(new_n878), .A2(new_n879), .ZN(G331));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n882));
  XNOR2_X1  g457(.A(G301), .B(G168), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n812), .B(new_n883), .Z(new_n884));
  NAND2_X1  g459(.A1(new_n884), .A2(new_n871), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n812), .B(new_n883), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n860), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n885), .A2(new_n864), .A3(new_n887), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n888), .A2(new_n848), .ZN(new_n889));
  XOR2_X1   g464(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n885), .A2(new_n887), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n889), .B(new_n891), .C1(new_n864), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n888), .A2(new_n848), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n868), .A2(KEYINPUT110), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n860), .A2(new_n896), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n884), .B(new_n895), .C1(KEYINPUT110), .C2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n864), .B1(new_n898), .B2(new_n887), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT43), .B1(new_n894), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n882), .B1(new_n893), .B2(new_n900), .ZN(new_n901));
  OR3_X1    g476(.A1(new_n894), .A2(new_n899), .A3(new_n890), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n892), .A2(new_n864), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n890), .B1(new_n903), .B2(new_n894), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n901), .B1(new_n905), .B2(new_n882), .ZN(G397));
  INV_X1    g481(.A(KEYINPUT45), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n907), .B1(new_n836), .B2(G1384), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  OAI211_X1 g484(.A(new_n465), .B(G40), .C1(new_n466), .C2(new_n471), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n910), .A2(new_n475), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT46), .ZN(new_n913));
  OR3_X1    g488(.A1(new_n912), .A2(new_n913), .A3(G1996), .ZN(new_n914));
  INV_X1    g489(.A(new_n912), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n723), .B(new_n729), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n915), .B1(new_n783), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n913), .B1(new_n912), .B2(G1996), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n914), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT47), .ZN(new_n921));
  NOR3_X1   g496(.A1(new_n912), .A2(G1986), .A3(G290), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n922), .B(KEYINPUT48), .Z(new_n923));
  OAI21_X1  g498(.A(new_n916), .B1(new_n784), .B2(G1996), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n924), .B1(G1996), .B2(new_n783), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(new_n683), .B2(new_n680), .ZN(new_n926));
  INV_X1    g501(.A(new_n680), .ZN(new_n927));
  INV_X1    g502(.A(new_n683), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n915), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n923), .A2(new_n930), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n925), .A2(new_n928), .A3(new_n927), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n723), .A2(G2067), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n915), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n921), .A2(new_n931), .A3(new_n934), .ZN(new_n935));
  XOR2_X1   g510(.A(new_n935), .B(KEYINPUT127), .Z(new_n936));
  INV_X1    g511(.A(KEYINPUT112), .ZN(new_n937));
  OR3_X1    g512(.A1(G305), .A2(new_n937), .A3(G1981), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n937), .B1(G305), .B2(G1981), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g515(.A(KEYINPUT113), .B(G86), .Z(new_n941));
  OAI21_X1  g516(.A(new_n576), .B1(new_n566), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(G1981), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT49), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n833), .A2(new_n835), .ZN(new_n947));
  INV_X1    g522(.A(new_n497), .ZN(new_n948));
  INV_X1    g523(.A(new_n500), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n948), .B1(new_n949), .B2(new_n498), .ZN(new_n950));
  AOI21_X1  g525(.A(G1384), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n911), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(G8), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n940), .A2(KEYINPUT49), .A3(new_n943), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n946), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(G1976), .ZN(new_n957));
  AND2_X1   g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n958), .A2(new_n569), .B1(new_n939), .B2(new_n938), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT55), .ZN(new_n960));
  INV_X1    g535(.A(G8), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n960), .B1(G166), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n965));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n492), .A2(new_n834), .ZN(new_n967));
  AOI211_X1 g542(.A(KEYINPUT104), .B(new_n486), .C1(new_n489), .C2(new_n491), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n965), .B(new_n966), .C1(new_n969), .C2(new_n828), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n501), .A2(new_n966), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT50), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n970), .A2(new_n911), .A3(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n973), .A2(G2090), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT45), .B1(new_n501), .B2(new_n966), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(new_n951), .B2(KEYINPUT45), .ZN(new_n976));
  AOI21_X1  g551(.A(G1971), .B1(new_n976), .B2(new_n911), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n964), .B(G8), .C1(new_n974), .C2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT52), .B1(G288), .B2(new_n957), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n954), .B(new_n979), .C1(new_n957), .C2(G288), .ZN(new_n980));
  NOR2_X1   g555(.A1(G288), .A2(new_n957), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT52), .B1(new_n953), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n980), .A2(new_n956), .A3(new_n982), .ZN(new_n983));
  OAI22_X1  g558(.A1(new_n959), .A2(new_n953), .B1(new_n978), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n951), .A2(KEYINPUT45), .ZN(new_n985));
  INV_X1    g560(.A(new_n975), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n985), .A2(new_n713), .A3(new_n911), .A4(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n988));
  AOI22_X1  g563(.A1(new_n987), .A2(new_n988), .B1(new_n791), .B2(new_n973), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n966), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n988), .A2(G2078), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n908), .A2(new_n911), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(G171), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n970), .A2(new_n911), .A3(new_n972), .ZN(new_n995));
  INV_X1    g570(.A(G2084), .ZN(new_n996));
  OAI211_X1 g571(.A(new_n911), .B(new_n990), .C1(new_n951), .C2(KEYINPUT45), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n995), .A2(new_n996), .B1(new_n997), .B2(new_n761), .ZN(new_n998));
  NAND2_X1  g573(.A1(G286), .A2(G8), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n1001), .B(new_n999), .C1(new_n998), .C2(new_n961), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n997), .A2(new_n761), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n970), .A2(new_n996), .A3(new_n911), .A4(new_n972), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g580(.A(KEYINPUT51), .B(G8), .C1(new_n1005), .C2(G286), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1000), .B1(new_n1002), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n1007), .B(KEYINPUT122), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n994), .B1(new_n1008), .B2(KEYINPUT62), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n501), .A2(new_n965), .A3(new_n966), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n911), .B(new_n1010), .C1(new_n951), .C2(new_n965), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G2090), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT50), .B1(new_n836), .B2(G1384), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n1015), .A2(KEYINPUT114), .A3(new_n911), .A4(new_n1010), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n977), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n964), .B1(new_n1019), .B2(G8), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n983), .B1(new_n1020), .B2(KEYINPUT115), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n978), .A2(KEYINPUT115), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n961), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1022), .B1(new_n964), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1021), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1002), .A2(new_n1006), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1000), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT122), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT122), .ZN(new_n1029));
  AOI211_X1 g604(.A(new_n1029), .B(new_n1000), .C1(new_n1002), .C2(new_n1006), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT62), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1025), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n984), .B1(new_n1009), .B2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(G299), .B(KEYINPUT57), .ZN(new_n1035));
  INV_X1    g610(.A(G1956), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1011), .A2(new_n1036), .ZN(new_n1037));
  XNOR2_X1  g612(.A(KEYINPUT56), .B(G2072), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n985), .A2(new_n911), .A3(new_n986), .A4(new_n1038), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1037), .A2(KEYINPUT118), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT118), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1035), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  OAI211_X1 g619(.A(KEYINPUT119), .B(new_n1035), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT117), .ZN(new_n1046));
  OAI22_X1  g621(.A1(new_n995), .A2(G1348), .B1(G2067), .B2(new_n952), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1046), .B1(new_n1047), .B2(new_n859), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n951), .A2(new_n911), .ZN(new_n1049));
  AOI22_X1  g624(.A1(new_n717), .A2(new_n973), .B1(new_n1049), .B2(new_n729), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1050), .A2(KEYINPUT117), .A3(new_n591), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1044), .A2(new_n1045), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(new_n1035), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1053), .A2(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1055), .B(KEYINPUT61), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1054), .A2(new_n1035), .ZN(new_n1059));
  XOR2_X1   g634(.A(KEYINPUT58), .B(G1341), .Z(new_n1060));
  NAND2_X1  g635(.A1(new_n952), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n985), .A2(new_n911), .A3(new_n986), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(new_n1062), .B2(G1996), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1063), .A2(new_n1064), .A3(new_n549), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT59), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1063), .A2(new_n1064), .A3(new_n1067), .A4(new_n549), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1059), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1050), .A2(KEYINPUT60), .A3(new_n591), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT60), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n591), .B1(new_n1047), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1072), .B1(new_n1071), .B2(new_n1047), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1058), .A2(new_n1069), .A3(new_n1070), .A4(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1057), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n910), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT123), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n462), .B1(new_n474), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1079), .B2(new_n474), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1078), .B(new_n1081), .C1(new_n951), .C2(KEYINPUT45), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT124), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT124), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n908), .A2(new_n1084), .A3(new_n1078), .A4(new_n1081), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1083), .A2(new_n1085), .A3(new_n985), .A4(new_n991), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1086), .A2(new_n989), .A3(G301), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n994), .A2(new_n1087), .ZN(new_n1088));
  OAI22_X1  g663(.A1(new_n1028), .A2(new_n1030), .B1(KEYINPUT54), .B2(new_n1088), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1086), .A2(new_n989), .A3(KEYINPUT125), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT125), .B1(new_n1086), .B2(new_n989), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1090), .A2(new_n1091), .A3(G301), .ZN(new_n1092));
  OAI21_X1  g667(.A(KEYINPUT54), .B1(new_n993), .B2(G171), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1021), .B(new_n1024), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1089), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1057), .A2(new_n1074), .A3(KEYINPUT121), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1077), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n998), .A2(new_n961), .A3(G286), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1021), .A2(new_n1098), .A3(new_n1024), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT116), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT63), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT116), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1021), .A2(new_n1102), .A3(new_n1098), .A4(new_n1024), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1100), .A2(new_n1101), .A3(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(G8), .B1(new_n977), .B2(new_n974), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1105), .A2(new_n962), .A3(new_n963), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n1106), .A2(new_n1098), .ZN(new_n1107));
  INV_X1    g682(.A(new_n983), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1107), .A2(KEYINPUT63), .A3(new_n978), .A4(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1104), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1034), .A2(new_n1097), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT126), .ZN(new_n1112));
  XOR2_X1   g687(.A(G290), .B(G1986), .Z(new_n1113));
  OAI21_X1  g688(.A(new_n930), .B1(new_n912), .B2(new_n1113), .ZN(new_n1114));
  XOR2_X1   g689(.A(new_n1114), .B(KEYINPUT111), .Z(new_n1115));
  AND3_X1   g690(.A1(new_n1111), .A2(new_n1112), .A3(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1112), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n936), .B1(new_n1116), .B2(new_n1117), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g693(.A1(new_n851), .A2(new_n636), .A3(new_n653), .ZN(new_n1120));
  NAND2_X1  g694(.A1(new_n902), .A2(new_n904), .ZN(new_n1121));
  NOR2_X1   g695(.A1(G229), .A2(new_n460), .ZN(new_n1122));
  AND3_X1   g696(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(G308));
  NAND3_X1  g697(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(G225));
endmodule


