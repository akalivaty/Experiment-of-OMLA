//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 0 1 0 0 1 0 0 0 1 1 0 1 0 1 0 1 0 1 0 0 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n823, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT22), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n202), .A3(new_n206), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G148gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT82), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT82), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G141gat), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT83), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(KEYINPUT80), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT80), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G141gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n222), .A3(G148gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT81), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT82), .B(G148gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT83), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(new_n227), .A3(G141gat), .ZN(new_n228));
  NAND4_X1  g027(.A1(new_n220), .A2(new_n222), .A3(KEYINPUT81), .A4(G148gat), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n219), .A2(new_n225), .A3(new_n228), .A4(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G155gat), .B(G162gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(KEYINPUT84), .A2(G155gat), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n232), .B1(KEYINPUT2), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n236));
  XOR2_X1   g035(.A(G141gat), .B(G148gat), .Z(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT79), .B(KEYINPUT2), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n231), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n235), .A2(new_n236), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT85), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n239), .B1(new_n230), .B2(new_n234), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n244), .A2(KEYINPUT85), .A3(new_n236), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT29), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n212), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G228gat), .ZN(new_n249));
  INV_X1    g048(.A(G233gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT3), .B1(new_n212), .B2(new_n247), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n244), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(KEYINPUT89), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT89), .ZN(new_n255));
  NOR3_X1   g054(.A1(new_n244), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n251), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n248), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT88), .ZN(new_n259));
  AND4_X1   g058(.A1(KEYINPUT85), .A2(new_n235), .A3(new_n236), .A4(new_n240), .ZN(new_n260));
  AOI21_X1  g059(.A(KEYINPUT85), .B1(new_n244), .B2(new_n236), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n247), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n212), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n253), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n259), .B1(new_n264), .B2(new_n251), .ZN(new_n265));
  INV_X1    g064(.A(new_n251), .ZN(new_n266));
  OAI211_X1 g065(.A(KEYINPUT88), .B(new_n266), .C1(new_n248), .C2(new_n253), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n258), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(G22gat), .ZN(new_n269));
  AOI21_X1  g068(.A(KEYINPUT90), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G78gat), .B(G106gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT31), .B(G50gat), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n271), .B(new_n272), .Z(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n265), .A2(new_n267), .ZN(new_n275));
  INV_X1    g074(.A(new_n258), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n269), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AOI211_X1 g076(.A(G22gat), .B(new_n258), .C1(new_n265), .C2(new_n267), .ZN(new_n278));
  OAI22_X1  g077(.A1(new_n270), .A2(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(new_n276), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(G22gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n268), .A2(new_n269), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n281), .A2(KEYINPUT90), .A3(new_n282), .A4(new_n273), .ZN(new_n283));
  INV_X1    g082(.A(G134gat), .ZN(new_n284));
  NOR3_X1   g083(.A1(new_n284), .A2(KEYINPUT70), .A3(G127gat), .ZN(new_n285));
  XNOR2_X1  g084(.A(G127gat), .B(G134gat), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n285), .B1(new_n286), .B2(KEYINPUT70), .ZN(new_n287));
  XNOR2_X1  g086(.A(G113gat), .B(G120gat), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n287), .B1(KEYINPUT1), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G113gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(G120gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT71), .B(G120gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n291), .B1(new_n292), .B2(new_n290), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT1), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n293), .A2(new_n294), .A3(new_n286), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n296), .B1(new_n244), .B2(new_n236), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n297), .B1(new_n243), .B2(new_n245), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n296), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(new_n244), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT4), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n300), .A2(new_n244), .A3(KEYINPUT4), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(G225gat), .A2(G233gat), .ZN(new_n307));
  NAND4_X1  g106(.A1(new_n299), .A2(new_n306), .A3(KEYINPUT5), .A4(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n307), .ZN(new_n309));
  NOR3_X1   g108(.A1(new_n298), .A2(new_n305), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT5), .ZN(new_n311));
  INV_X1    g110(.A(new_n244), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n296), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n301), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n311), .B1(new_n314), .B2(new_n309), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n308), .B1(new_n310), .B2(new_n315), .ZN(new_n316));
  XNOR2_X1  g115(.A(G57gat), .B(G85gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT87), .ZN(new_n318));
  XNOR2_X1  g117(.A(new_n317), .B(new_n318), .ZN(new_n319));
  XOR2_X1   g118(.A(G1gat), .B(G29gat), .Z(new_n320));
  XNOR2_X1  g119(.A(new_n319), .B(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n316), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT92), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n323), .B(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n327), .B(new_n308), .C1(new_n310), .C2(new_n315), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT6), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n325), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n316), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(KEYINPUT6), .A3(new_n323), .ZN(new_n332));
  AOI21_X1  g131(.A(KEYINPUT35), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n279), .A2(new_n283), .A3(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G8gat), .B(G36gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(G64gat), .B(G92gat), .ZN(new_n336));
  XOR2_X1   g135(.A(new_n335), .B(new_n336), .Z(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(G183gat), .ZN(new_n339));
  INV_X1    g138(.A(G190gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n339), .A2(new_n340), .A3(KEYINPUT67), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT67), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n342), .B1(G183gat), .B2(G190gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  AND3_X1   g143(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT23), .ZN(new_n349));
  NOR3_X1   g148(.A1(new_n349), .A2(G169gat), .A3(G176gat), .ZN(new_n350));
  INV_X1    g149(.A(G169gat), .ZN(new_n351));
  INV_X1    g150(.A(G176gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT23), .B1(new_n351), .B2(new_n352), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n350), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n348), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT25), .ZN(new_n357));
  NOR2_X1   g156(.A1(G183gat), .A2(G190gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(G183gat), .A2(G190gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT24), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT66), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n358), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(KEYINPUT65), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT65), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n366), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n346), .A2(KEYINPUT66), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n363), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT25), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(new_n371), .A3(new_n355), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT69), .A4(KEYINPUT26), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT69), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT26), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n376), .B1(new_n351), .B2(new_n352), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n359), .B(new_n374), .C1(new_n375), .C2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT28), .ZN(new_n379));
  XNOR2_X1  g178(.A(KEYINPUT27), .B(G183gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(KEYINPUT68), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n339), .A2(KEYINPUT27), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(KEYINPUT68), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(new_n340), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n379), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT27), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(G183gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n382), .A2(new_n387), .ZN(new_n388));
  NOR3_X1   g187(.A1(new_n388), .A2(new_n379), .A3(G190gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n378), .B1(new_n385), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n373), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G226gat), .A2(G233gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT76), .B1(new_n373), .B2(new_n391), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n375), .A2(new_n377), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n374), .A2(new_n359), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT68), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n388), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(G190gat), .B1(new_n382), .B2(KEYINPUT68), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT28), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n396), .B(new_n397), .C1(new_n401), .C2(new_n389), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT76), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n402), .A2(new_n403), .A3(new_n357), .A4(new_n372), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n395), .A2(new_n247), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n393), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n394), .B1(new_n406), .B2(KEYINPUT77), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT77), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n405), .A2(new_n408), .A3(new_n393), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n212), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n404), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n411), .A2(G226gat), .A3(G233gat), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n247), .B(new_n393), .C1(new_n373), .C2(new_n391), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n263), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n338), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n414), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n405), .A2(new_n408), .A3(new_n393), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n408), .B1(new_n405), .B2(new_n393), .ZN(new_n418));
  NOR3_X1   g217(.A1(new_n417), .A2(new_n418), .A3(new_n394), .ZN(new_n419));
  OAI211_X1 g218(.A(new_n416), .B(new_n337), .C1(new_n419), .C2(new_n212), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT30), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n421), .A2(KEYINPUT78), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n415), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n410), .A2(new_n414), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT78), .B(KEYINPUT30), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n337), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT91), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n423), .A2(new_n426), .A3(KEYINPUT91), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n300), .B1(new_n373), .B2(new_n391), .ZN(new_n432));
  NAND2_X1  g231(.A1(G227gat), .A2(G233gat), .ZN(new_n433));
  XOR2_X1   g232(.A(new_n433), .B(KEYINPUT64), .Z(new_n434));
  NAND4_X1  g233(.A1(new_n402), .A2(new_n296), .A3(new_n357), .A4(new_n372), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT72), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n432), .A2(new_n435), .A3(KEYINPUT72), .A4(new_n434), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT33), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OR2_X1    g239(.A1(new_n440), .A2(KEYINPUT73), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n438), .A2(new_n439), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT32), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT74), .ZN(new_n444));
  XNOR2_X1  g243(.A(G15gat), .B(G43gat), .ZN(new_n445));
  XNOR2_X1  g244(.A(new_n445), .B(KEYINPUT75), .ZN(new_n446));
  XNOR2_X1  g245(.A(G71gat), .B(G99gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n448), .B1(new_n440), .B2(KEYINPUT73), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT74), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n442), .A2(new_n450), .A3(KEYINPUT32), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n441), .A2(new_n444), .A3(new_n449), .A4(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT33), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n442), .B(KEYINPUT32), .C1(new_n453), .C2(new_n448), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT34), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n432), .A2(new_n435), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n457), .A2(new_n434), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT34), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n452), .A2(new_n459), .A3(new_n454), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n456), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n458), .ZN(new_n462));
  INV_X1    g261(.A(new_n460), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n459), .B1(new_n452), .B2(new_n454), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n334), .A2(new_n431), .A3(new_n461), .A4(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT93), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n279), .A2(new_n283), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n331), .A2(new_n323), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n469), .A2(new_n329), .A3(new_n325), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n470), .A2(new_n332), .B1(new_n423), .B2(new_n426), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n468), .A2(new_n461), .A3(new_n465), .A4(new_n471), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n466), .A2(new_n467), .B1(new_n472), .B2(KEYINPUT35), .ZN(new_n473));
  NOR3_X1   g272(.A1(new_n463), .A2(new_n464), .A3(new_n462), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n458), .B1(new_n456), .B2(new_n460), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n476), .A2(KEYINPUT93), .A3(new_n431), .A4(new_n334), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n309), .B1(new_n298), .B2(new_n305), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n313), .A2(new_n307), .A3(new_n301), .ZN(new_n479));
  AND2_X1   g278(.A1(new_n479), .A2(KEYINPUT39), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n327), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n481), .B1(KEYINPUT39), .B2(new_n478), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT40), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n328), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n484), .B1(new_n483), .B2(new_n482), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n485), .A2(new_n429), .A3(new_n430), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT37), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n337), .B1(new_n424), .B2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n488), .B1(new_n487), .B2(new_n424), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT38), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n419), .A2(new_n263), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n412), .A2(new_n413), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n487), .B1(new_n492), .B2(new_n263), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT38), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(new_n488), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n330), .A2(new_n332), .A3(new_n420), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n490), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n486), .A2(new_n497), .A3(new_n468), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n471), .B1(new_n283), .B2(new_n279), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT36), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n474), .B2(new_n475), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n465), .A2(new_n461), .A3(KEYINPUT36), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n473), .A2(new_n477), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G43gat), .B(G50gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT15), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT98), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n506), .B(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(KEYINPUT97), .B(G36gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(G29gat), .ZN(new_n510));
  OR3_X1    g309(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n510), .B(new_n513), .C1(KEYINPUT15), .C2(new_n505), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n508), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n512), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n516), .B1(new_n511), .B2(KEYINPUT96), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n517), .B1(KEYINPUT96), .B2(new_n511), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n506), .B1(new_n518), .B2(new_n510), .ZN(new_n519));
  OR2_X1    g318(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT17), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G15gat), .B(G22gat), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT16), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n523), .B1(new_n524), .B2(G1gat), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n525), .B1(G1gat), .B2(new_n523), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n526), .B(G8gat), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n515), .A2(new_n519), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT17), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n522), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(G229gat), .A2(G233gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n520), .A2(new_n527), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(KEYINPUT99), .A2(KEYINPUT18), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n527), .B1(new_n520), .B2(new_n521), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n537), .A2(new_n530), .B1(new_n520), .B2(new_n527), .ZN(new_n538));
  INV_X1    g337(.A(new_n535), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(new_n532), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n529), .A2(new_n528), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n533), .A2(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n532), .B(KEYINPUT13), .Z(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n536), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT95), .ZN(new_n546));
  XNOR2_X1  g345(.A(G113gat), .B(G141gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT94), .B(G197gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT11), .B(G169gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT12), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n545), .A2(new_n546), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n552), .B1(new_n545), .B2(new_n546), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n504), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G71gat), .B(G78gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n559), .A2(KEYINPUT100), .ZN(new_n560));
  AOI21_X1  g359(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(G57gat), .B(G64gat), .ZN(new_n562));
  NOR3_X1   g361(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n559), .A2(KEYINPUT100), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI211_X1 g364(.A(KEYINPUT100), .B(new_n559), .C1(new_n562), .C2(new_n561), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n567), .A2(KEYINPUT21), .ZN(new_n568));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G127gat), .B(G155gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT20), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n570), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G183gat), .B(G211gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT102), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n573), .B(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n527), .B1(KEYINPUT21), .B2(new_n567), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT101), .B(KEYINPUT19), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n576), .B(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G85gat), .A2(G92gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT7), .ZN(new_n583));
  NAND2_X1  g382(.A1(G99gat), .A2(G106gat), .ZN(new_n584));
  INV_X1    g383(.A(G85gat), .ZN(new_n585));
  INV_X1    g384(.A(G92gat), .ZN(new_n586));
  AOI22_X1  g385(.A1(KEYINPUT8), .A2(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G99gat), .B(G106gat), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n588), .B(new_n589), .Z(new_n590));
  NAND3_X1  g389(.A1(new_n522), .A2(new_n530), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n588), .B(new_n589), .ZN(new_n592));
  AND2_X1   g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(new_n520), .A2(new_n592), .B1(KEYINPUT41), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G190gat), .B(G218gat), .Z(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n593), .A2(KEYINPUT41), .ZN(new_n598));
  XNOR2_X1  g397(.A(G134gat), .B(G162gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n595), .A2(new_n596), .ZN(new_n602));
  OR3_X1    g401(.A1(new_n597), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n601), .B1(new_n602), .B2(new_n597), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n567), .A2(KEYINPUT10), .A3(new_n592), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT104), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n583), .A2(new_n589), .A3(new_n587), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(KEYINPUT103), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n567), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(new_n592), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT10), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n608), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n611), .A2(new_n592), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n590), .B1(new_n567), .B2(new_n610), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n617), .A2(KEYINPUT104), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n607), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G230gat), .A2(G233gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n612), .A2(new_n620), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G120gat), .B(G148gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(G176gat), .B(G204gat), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n625), .B(new_n626), .Z(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n621), .A2(new_n623), .A3(new_n627), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NOR3_X1   g430(.A1(new_n581), .A2(new_n606), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n558), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n470), .A2(new_n332), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g437(.A1(new_n633), .A2(new_n431), .ZN(new_n639));
  XOR2_X1   g438(.A(KEYINPUT16), .B(G8gat), .Z(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT42), .ZN(new_n642));
  INV_X1    g441(.A(new_n639), .ZN(new_n643));
  AOI22_X1  g442(.A1(new_n641), .A2(new_n642), .B1(new_n643), .B2(G8gat), .ZN(new_n644));
  OAI21_X1  g443(.A(KEYINPUT105), .B1(new_n641), .B2(new_n642), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT105), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n639), .A2(new_n646), .A3(KEYINPUT42), .A4(new_n640), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(G1325gat));
  NAND2_X1  g447(.A1(new_n501), .A2(new_n502), .ZN(new_n649));
  OAI21_X1  g448(.A(G15gat), .B1(new_n633), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n476), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n651), .A2(G15gat), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n650), .B1(new_n633), .B2(new_n652), .ZN(G1326gat));
  NOR2_X1   g452(.A1(new_n633), .A2(new_n468), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT43), .B(G22gat), .Z(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(G1327gat));
  NOR2_X1   g455(.A1(new_n580), .A2(new_n631), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n658), .A2(new_n557), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n504), .B2(new_n605), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n466), .A2(new_n467), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n472), .A2(KEYINPUT35), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n664), .A2(new_n477), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n503), .A2(new_n498), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n668), .A2(new_n606), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n660), .B1(new_n663), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n636), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(G29gat), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n605), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n675), .A2(G29gat), .A3(new_n635), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n558), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT45), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n673), .A2(new_n678), .ZN(G1328gat));
  NOR3_X1   g478(.A1(new_n675), .A2(new_n509), .A3(new_n431), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n558), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(KEYINPUT46), .Z(new_n682));
  INV_X1    g481(.A(new_n431), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n671), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT107), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n509), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n684), .A2(KEYINPUT107), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n682), .B1(new_n686), .B2(new_n687), .ZN(G1329gat));
  INV_X1    g487(.A(G43gat), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n558), .A2(new_n689), .A3(new_n476), .A4(new_n674), .ZN(new_n690));
  INV_X1    g489(.A(new_n649), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n671), .A2(new_n691), .ZN(new_n692));
  OAI211_X1 g491(.A(KEYINPUT47), .B(new_n690), .C1(new_n692), .C2(new_n689), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT47), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n689), .B1(new_n671), .B2(new_n691), .ZN(new_n695));
  INV_X1    g494(.A(new_n690), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n694), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n693), .A2(new_n697), .ZN(G1330gat));
  INV_X1    g497(.A(new_n468), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n671), .A2(G50gat), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n558), .A2(new_n699), .A3(new_n674), .ZN(new_n701));
  INV_X1    g500(.A(G50gat), .ZN(new_n702));
  AOI22_X1  g501(.A1(new_n701), .A2(new_n702), .B1(KEYINPUT108), .B2(KEYINPUT48), .ZN(new_n703));
  OR2_X1    g502(.A1(KEYINPUT108), .A2(KEYINPUT48), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n700), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n704), .B1(new_n700), .B2(new_n703), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(G1331gat));
  NAND3_X1  g506(.A1(new_n580), .A2(new_n557), .A3(new_n605), .ZN(new_n708));
  INV_X1    g507(.A(new_n631), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n710), .B(KEYINPUT109), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n504), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(new_n636), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g513(.A(new_n431), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n715), .B(KEYINPUT110), .Z(new_n716));
  NAND2_X1  g515(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT111), .ZN(new_n718));
  NOR2_X1   g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1333gat));
  XOR2_X1   g519(.A(new_n476), .B(KEYINPUT112), .Z(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(G71gat), .B1(new_n712), .B2(new_n722), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n691), .A2(G71gat), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n723), .B1(new_n712), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT50), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1334gat));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n699), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g528(.A1(new_n581), .A2(KEYINPUT113), .A3(new_n557), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT113), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n731), .B1(new_n580), .B2(new_n556), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT114), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT51), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n730), .A2(new_n732), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n668), .A2(new_n606), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n733), .A2(new_n734), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n737), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n668), .A2(new_n606), .A3(new_n735), .A4(new_n739), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n709), .A2(new_n635), .A3(G85gat), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n738), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n730), .A2(new_n732), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n631), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n744), .B1(new_n663), .B2(new_n670), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n745), .A2(new_n636), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n742), .B1(new_n746), .B2(new_n585), .ZN(G1336gat));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n709), .A2(G92gat), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n738), .A2(new_n683), .A3(new_n740), .A4(new_n749), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n745), .A2(new_n683), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n748), .B(new_n750), .C1(new_n751), .C2(new_n586), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n586), .B1(new_n745), .B2(new_n683), .ZN(new_n753));
  INV_X1    g552(.A(new_n750), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT52), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n752), .A2(new_n755), .ZN(G1337gat));
  NOR3_X1   g555(.A1(new_n651), .A2(G99gat), .A3(new_n709), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT116), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n738), .A2(new_n740), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n745), .A2(new_n691), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT115), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G99gat), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n760), .A2(KEYINPUT115), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n759), .B1(new_n762), .B2(new_n763), .ZN(G1338gat));
  INV_X1    g563(.A(KEYINPUT117), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n765), .A2(KEYINPUT53), .ZN(new_n766));
  INV_X1    g565(.A(G106gat), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n468), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n766), .B1(new_n745), .B2(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n468), .A2(new_n709), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n738), .A2(new_n740), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n767), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n765), .A2(KEYINPUT53), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n769), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n773), .B1(new_n769), .B2(new_n772), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(G1339gat));
  NOR2_X1   g575(.A1(new_n708), .A2(new_n631), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779));
  INV_X1    g578(.A(new_n607), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n612), .A2(new_n608), .A3(new_n613), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n617), .A2(KEYINPUT104), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n620), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(KEYINPUT54), .B1(new_n783), .B2(new_n784), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n619), .A2(new_n789), .A3(new_n620), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n628), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n779), .B1(new_n788), .B2(new_n791), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n621), .A2(KEYINPUT54), .A3(new_n785), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n793), .A2(KEYINPUT55), .A3(new_n628), .A4(new_n790), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n792), .A2(new_n630), .A3(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n536), .A2(new_n540), .A3(new_n544), .A4(new_n552), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n538), .A2(new_n532), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n542), .A2(new_n543), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n551), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n606), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n795), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n792), .A2(new_n556), .A3(new_n630), .A4(new_n794), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n627), .B1(new_n621), .B2(new_n623), .ZN(new_n804));
  AOI211_X1 g603(.A(new_n622), .B(new_n628), .C1(new_n619), .C2(new_n620), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n800), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT118), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n631), .A2(new_n808), .A3(new_n800), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n803), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n802), .B1(new_n810), .B2(new_n605), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n778), .B1(new_n811), .B2(new_n580), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n813), .A2(new_n699), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n431), .A2(new_n636), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n651), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n817), .A2(new_n557), .ZN(new_n818));
  XNOR2_X1  g617(.A(new_n818), .B(new_n290), .ZN(G1340gat));
  NOR2_X1   g618(.A1(new_n817), .A2(new_n709), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(G120gat), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(new_n292), .B2(new_n820), .ZN(G1341gat));
  NOR2_X1   g621(.A1(new_n817), .A2(new_n581), .ZN(new_n823));
  XOR2_X1   g622(.A(KEYINPUT119), .B(G127gat), .Z(new_n824));
  XNOR2_X1  g623(.A(new_n823), .B(new_n824), .ZN(G1342gat));
  NOR2_X1   g624(.A1(new_n817), .A2(new_n605), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n284), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT56), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n826), .A2(new_n829), .A3(new_n284), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n828), .B(new_n830), .C1(new_n284), .C2(new_n826), .ZN(G1343gat));
  NAND2_X1  g630(.A1(new_n812), .A2(new_n699), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n649), .A2(new_n636), .A3(new_n431), .ZN(new_n833));
  NOR4_X1   g632(.A1(new_n832), .A2(G141gat), .A3(new_n557), .A4(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(new_n833), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n699), .A2(KEYINPUT57), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n606), .B1(new_n803), .B2(new_n806), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n581), .B1(new_n838), .B2(new_n802), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n777), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI211_X1 g640(.A(KEYINPUT120), .B(new_n581), .C1(new_n838), .C2(new_n802), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n837), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT57), .B1(new_n812), .B2(new_n699), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n556), .B(new_n835), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n220), .A2(new_n222), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n834), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n847), .A2(new_n848), .A3(KEYINPUT58), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(KEYINPUT58), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n848), .A2(KEYINPUT58), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n847), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n849), .A2(new_n852), .ZN(G1344gat));
  NOR2_X1   g652(.A1(new_n832), .A2(new_n833), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n226), .A3(new_n631), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n843), .A2(new_n844), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n856), .A2(new_n833), .ZN(new_n857));
  AOI211_X1 g656(.A(KEYINPUT59), .B(new_n226), .C1(new_n857), .C2(new_n631), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n813), .A2(new_n837), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n839), .A2(new_n778), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT57), .B1(new_n861), .B2(new_n699), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n631), .B(new_n835), .C1(new_n860), .C2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n859), .B1(new_n863), .B2(G148gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n855), .B1(new_n858), .B2(new_n864), .ZN(G1345gat));
  NAND2_X1  g664(.A1(new_n854), .A2(new_n580), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n866), .B(KEYINPUT122), .ZN(new_n867));
  XOR2_X1   g666(.A(KEYINPUT84), .B(G155gat), .Z(new_n868));
  NOR2_X1   g667(.A1(new_n581), .A2(new_n868), .ZN(new_n869));
  AOI22_X1  g668(.A1(new_n867), .A2(new_n868), .B1(new_n857), .B2(new_n869), .ZN(G1346gat));
  INV_X1    g669(.A(G162gat), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n606), .B(new_n835), .C1(new_n843), .C2(new_n844), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n873), .B2(new_n872), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n635), .A2(new_n605), .A3(G162gat), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n649), .A2(new_n431), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n875), .B1(new_n832), .B2(new_n877), .ZN(G1347gat));
  NOR3_X1   g677(.A1(new_n721), .A2(new_n636), .A3(new_n431), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n814), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n880), .A2(new_n351), .A3(new_n557), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n813), .A2(new_n636), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n651), .A2(new_n699), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(KEYINPUT124), .A3(new_n683), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT124), .ZN(new_n885));
  INV_X1    g684(.A(new_n883), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n885), .B1(new_n886), .B2(new_n431), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n882), .A2(new_n884), .A3(new_n887), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n888), .A2(KEYINPUT125), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(KEYINPUT125), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n889), .A2(new_n556), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n881), .B1(new_n891), .B2(new_n351), .ZN(G1348gat));
  OAI21_X1  g691(.A(G176gat), .B1(new_n880), .B2(new_n709), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n889), .A2(new_n890), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n631), .A2(new_n352), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(G1349gat));
  OAI21_X1  g695(.A(G183gat), .B1(new_n880), .B2(new_n581), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n581), .A2(new_n388), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n897), .B1(new_n888), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT60), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT60), .ZN(new_n902));
  OAI211_X1 g701(.A(new_n897), .B(new_n902), .C1(new_n888), .C2(new_n899), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n880), .B2(new_n605), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(KEYINPUT61), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n905), .A2(KEYINPUT61), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n606), .A2(new_n340), .ZN(new_n908));
  OAI22_X1  g707(.A1(new_n906), .A2(new_n907), .B1(new_n894), .B2(new_n908), .ZN(G1351gat));
  NAND3_X1  g708(.A1(new_n649), .A2(new_n635), .A3(new_n683), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n832), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(G197gat), .B1(new_n911), .B2(new_n556), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n860), .A2(new_n862), .ZN(new_n913));
  INV_X1    g712(.A(G197gat), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n913), .A2(new_n914), .A3(new_n557), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n910), .B(KEYINPUT126), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n912), .B1(new_n915), .B2(new_n917), .ZN(G1352gat));
  NOR4_X1   g717(.A1(new_n832), .A2(G204gat), .A3(new_n709), .A4(new_n910), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT62), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n631), .B1(new_n860), .B2(new_n862), .ZN(new_n921));
  OAI21_X1  g720(.A(G204gat), .B1(new_n921), .B2(new_n916), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1353gat));
  NAND3_X1  g722(.A1(new_n911), .A2(new_n204), .A3(new_n580), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n910), .A2(new_n581), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n925), .B1(new_n860), .B2(new_n862), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n926), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT63), .B1(new_n926), .B2(G211gat), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n924), .B1(new_n927), .B2(new_n928), .ZN(G1354gat));
  AOI21_X1  g728(.A(G218gat), .B1(new_n911), .B2(new_n606), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n913), .A2(new_n205), .A3(new_n605), .ZN(new_n934));
  AOI22_X1  g733(.A1(new_n932), .A2(new_n933), .B1(new_n934), .B2(new_n917), .ZN(G1355gat));
endmodule


